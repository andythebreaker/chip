`define size_minus_1(x) (x-1)
`define matrix_size_1 100
`define matrix_size_2 400
`define vector_size `matrix_size_1

module vector_add_vector_genED_X_100_400_V_100 (
input logic signed [31:0] a[0:`size_minus_1(`vector_size)],
input logic signed [31:0] b[0:`size_minus_1(`vector_size)],
output logic signed [31:0] result[0:`size_minus_1(`vector_size)]
);
assign result[0] = a[0] + b[0];
assign result[1] = a[1] + b[1];
assign result[2] = a[2] + b[2];
assign result[3] = a[3] + b[3];
assign result[4] = a[4] + b[4];
assign result[5] = a[5] + b[5];
assign result[6] = a[6] + b[6];
assign result[7] = a[7] + b[7];
assign result[8] = a[8] + b[8];
assign result[9] = a[9] + b[9];
assign result[10] = a[10] + b[10];
assign result[11] = a[11] + b[11];
assign result[12] = a[12] + b[12];
assign result[13] = a[13] + b[13];
assign result[14] = a[14] + b[14];
assign result[15] = a[15] + b[15];
assign result[16] = a[16] + b[16];
assign result[17] = a[17] + b[17];
assign result[18] = a[18] + b[18];
assign result[19] = a[19] + b[19];
assign result[20] = a[20] + b[20];
assign result[21] = a[21] + b[21];
assign result[22] = a[22] + b[22];
assign result[23] = a[23] + b[23];
assign result[24] = a[24] + b[24];
assign result[25] = a[25] + b[25];
assign result[26] = a[26] + b[26];
assign result[27] = a[27] + b[27];
assign result[28] = a[28] + b[28];
assign result[29] = a[29] + b[29];
assign result[30] = a[30] + b[30];
assign result[31] = a[31] + b[31];
assign result[32] = a[32] + b[32];
assign result[33] = a[33] + b[33];
assign result[34] = a[34] + b[34];
assign result[35] = a[35] + b[35];
assign result[36] = a[36] + b[36];
assign result[37] = a[37] + b[37];
assign result[38] = a[38] + b[38];
assign result[39] = a[39] + b[39];
assign result[40] = a[40] + b[40];
assign result[41] = a[41] + b[41];
assign result[42] = a[42] + b[42];
assign result[43] = a[43] + b[43];
assign result[44] = a[44] + b[44];
assign result[45] = a[45] + b[45];
assign result[46] = a[46] + b[46];
assign result[47] = a[47] + b[47];
assign result[48] = a[48] + b[48];
assign result[49] = a[49] + b[49];
assign result[50] = a[50] + b[50];
assign result[51] = a[51] + b[51];
assign result[52] = a[52] + b[52];
assign result[53] = a[53] + b[53];
assign result[54] = a[54] + b[54];
assign result[55] = a[55] + b[55];
assign result[56] = a[56] + b[56];
assign result[57] = a[57] + b[57];
assign result[58] = a[58] + b[58];
assign result[59] = a[59] + b[59];
assign result[60] = a[60] + b[60];
assign result[61] = a[61] + b[61];
assign result[62] = a[62] + b[62];
assign result[63] = a[63] + b[63];
assign result[64] = a[64] + b[64];
assign result[65] = a[65] + b[65];
assign result[66] = a[66] + b[66];
assign result[67] = a[67] + b[67];
assign result[68] = a[68] + b[68];
assign result[69] = a[69] + b[69];
assign result[70] = a[70] + b[70];
assign result[71] = a[71] + b[71];
assign result[72] = a[72] + b[72];
assign result[73] = a[73] + b[73];
assign result[74] = a[74] + b[74];
assign result[75] = a[75] + b[75];
assign result[76] = a[76] + b[76];
assign result[77] = a[77] + b[77];
assign result[78] = a[78] + b[78];
assign result[79] = a[79] + b[79];
assign result[80] = a[80] + b[80];
assign result[81] = a[81] + b[81];
assign result[82] = a[82] + b[82];
assign result[83] = a[83] + b[83];
assign result[84] = a[84] + b[84];
assign result[85] = a[85] + b[85];
assign result[86] = a[86] + b[86];
assign result[87] = a[87] + b[87];
assign result[88] = a[88] + b[88];
assign result[89] = a[89] + b[89];
assign result[90] = a[90] + b[90];
assign result[91] = a[91] + b[91];
assign result[92] = a[92] + b[92];
assign result[93] = a[93] + b[93];
assign result[94] = a[94] + b[94];
assign result[95] = a[95] + b[95];
assign result[96] = a[96] + b[96];
assign result[97] = a[97] + b[97];
assign result[98] = a[98] + b[98];
assign result[99] = a[99] + b[99];

endmodule
