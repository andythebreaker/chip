module float_mat_mux(
    input a,
    input b,
    output c
);
    
endmodule