`define size_minus_1(x) (x-1)
`define matrix_size_1 100
`define matrix_size_2 400
`define vector_size `matrix_size_1

module vector_add_vector_genED_M_100_400_X_400 (
input logic signed [31:0] a[0:`size_minus_1(`matrix_size_2)],
input logic signed [31:0] b[0:`size_minus_1(`matrix_size_2)],
output logic signed [31:0] result[0:`size_minus_1(`matrix_size_2)]
);
assign result[0] = a[0] + b[0];
assign result[1] = a[1] + b[1];
assign result[2] = a[2] + b[2];
assign result[3] = a[3] + b[3];
assign result[4] = a[4] + b[4];
assign result[5] = a[5] + b[5];
assign result[6] = a[6] + b[6];
assign result[7] = a[7] + b[7];
assign result[8] = a[8] + b[8];
assign result[9] = a[9] + b[9];
assign result[10] = a[10] + b[10];
assign result[11] = a[11] + b[11];
assign result[12] = a[12] + b[12];
assign result[13] = a[13] + b[13];
assign result[14] = a[14] + b[14];
assign result[15] = a[15] + b[15];
assign result[16] = a[16] + b[16];
assign result[17] = a[17] + b[17];
assign result[18] = a[18] + b[18];
assign result[19] = a[19] + b[19];
assign result[20] = a[20] + b[20];
assign result[21] = a[21] + b[21];
assign result[22] = a[22] + b[22];
assign result[23] = a[23] + b[23];
assign result[24] = a[24] + b[24];
assign result[25] = a[25] + b[25];
assign result[26] = a[26] + b[26];
assign result[27] = a[27] + b[27];
assign result[28] = a[28] + b[28];
assign result[29] = a[29] + b[29];
assign result[30] = a[30] + b[30];
assign result[31] = a[31] + b[31];
assign result[32] = a[32] + b[32];
assign result[33] = a[33] + b[33];
assign result[34] = a[34] + b[34];
assign result[35] = a[35] + b[35];
assign result[36] = a[36] + b[36];
assign result[37] = a[37] + b[37];
assign result[38] = a[38] + b[38];
assign result[39] = a[39] + b[39];
assign result[40] = a[40] + b[40];
assign result[41] = a[41] + b[41];
assign result[42] = a[42] + b[42];
assign result[43] = a[43] + b[43];
assign result[44] = a[44] + b[44];
assign result[45] = a[45] + b[45];
assign result[46] = a[46] + b[46];
assign result[47] = a[47] + b[47];
assign result[48] = a[48] + b[48];
assign result[49] = a[49] + b[49];
assign result[50] = a[50] + b[50];
assign result[51] = a[51] + b[51];
assign result[52] = a[52] + b[52];
assign result[53] = a[53] + b[53];
assign result[54] = a[54] + b[54];
assign result[55] = a[55] + b[55];
assign result[56] = a[56] + b[56];
assign result[57] = a[57] + b[57];
assign result[58] = a[58] + b[58];
assign result[59] = a[59] + b[59];
assign result[60] = a[60] + b[60];
assign result[61] = a[61] + b[61];
assign result[62] = a[62] + b[62];
assign result[63] = a[63] + b[63];
assign result[64] = a[64] + b[64];
assign result[65] = a[65] + b[65];
assign result[66] = a[66] + b[66];
assign result[67] = a[67] + b[67];
assign result[68] = a[68] + b[68];
assign result[69] = a[69] + b[69];
assign result[70] = a[70] + b[70];
assign result[71] = a[71] + b[71];
assign result[72] = a[72] + b[72];
assign result[73] = a[73] + b[73];
assign result[74] = a[74] + b[74];
assign result[75] = a[75] + b[75];
assign result[76] = a[76] + b[76];
assign result[77] = a[77] + b[77];
assign result[78] = a[78] + b[78];
assign result[79] = a[79] + b[79];
assign result[80] = a[80] + b[80];
assign result[81] = a[81] + b[81];
assign result[82] = a[82] + b[82];
assign result[83] = a[83] + b[83];
assign result[84] = a[84] + b[84];
assign result[85] = a[85] + b[85];
assign result[86] = a[86] + b[86];
assign result[87] = a[87] + b[87];
assign result[88] = a[88] + b[88];
assign result[89] = a[89] + b[89];
assign result[90] = a[90] + b[90];
assign result[91] = a[91] + b[91];
assign result[92] = a[92] + b[92];
assign result[93] = a[93] + b[93];
assign result[94] = a[94] + b[94];
assign result[95] = a[95] + b[95];
assign result[96] = a[96] + b[96];
assign result[97] = a[97] + b[97];
assign result[98] = a[98] + b[98];
assign result[99] = a[99] + b[99];
assign result[100] = a[100] + b[100];
assign result[101] = a[101] + b[101];
assign result[102] = a[102] + b[102];
assign result[103] = a[103] + b[103];
assign result[104] = a[104] + b[104];
assign result[105] = a[105] + b[105];
assign result[106] = a[106] + b[106];
assign result[107] = a[107] + b[107];
assign result[108] = a[108] + b[108];
assign result[109] = a[109] + b[109];
assign result[110] = a[110] + b[110];
assign result[111] = a[111] + b[111];
assign result[112] = a[112] + b[112];
assign result[113] = a[113] + b[113];
assign result[114] = a[114] + b[114];
assign result[115] = a[115] + b[115];
assign result[116] = a[116] + b[116];
assign result[117] = a[117] + b[117];
assign result[118] = a[118] + b[118];
assign result[119] = a[119] + b[119];
assign result[120] = a[120] + b[120];
assign result[121] = a[121] + b[121];
assign result[122] = a[122] + b[122];
assign result[123] = a[123] + b[123];
assign result[124] = a[124] + b[124];
assign result[125] = a[125] + b[125];
assign result[126] = a[126] + b[126];
assign result[127] = a[127] + b[127];
assign result[128] = a[128] + b[128];
assign result[129] = a[129] + b[129];
assign result[130] = a[130] + b[130];
assign result[131] = a[131] + b[131];
assign result[132] = a[132] + b[132];
assign result[133] = a[133] + b[133];
assign result[134] = a[134] + b[134];
assign result[135] = a[135] + b[135];
assign result[136] = a[136] + b[136];
assign result[137] = a[137] + b[137];
assign result[138] = a[138] + b[138];
assign result[139] = a[139] + b[139];
assign result[140] = a[140] + b[140];
assign result[141] = a[141] + b[141];
assign result[142] = a[142] + b[142];
assign result[143] = a[143] + b[143];
assign result[144] = a[144] + b[144];
assign result[145] = a[145] + b[145];
assign result[146] = a[146] + b[146];
assign result[147] = a[147] + b[147];
assign result[148] = a[148] + b[148];
assign result[149] = a[149] + b[149];
assign result[150] = a[150] + b[150];
assign result[151] = a[151] + b[151];
assign result[152] = a[152] + b[152];
assign result[153] = a[153] + b[153];
assign result[154] = a[154] + b[154];
assign result[155] = a[155] + b[155];
assign result[156] = a[156] + b[156];
assign result[157] = a[157] + b[157];
assign result[158] = a[158] + b[158];
assign result[159] = a[159] + b[159];
assign result[160] = a[160] + b[160];
assign result[161] = a[161] + b[161];
assign result[162] = a[162] + b[162];
assign result[163] = a[163] + b[163];
assign result[164] = a[164] + b[164];
assign result[165] = a[165] + b[165];
assign result[166] = a[166] + b[166];
assign result[167] = a[167] + b[167];
assign result[168] = a[168] + b[168];
assign result[169] = a[169] + b[169];
assign result[170] = a[170] + b[170];
assign result[171] = a[171] + b[171];
assign result[172] = a[172] + b[172];
assign result[173] = a[173] + b[173];
assign result[174] = a[174] + b[174];
assign result[175] = a[175] + b[175];
assign result[176] = a[176] + b[176];
assign result[177] = a[177] + b[177];
assign result[178] = a[178] + b[178];
assign result[179] = a[179] + b[179];
assign result[180] = a[180] + b[180];
assign result[181] = a[181] + b[181];
assign result[182] = a[182] + b[182];
assign result[183] = a[183] + b[183];
assign result[184] = a[184] + b[184];
assign result[185] = a[185] + b[185];
assign result[186] = a[186] + b[186];
assign result[187] = a[187] + b[187];
assign result[188] = a[188] + b[188];
assign result[189] = a[189] + b[189];
assign result[190] = a[190] + b[190];
assign result[191] = a[191] + b[191];
assign result[192] = a[192] + b[192];
assign result[193] = a[193] + b[193];
assign result[194] = a[194] + b[194];
assign result[195] = a[195] + b[195];
assign result[196] = a[196] + b[196];
assign result[197] = a[197] + b[197];
assign result[198] = a[198] + b[198];
assign result[199] = a[199] + b[199];
assign result[200] = a[200] + b[200];
assign result[201] = a[201] + b[201];
assign result[202] = a[202] + b[202];
assign result[203] = a[203] + b[203];
assign result[204] = a[204] + b[204];
assign result[205] = a[205] + b[205];
assign result[206] = a[206] + b[206];
assign result[207] = a[207] + b[207];
assign result[208] = a[208] + b[208];
assign result[209] = a[209] + b[209];
assign result[210] = a[210] + b[210];
assign result[211] = a[211] + b[211];
assign result[212] = a[212] + b[212];
assign result[213] = a[213] + b[213];
assign result[214] = a[214] + b[214];
assign result[215] = a[215] + b[215];
assign result[216] = a[216] + b[216];
assign result[217] = a[217] + b[217];
assign result[218] = a[218] + b[218];
assign result[219] = a[219] + b[219];
assign result[220] = a[220] + b[220];
assign result[221] = a[221] + b[221];
assign result[222] = a[222] + b[222];
assign result[223] = a[223] + b[223];
assign result[224] = a[224] + b[224];
assign result[225] = a[225] + b[225];
assign result[226] = a[226] + b[226];
assign result[227] = a[227] + b[227];
assign result[228] = a[228] + b[228];
assign result[229] = a[229] + b[229];
assign result[230] = a[230] + b[230];
assign result[231] = a[231] + b[231];
assign result[232] = a[232] + b[232];
assign result[233] = a[233] + b[233];
assign result[234] = a[234] + b[234];
assign result[235] = a[235] + b[235];
assign result[236] = a[236] + b[236];
assign result[237] = a[237] + b[237];
assign result[238] = a[238] + b[238];
assign result[239] = a[239] + b[239];
assign result[240] = a[240] + b[240];
assign result[241] = a[241] + b[241];
assign result[242] = a[242] + b[242];
assign result[243] = a[243] + b[243];
assign result[244] = a[244] + b[244];
assign result[245] = a[245] + b[245];
assign result[246] = a[246] + b[246];
assign result[247] = a[247] + b[247];
assign result[248] = a[248] + b[248];
assign result[249] = a[249] + b[249];
assign result[250] = a[250] + b[250];
assign result[251] = a[251] + b[251];
assign result[252] = a[252] + b[252];
assign result[253] = a[253] + b[253];
assign result[254] = a[254] + b[254];
assign result[255] = a[255] + b[255];
assign result[256] = a[256] + b[256];
assign result[257] = a[257] + b[257];
assign result[258] = a[258] + b[258];
assign result[259] = a[259] + b[259];
assign result[260] = a[260] + b[260];
assign result[261] = a[261] + b[261];
assign result[262] = a[262] + b[262];
assign result[263] = a[263] + b[263];
assign result[264] = a[264] + b[264];
assign result[265] = a[265] + b[265];
assign result[266] = a[266] + b[266];
assign result[267] = a[267] + b[267];
assign result[268] = a[268] + b[268];
assign result[269] = a[269] + b[269];
assign result[270] = a[270] + b[270];
assign result[271] = a[271] + b[271];
assign result[272] = a[272] + b[272];
assign result[273] = a[273] + b[273];
assign result[274] = a[274] + b[274];
assign result[275] = a[275] + b[275];
assign result[276] = a[276] + b[276];
assign result[277] = a[277] + b[277];
assign result[278] = a[278] + b[278];
assign result[279] = a[279] + b[279];
assign result[280] = a[280] + b[280];
assign result[281] = a[281] + b[281];
assign result[282] = a[282] + b[282];
assign result[283] = a[283] + b[283];
assign result[284] = a[284] + b[284];
assign result[285] = a[285] + b[285];
assign result[286] = a[286] + b[286];
assign result[287] = a[287] + b[287];
assign result[288] = a[288] + b[288];
assign result[289] = a[289] + b[289];
assign result[290] = a[290] + b[290];
assign result[291] = a[291] + b[291];
assign result[292] = a[292] + b[292];
assign result[293] = a[293] + b[293];
assign result[294] = a[294] + b[294];
assign result[295] = a[295] + b[295];
assign result[296] = a[296] + b[296];
assign result[297] = a[297] + b[297];
assign result[298] = a[298] + b[298];
assign result[299] = a[299] + b[299];
assign result[300] = a[300] + b[300];
assign result[301] = a[301] + b[301];
assign result[302] = a[302] + b[302];
assign result[303] = a[303] + b[303];
assign result[304] = a[304] + b[304];
assign result[305] = a[305] + b[305];
assign result[306] = a[306] + b[306];
assign result[307] = a[307] + b[307];
assign result[308] = a[308] + b[308];
assign result[309] = a[309] + b[309];
assign result[310] = a[310] + b[310];
assign result[311] = a[311] + b[311];
assign result[312] = a[312] + b[312];
assign result[313] = a[313] + b[313];
assign result[314] = a[314] + b[314];
assign result[315] = a[315] + b[315];
assign result[316] = a[316] + b[316];
assign result[317] = a[317] + b[317];
assign result[318] = a[318] + b[318];
assign result[319] = a[319] + b[319];
assign result[320] = a[320] + b[320];
assign result[321] = a[321] + b[321];
assign result[322] = a[322] + b[322];
assign result[323] = a[323] + b[323];
assign result[324] = a[324] + b[324];
assign result[325] = a[325] + b[325];
assign result[326] = a[326] + b[326];
assign result[327] = a[327] + b[327];
assign result[328] = a[328] + b[328];
assign result[329] = a[329] + b[329];
assign result[330] = a[330] + b[330];
assign result[331] = a[331] + b[331];
assign result[332] = a[332] + b[332];
assign result[333] = a[333] + b[333];
assign result[334] = a[334] + b[334];
assign result[335] = a[335] + b[335];
assign result[336] = a[336] + b[336];
assign result[337] = a[337] + b[337];
assign result[338] = a[338] + b[338];
assign result[339] = a[339] + b[339];
assign result[340] = a[340] + b[340];
assign result[341] = a[341] + b[341];
assign result[342] = a[342] + b[342];
assign result[343] = a[343] + b[343];
assign result[344] = a[344] + b[344];
assign result[345] = a[345] + b[345];
assign result[346] = a[346] + b[346];
assign result[347] = a[347] + b[347];
assign result[348] = a[348] + b[348];
assign result[349] = a[349] + b[349];
assign result[350] = a[350] + b[350];
assign result[351] = a[351] + b[351];
assign result[352] = a[352] + b[352];
assign result[353] = a[353] + b[353];
assign result[354] = a[354] + b[354];
assign result[355] = a[355] + b[355];
assign result[356] = a[356] + b[356];
assign result[357] = a[357] + b[357];
assign result[358] = a[358] + b[358];
assign result[359] = a[359] + b[359];
assign result[360] = a[360] + b[360];
assign result[361] = a[361] + b[361];
assign result[362] = a[362] + b[362];
assign result[363] = a[363] + b[363];
assign result[364] = a[364] + b[364];
assign result[365] = a[365] + b[365];
assign result[366] = a[366] + b[366];
assign result[367] = a[367] + b[367];
assign result[368] = a[368] + b[368];
assign result[369] = a[369] + b[369];
assign result[370] = a[370] + b[370];
assign result[371] = a[371] + b[371];
assign result[372] = a[372] + b[372];
assign result[373] = a[373] + b[373];
assign result[374] = a[374] + b[374];
assign result[375] = a[375] + b[375];
assign result[376] = a[376] + b[376];
assign result[377] = a[377] + b[377];
assign result[378] = a[378] + b[378];
assign result[379] = a[379] + b[379];
assign result[380] = a[380] + b[380];
assign result[381] = a[381] + b[381];
assign result[382] = a[382] + b[382];
assign result[383] = a[383] + b[383];
assign result[384] = a[384] + b[384];
assign result[385] = a[385] + b[385];
assign result[386] = a[386] + b[386];
assign result[387] = a[387] + b[387];
assign result[388] = a[388] + b[388];
assign result[389] = a[389] + b[389];
assign result[390] = a[390] + b[390];
assign result[391] = a[391] + b[391];
assign result[392] = a[392] + b[392];
assign result[393] = a[393] + b[393];
assign result[394] = a[394] + b[394];
assign result[395] = a[395] + b[395];
assign result[396] = a[396] + b[396];
assign result[397] = a[397] + b[397];
assign result[398] = a[398] + b[398];
assign result[399] = a[399] + b[399];

endmodule
