`define size_minus_1(x) (x-1)
`define matrix_size_1 100
`define matrix_size_2 400
`define vector_size `matrix_size_1

module matrix_times_vector_genED_M_100_400_V_100 (
input logic signed [31:0] matrix[0:`size_minus_1(`matrix_size_1)][0:`size_minus_1(`matrix_size_2)],
input logic signed [31:0] vector[0:`size_minus_1(`vector_size)],
output logic signed [31:0] result[0:`size_minus_1(`matrix_size_2)]
);
assign result[0] = matrix[0][0] * vector[0] +matrix[1][0] * vector[1] +matrix[2][0] * vector[2] +matrix[3][0] * vector[3] +matrix[4][0] * vector[4] +matrix[5][0] * vector[5] +matrix[6][0] * vector[6] +matrix[7][0] * vector[7] +matrix[8][0] * vector[8] +matrix[9][0] * vector[9] +matrix[10][0] * vector[10] +matrix[11][0] * vector[11] +matrix[12][0] * vector[12] +matrix[13][0] * vector[13] +matrix[14][0] * vector[14] +matrix[15][0] * vector[15] +matrix[16][0] * vector[16] +matrix[17][0] * vector[17] +matrix[18][0] * vector[18] +matrix[19][0] * vector[19] +matrix[20][0] * vector[20] +matrix[21][0] * vector[21] +matrix[22][0] * vector[22] +matrix[23][0] * vector[23] +matrix[24][0] * vector[24] +matrix[25][0] * vector[25] +matrix[26][0] * vector[26] +matrix[27][0] * vector[27] +matrix[28][0] * vector[28] +matrix[29][0] * vector[29] +matrix[30][0] * vector[30] +matrix[31][0] * vector[31] +matrix[32][0] * vector[32] +matrix[33][0] * vector[33] +matrix[34][0] * vector[34] +matrix[35][0] * vector[35] +matrix[36][0] * vector[36] +matrix[37][0] * vector[37] +matrix[38][0] * vector[38] +matrix[39][0] * vector[39] +matrix[40][0] * vector[40] +matrix[41][0] * vector[41] +matrix[42][0] * vector[42] +matrix[43][0] * vector[43] +matrix[44][0] * vector[44] +matrix[45][0] * vector[45] +matrix[46][0] * vector[46] +matrix[47][0] * vector[47] +matrix[48][0] * vector[48] +matrix[49][0] * vector[49] +matrix[50][0] * vector[50] +matrix[51][0] * vector[51] +matrix[52][0] * vector[52] +matrix[53][0] * vector[53] +matrix[54][0] * vector[54] +matrix[55][0] * vector[55] +matrix[56][0] * vector[56] +matrix[57][0] * vector[57] +matrix[58][0] * vector[58] +matrix[59][0] * vector[59] +matrix[60][0] * vector[60] +matrix[61][0] * vector[61] +matrix[62][0] * vector[62] +matrix[63][0] * vector[63] +matrix[64][0] * vector[64] +matrix[65][0] * vector[65] +matrix[66][0] * vector[66] +matrix[67][0] * vector[67] +matrix[68][0] * vector[68] +matrix[69][0] * vector[69] +matrix[70][0] * vector[70] +matrix[71][0] * vector[71] +matrix[72][0] * vector[72] +matrix[73][0] * vector[73] +matrix[74][0] * vector[74] +matrix[75][0] * vector[75] +matrix[76][0] * vector[76] +matrix[77][0] * vector[77] +matrix[78][0] * vector[78] +matrix[79][0] * vector[79] +matrix[80][0] * vector[80] +matrix[81][0] * vector[81] +matrix[82][0] * vector[82] +matrix[83][0] * vector[83] +matrix[84][0] * vector[84] +matrix[85][0] * vector[85] +matrix[86][0] * vector[86] +matrix[87][0] * vector[87] +matrix[88][0] * vector[88] +matrix[89][0] * vector[89] +matrix[90][0] * vector[90] +matrix[91][0] * vector[91] +matrix[92][0] * vector[92] +matrix[93][0] * vector[93] +matrix[94][0] * vector[94] +matrix[95][0] * vector[95] +matrix[96][0] * vector[96] +matrix[97][0] * vector[97] +matrix[98][0] * vector[98] +matrix[99][0] * vector[99] +b[0];
assign result[1] = matrix[0][1] * vector[0] +matrix[1][1] * vector[1] +matrix[2][1] * vector[2] +matrix[3][1] * vector[3] +matrix[4][1] * vector[4] +matrix[5][1] * vector[5] +matrix[6][1] * vector[6] +matrix[7][1] * vector[7] +matrix[8][1] * vector[8] +matrix[9][1] * vector[9] +matrix[10][1] * vector[10] +matrix[11][1] * vector[11] +matrix[12][1] * vector[12] +matrix[13][1] * vector[13] +matrix[14][1] * vector[14] +matrix[15][1] * vector[15] +matrix[16][1] * vector[16] +matrix[17][1] * vector[17] +matrix[18][1] * vector[18] +matrix[19][1] * vector[19] +matrix[20][1] * vector[20] +matrix[21][1] * vector[21] +matrix[22][1] * vector[22] +matrix[23][1] * vector[23] +matrix[24][1] * vector[24] +matrix[25][1] * vector[25] +matrix[26][1] * vector[26] +matrix[27][1] * vector[27] +matrix[28][1] * vector[28] +matrix[29][1] * vector[29] +matrix[30][1] * vector[30] +matrix[31][1] * vector[31] +matrix[32][1] * vector[32] +matrix[33][1] * vector[33] +matrix[34][1] * vector[34] +matrix[35][1] * vector[35] +matrix[36][1] * vector[36] +matrix[37][1] * vector[37] +matrix[38][1] * vector[38] +matrix[39][1] * vector[39] +matrix[40][1] * vector[40] +matrix[41][1] * vector[41] +matrix[42][1] * vector[42] +matrix[43][1] * vector[43] +matrix[44][1] * vector[44] +matrix[45][1] * vector[45] +matrix[46][1] * vector[46] +matrix[47][1] * vector[47] +matrix[48][1] * vector[48] +matrix[49][1] * vector[49] +matrix[50][1] * vector[50] +matrix[51][1] * vector[51] +matrix[52][1] * vector[52] +matrix[53][1] * vector[53] +matrix[54][1] * vector[54] +matrix[55][1] * vector[55] +matrix[56][1] * vector[56] +matrix[57][1] * vector[57] +matrix[58][1] * vector[58] +matrix[59][1] * vector[59] +matrix[60][1] * vector[60] +matrix[61][1] * vector[61] +matrix[62][1] * vector[62] +matrix[63][1] * vector[63] +matrix[64][1] * vector[64] +matrix[65][1] * vector[65] +matrix[66][1] * vector[66] +matrix[67][1] * vector[67] +matrix[68][1] * vector[68] +matrix[69][1] * vector[69] +matrix[70][1] * vector[70] +matrix[71][1] * vector[71] +matrix[72][1] * vector[72] +matrix[73][1] * vector[73] +matrix[74][1] * vector[74] +matrix[75][1] * vector[75] +matrix[76][1] * vector[76] +matrix[77][1] * vector[77] +matrix[78][1] * vector[78] +matrix[79][1] * vector[79] +matrix[80][1] * vector[80] +matrix[81][1] * vector[81] +matrix[82][1] * vector[82] +matrix[83][1] * vector[83] +matrix[84][1] * vector[84] +matrix[85][1] * vector[85] +matrix[86][1] * vector[86] +matrix[87][1] * vector[87] +matrix[88][1] * vector[88] +matrix[89][1] * vector[89] +matrix[90][1] * vector[90] +matrix[91][1] * vector[91] +matrix[92][1] * vector[92] +matrix[93][1] * vector[93] +matrix[94][1] * vector[94] +matrix[95][1] * vector[95] +matrix[96][1] * vector[96] +matrix[97][1] * vector[97] +matrix[98][1] * vector[98] +matrix[99][1] * vector[99] +b[1];
assign result[2] = matrix[0][2] * vector[0] +matrix[1][2] * vector[1] +matrix[2][2] * vector[2] +matrix[3][2] * vector[3] +matrix[4][2] * vector[4] +matrix[5][2] * vector[5] +matrix[6][2] * vector[6] +matrix[7][2] * vector[7] +matrix[8][2] * vector[8] +matrix[9][2] * vector[9] +matrix[10][2] * vector[10] +matrix[11][2] * vector[11] +matrix[12][2] * vector[12] +matrix[13][2] * vector[13] +matrix[14][2] * vector[14] +matrix[15][2] * vector[15] +matrix[16][2] * vector[16] +matrix[17][2] * vector[17] +matrix[18][2] * vector[18] +matrix[19][2] * vector[19] +matrix[20][2] * vector[20] +matrix[21][2] * vector[21] +matrix[22][2] * vector[22] +matrix[23][2] * vector[23] +matrix[24][2] * vector[24] +matrix[25][2] * vector[25] +matrix[26][2] * vector[26] +matrix[27][2] * vector[27] +matrix[28][2] * vector[28] +matrix[29][2] * vector[29] +matrix[30][2] * vector[30] +matrix[31][2] * vector[31] +matrix[32][2] * vector[32] +matrix[33][2] * vector[33] +matrix[34][2] * vector[34] +matrix[35][2] * vector[35] +matrix[36][2] * vector[36] +matrix[37][2] * vector[37] +matrix[38][2] * vector[38] +matrix[39][2] * vector[39] +matrix[40][2] * vector[40] +matrix[41][2] * vector[41] +matrix[42][2] * vector[42] +matrix[43][2] * vector[43] +matrix[44][2] * vector[44] +matrix[45][2] * vector[45] +matrix[46][2] * vector[46] +matrix[47][2] * vector[47] +matrix[48][2] * vector[48] +matrix[49][2] * vector[49] +matrix[50][2] * vector[50] +matrix[51][2] * vector[51] +matrix[52][2] * vector[52] +matrix[53][2] * vector[53] +matrix[54][2] * vector[54] +matrix[55][2] * vector[55] +matrix[56][2] * vector[56] +matrix[57][2] * vector[57] +matrix[58][2] * vector[58] +matrix[59][2] * vector[59] +matrix[60][2] * vector[60] +matrix[61][2] * vector[61] +matrix[62][2] * vector[62] +matrix[63][2] * vector[63] +matrix[64][2] * vector[64] +matrix[65][2] * vector[65] +matrix[66][2] * vector[66] +matrix[67][2] * vector[67] +matrix[68][2] * vector[68] +matrix[69][2] * vector[69] +matrix[70][2] * vector[70] +matrix[71][2] * vector[71] +matrix[72][2] * vector[72] +matrix[73][2] * vector[73] +matrix[74][2] * vector[74] +matrix[75][2] * vector[75] +matrix[76][2] * vector[76] +matrix[77][2] * vector[77] +matrix[78][2] * vector[78] +matrix[79][2] * vector[79] +matrix[80][2] * vector[80] +matrix[81][2] * vector[81] +matrix[82][2] * vector[82] +matrix[83][2] * vector[83] +matrix[84][2] * vector[84] +matrix[85][2] * vector[85] +matrix[86][2] * vector[86] +matrix[87][2] * vector[87] +matrix[88][2] * vector[88] +matrix[89][2] * vector[89] +matrix[90][2] * vector[90] +matrix[91][2] * vector[91] +matrix[92][2] * vector[92] +matrix[93][2] * vector[93] +matrix[94][2] * vector[94] +matrix[95][2] * vector[95] +matrix[96][2] * vector[96] +matrix[97][2] * vector[97] +matrix[98][2] * vector[98] +matrix[99][2] * vector[99] +b[2];
assign result[3] = matrix[0][3] * vector[0] +matrix[1][3] * vector[1] +matrix[2][3] * vector[2] +matrix[3][3] * vector[3] +matrix[4][3] * vector[4] +matrix[5][3] * vector[5] +matrix[6][3] * vector[6] +matrix[7][3] * vector[7] +matrix[8][3] * vector[8] +matrix[9][3] * vector[9] +matrix[10][3] * vector[10] +matrix[11][3] * vector[11] +matrix[12][3] * vector[12] +matrix[13][3] * vector[13] +matrix[14][3] * vector[14] +matrix[15][3] * vector[15] +matrix[16][3] * vector[16] +matrix[17][3] * vector[17] +matrix[18][3] * vector[18] +matrix[19][3] * vector[19] +matrix[20][3] * vector[20] +matrix[21][3] * vector[21] +matrix[22][3] * vector[22] +matrix[23][3] * vector[23] +matrix[24][3] * vector[24] +matrix[25][3] * vector[25] +matrix[26][3] * vector[26] +matrix[27][3] * vector[27] +matrix[28][3] * vector[28] +matrix[29][3] * vector[29] +matrix[30][3] * vector[30] +matrix[31][3] * vector[31] +matrix[32][3] * vector[32] +matrix[33][3] * vector[33] +matrix[34][3] * vector[34] +matrix[35][3] * vector[35] +matrix[36][3] * vector[36] +matrix[37][3] * vector[37] +matrix[38][3] * vector[38] +matrix[39][3] * vector[39] +matrix[40][3] * vector[40] +matrix[41][3] * vector[41] +matrix[42][3] * vector[42] +matrix[43][3] * vector[43] +matrix[44][3] * vector[44] +matrix[45][3] * vector[45] +matrix[46][3] * vector[46] +matrix[47][3] * vector[47] +matrix[48][3] * vector[48] +matrix[49][3] * vector[49] +matrix[50][3] * vector[50] +matrix[51][3] * vector[51] +matrix[52][3] * vector[52] +matrix[53][3] * vector[53] +matrix[54][3] * vector[54] +matrix[55][3] * vector[55] +matrix[56][3] * vector[56] +matrix[57][3] * vector[57] +matrix[58][3] * vector[58] +matrix[59][3] * vector[59] +matrix[60][3] * vector[60] +matrix[61][3] * vector[61] +matrix[62][3] * vector[62] +matrix[63][3] * vector[63] +matrix[64][3] * vector[64] +matrix[65][3] * vector[65] +matrix[66][3] * vector[66] +matrix[67][3] * vector[67] +matrix[68][3] * vector[68] +matrix[69][3] * vector[69] +matrix[70][3] * vector[70] +matrix[71][3] * vector[71] +matrix[72][3] * vector[72] +matrix[73][3] * vector[73] +matrix[74][3] * vector[74] +matrix[75][3] * vector[75] +matrix[76][3] * vector[76] +matrix[77][3] * vector[77] +matrix[78][3] * vector[78] +matrix[79][3] * vector[79] +matrix[80][3] * vector[80] +matrix[81][3] * vector[81] +matrix[82][3] * vector[82] +matrix[83][3] * vector[83] +matrix[84][3] * vector[84] +matrix[85][3] * vector[85] +matrix[86][3] * vector[86] +matrix[87][3] * vector[87] +matrix[88][3] * vector[88] +matrix[89][3] * vector[89] +matrix[90][3] * vector[90] +matrix[91][3] * vector[91] +matrix[92][3] * vector[92] +matrix[93][3] * vector[93] +matrix[94][3] * vector[94] +matrix[95][3] * vector[95] +matrix[96][3] * vector[96] +matrix[97][3] * vector[97] +matrix[98][3] * vector[98] +matrix[99][3] * vector[99] +b[3];
assign result[4] = matrix[0][4] * vector[0] +matrix[1][4] * vector[1] +matrix[2][4] * vector[2] +matrix[3][4] * vector[3] +matrix[4][4] * vector[4] +matrix[5][4] * vector[5] +matrix[6][4] * vector[6] +matrix[7][4] * vector[7] +matrix[8][4] * vector[8] +matrix[9][4] * vector[9] +matrix[10][4] * vector[10] +matrix[11][4] * vector[11] +matrix[12][4] * vector[12] +matrix[13][4] * vector[13] +matrix[14][4] * vector[14] +matrix[15][4] * vector[15] +matrix[16][4] * vector[16] +matrix[17][4] * vector[17] +matrix[18][4] * vector[18] +matrix[19][4] * vector[19] +matrix[20][4] * vector[20] +matrix[21][4] * vector[21] +matrix[22][4] * vector[22] +matrix[23][4] * vector[23] +matrix[24][4] * vector[24] +matrix[25][4] * vector[25] +matrix[26][4] * vector[26] +matrix[27][4] * vector[27] +matrix[28][4] * vector[28] +matrix[29][4] * vector[29] +matrix[30][4] * vector[30] +matrix[31][4] * vector[31] +matrix[32][4] * vector[32] +matrix[33][4] * vector[33] +matrix[34][4] * vector[34] +matrix[35][4] * vector[35] +matrix[36][4] * vector[36] +matrix[37][4] * vector[37] +matrix[38][4] * vector[38] +matrix[39][4] * vector[39] +matrix[40][4] * vector[40] +matrix[41][4] * vector[41] +matrix[42][4] * vector[42] +matrix[43][4] * vector[43] +matrix[44][4] * vector[44] +matrix[45][4] * vector[45] +matrix[46][4] * vector[46] +matrix[47][4] * vector[47] +matrix[48][4] * vector[48] +matrix[49][4] * vector[49] +matrix[50][4] * vector[50] +matrix[51][4] * vector[51] +matrix[52][4] * vector[52] +matrix[53][4] * vector[53] +matrix[54][4] * vector[54] +matrix[55][4] * vector[55] +matrix[56][4] * vector[56] +matrix[57][4] * vector[57] +matrix[58][4] * vector[58] +matrix[59][4] * vector[59] +matrix[60][4] * vector[60] +matrix[61][4] * vector[61] +matrix[62][4] * vector[62] +matrix[63][4] * vector[63] +matrix[64][4] * vector[64] +matrix[65][4] * vector[65] +matrix[66][4] * vector[66] +matrix[67][4] * vector[67] +matrix[68][4] * vector[68] +matrix[69][4] * vector[69] +matrix[70][4] * vector[70] +matrix[71][4] * vector[71] +matrix[72][4] * vector[72] +matrix[73][4] * vector[73] +matrix[74][4] * vector[74] +matrix[75][4] * vector[75] +matrix[76][4] * vector[76] +matrix[77][4] * vector[77] +matrix[78][4] * vector[78] +matrix[79][4] * vector[79] +matrix[80][4] * vector[80] +matrix[81][4] * vector[81] +matrix[82][4] * vector[82] +matrix[83][4] * vector[83] +matrix[84][4] * vector[84] +matrix[85][4] * vector[85] +matrix[86][4] * vector[86] +matrix[87][4] * vector[87] +matrix[88][4] * vector[88] +matrix[89][4] * vector[89] +matrix[90][4] * vector[90] +matrix[91][4] * vector[91] +matrix[92][4] * vector[92] +matrix[93][4] * vector[93] +matrix[94][4] * vector[94] +matrix[95][4] * vector[95] +matrix[96][4] * vector[96] +matrix[97][4] * vector[97] +matrix[98][4] * vector[98] +matrix[99][4] * vector[99] +b[4];
assign result[5] = matrix[0][5] * vector[0] +matrix[1][5] * vector[1] +matrix[2][5] * vector[2] +matrix[3][5] * vector[3] +matrix[4][5] * vector[4] +matrix[5][5] * vector[5] +matrix[6][5] * vector[6] +matrix[7][5] * vector[7] +matrix[8][5] * vector[8] +matrix[9][5] * vector[9] +matrix[10][5] * vector[10] +matrix[11][5] * vector[11] +matrix[12][5] * vector[12] +matrix[13][5] * vector[13] +matrix[14][5] * vector[14] +matrix[15][5] * vector[15] +matrix[16][5] * vector[16] +matrix[17][5] * vector[17] +matrix[18][5] * vector[18] +matrix[19][5] * vector[19] +matrix[20][5] * vector[20] +matrix[21][5] * vector[21] +matrix[22][5] * vector[22] +matrix[23][5] * vector[23] +matrix[24][5] * vector[24] +matrix[25][5] * vector[25] +matrix[26][5] * vector[26] +matrix[27][5] * vector[27] +matrix[28][5] * vector[28] +matrix[29][5] * vector[29] +matrix[30][5] * vector[30] +matrix[31][5] * vector[31] +matrix[32][5] * vector[32] +matrix[33][5] * vector[33] +matrix[34][5] * vector[34] +matrix[35][5] * vector[35] +matrix[36][5] * vector[36] +matrix[37][5] * vector[37] +matrix[38][5] * vector[38] +matrix[39][5] * vector[39] +matrix[40][5] * vector[40] +matrix[41][5] * vector[41] +matrix[42][5] * vector[42] +matrix[43][5] * vector[43] +matrix[44][5] * vector[44] +matrix[45][5] * vector[45] +matrix[46][5] * vector[46] +matrix[47][5] * vector[47] +matrix[48][5] * vector[48] +matrix[49][5] * vector[49] +matrix[50][5] * vector[50] +matrix[51][5] * vector[51] +matrix[52][5] * vector[52] +matrix[53][5] * vector[53] +matrix[54][5] * vector[54] +matrix[55][5] * vector[55] +matrix[56][5] * vector[56] +matrix[57][5] * vector[57] +matrix[58][5] * vector[58] +matrix[59][5] * vector[59] +matrix[60][5] * vector[60] +matrix[61][5] * vector[61] +matrix[62][5] * vector[62] +matrix[63][5] * vector[63] +matrix[64][5] * vector[64] +matrix[65][5] * vector[65] +matrix[66][5] * vector[66] +matrix[67][5] * vector[67] +matrix[68][5] * vector[68] +matrix[69][5] * vector[69] +matrix[70][5] * vector[70] +matrix[71][5] * vector[71] +matrix[72][5] * vector[72] +matrix[73][5] * vector[73] +matrix[74][5] * vector[74] +matrix[75][5] * vector[75] +matrix[76][5] * vector[76] +matrix[77][5] * vector[77] +matrix[78][5] * vector[78] +matrix[79][5] * vector[79] +matrix[80][5] * vector[80] +matrix[81][5] * vector[81] +matrix[82][5] * vector[82] +matrix[83][5] * vector[83] +matrix[84][5] * vector[84] +matrix[85][5] * vector[85] +matrix[86][5] * vector[86] +matrix[87][5] * vector[87] +matrix[88][5] * vector[88] +matrix[89][5] * vector[89] +matrix[90][5] * vector[90] +matrix[91][5] * vector[91] +matrix[92][5] * vector[92] +matrix[93][5] * vector[93] +matrix[94][5] * vector[94] +matrix[95][5] * vector[95] +matrix[96][5] * vector[96] +matrix[97][5] * vector[97] +matrix[98][5] * vector[98] +matrix[99][5] * vector[99] +b[5];
assign result[6] = matrix[0][6] * vector[0] +matrix[1][6] * vector[1] +matrix[2][6] * vector[2] +matrix[3][6] * vector[3] +matrix[4][6] * vector[4] +matrix[5][6] * vector[5] +matrix[6][6] * vector[6] +matrix[7][6] * vector[7] +matrix[8][6] * vector[8] +matrix[9][6] * vector[9] +matrix[10][6] * vector[10] +matrix[11][6] * vector[11] +matrix[12][6] * vector[12] +matrix[13][6] * vector[13] +matrix[14][6] * vector[14] +matrix[15][6] * vector[15] +matrix[16][6] * vector[16] +matrix[17][6] * vector[17] +matrix[18][6] * vector[18] +matrix[19][6] * vector[19] +matrix[20][6] * vector[20] +matrix[21][6] * vector[21] +matrix[22][6] * vector[22] +matrix[23][6] * vector[23] +matrix[24][6] * vector[24] +matrix[25][6] * vector[25] +matrix[26][6] * vector[26] +matrix[27][6] * vector[27] +matrix[28][6] * vector[28] +matrix[29][6] * vector[29] +matrix[30][6] * vector[30] +matrix[31][6] * vector[31] +matrix[32][6] * vector[32] +matrix[33][6] * vector[33] +matrix[34][6] * vector[34] +matrix[35][6] * vector[35] +matrix[36][6] * vector[36] +matrix[37][6] * vector[37] +matrix[38][6] * vector[38] +matrix[39][6] * vector[39] +matrix[40][6] * vector[40] +matrix[41][6] * vector[41] +matrix[42][6] * vector[42] +matrix[43][6] * vector[43] +matrix[44][6] * vector[44] +matrix[45][6] * vector[45] +matrix[46][6] * vector[46] +matrix[47][6] * vector[47] +matrix[48][6] * vector[48] +matrix[49][6] * vector[49] +matrix[50][6] * vector[50] +matrix[51][6] * vector[51] +matrix[52][6] * vector[52] +matrix[53][6] * vector[53] +matrix[54][6] * vector[54] +matrix[55][6] * vector[55] +matrix[56][6] * vector[56] +matrix[57][6] * vector[57] +matrix[58][6] * vector[58] +matrix[59][6] * vector[59] +matrix[60][6] * vector[60] +matrix[61][6] * vector[61] +matrix[62][6] * vector[62] +matrix[63][6] * vector[63] +matrix[64][6] * vector[64] +matrix[65][6] * vector[65] +matrix[66][6] * vector[66] +matrix[67][6] * vector[67] +matrix[68][6] * vector[68] +matrix[69][6] * vector[69] +matrix[70][6] * vector[70] +matrix[71][6] * vector[71] +matrix[72][6] * vector[72] +matrix[73][6] * vector[73] +matrix[74][6] * vector[74] +matrix[75][6] * vector[75] +matrix[76][6] * vector[76] +matrix[77][6] * vector[77] +matrix[78][6] * vector[78] +matrix[79][6] * vector[79] +matrix[80][6] * vector[80] +matrix[81][6] * vector[81] +matrix[82][6] * vector[82] +matrix[83][6] * vector[83] +matrix[84][6] * vector[84] +matrix[85][6] * vector[85] +matrix[86][6] * vector[86] +matrix[87][6] * vector[87] +matrix[88][6] * vector[88] +matrix[89][6] * vector[89] +matrix[90][6] * vector[90] +matrix[91][6] * vector[91] +matrix[92][6] * vector[92] +matrix[93][6] * vector[93] +matrix[94][6] * vector[94] +matrix[95][6] * vector[95] +matrix[96][6] * vector[96] +matrix[97][6] * vector[97] +matrix[98][6] * vector[98] +matrix[99][6] * vector[99] +b[6];
assign result[7] = matrix[0][7] * vector[0] +matrix[1][7] * vector[1] +matrix[2][7] * vector[2] +matrix[3][7] * vector[3] +matrix[4][7] * vector[4] +matrix[5][7] * vector[5] +matrix[6][7] * vector[6] +matrix[7][7] * vector[7] +matrix[8][7] * vector[8] +matrix[9][7] * vector[9] +matrix[10][7] * vector[10] +matrix[11][7] * vector[11] +matrix[12][7] * vector[12] +matrix[13][7] * vector[13] +matrix[14][7] * vector[14] +matrix[15][7] * vector[15] +matrix[16][7] * vector[16] +matrix[17][7] * vector[17] +matrix[18][7] * vector[18] +matrix[19][7] * vector[19] +matrix[20][7] * vector[20] +matrix[21][7] * vector[21] +matrix[22][7] * vector[22] +matrix[23][7] * vector[23] +matrix[24][7] * vector[24] +matrix[25][7] * vector[25] +matrix[26][7] * vector[26] +matrix[27][7] * vector[27] +matrix[28][7] * vector[28] +matrix[29][7] * vector[29] +matrix[30][7] * vector[30] +matrix[31][7] * vector[31] +matrix[32][7] * vector[32] +matrix[33][7] * vector[33] +matrix[34][7] * vector[34] +matrix[35][7] * vector[35] +matrix[36][7] * vector[36] +matrix[37][7] * vector[37] +matrix[38][7] * vector[38] +matrix[39][7] * vector[39] +matrix[40][7] * vector[40] +matrix[41][7] * vector[41] +matrix[42][7] * vector[42] +matrix[43][7] * vector[43] +matrix[44][7] * vector[44] +matrix[45][7] * vector[45] +matrix[46][7] * vector[46] +matrix[47][7] * vector[47] +matrix[48][7] * vector[48] +matrix[49][7] * vector[49] +matrix[50][7] * vector[50] +matrix[51][7] * vector[51] +matrix[52][7] * vector[52] +matrix[53][7] * vector[53] +matrix[54][7] * vector[54] +matrix[55][7] * vector[55] +matrix[56][7] * vector[56] +matrix[57][7] * vector[57] +matrix[58][7] * vector[58] +matrix[59][7] * vector[59] +matrix[60][7] * vector[60] +matrix[61][7] * vector[61] +matrix[62][7] * vector[62] +matrix[63][7] * vector[63] +matrix[64][7] * vector[64] +matrix[65][7] * vector[65] +matrix[66][7] * vector[66] +matrix[67][7] * vector[67] +matrix[68][7] * vector[68] +matrix[69][7] * vector[69] +matrix[70][7] * vector[70] +matrix[71][7] * vector[71] +matrix[72][7] * vector[72] +matrix[73][7] * vector[73] +matrix[74][7] * vector[74] +matrix[75][7] * vector[75] +matrix[76][7] * vector[76] +matrix[77][7] * vector[77] +matrix[78][7] * vector[78] +matrix[79][7] * vector[79] +matrix[80][7] * vector[80] +matrix[81][7] * vector[81] +matrix[82][7] * vector[82] +matrix[83][7] * vector[83] +matrix[84][7] * vector[84] +matrix[85][7] * vector[85] +matrix[86][7] * vector[86] +matrix[87][7] * vector[87] +matrix[88][7] * vector[88] +matrix[89][7] * vector[89] +matrix[90][7] * vector[90] +matrix[91][7] * vector[91] +matrix[92][7] * vector[92] +matrix[93][7] * vector[93] +matrix[94][7] * vector[94] +matrix[95][7] * vector[95] +matrix[96][7] * vector[96] +matrix[97][7] * vector[97] +matrix[98][7] * vector[98] +matrix[99][7] * vector[99] +b[7];
assign result[8] = matrix[0][8] * vector[0] +matrix[1][8] * vector[1] +matrix[2][8] * vector[2] +matrix[3][8] * vector[3] +matrix[4][8] * vector[4] +matrix[5][8] * vector[5] +matrix[6][8] * vector[6] +matrix[7][8] * vector[7] +matrix[8][8] * vector[8] +matrix[9][8] * vector[9] +matrix[10][8] * vector[10] +matrix[11][8] * vector[11] +matrix[12][8] * vector[12] +matrix[13][8] * vector[13] +matrix[14][8] * vector[14] +matrix[15][8] * vector[15] +matrix[16][8] * vector[16] +matrix[17][8] * vector[17] +matrix[18][8] * vector[18] +matrix[19][8] * vector[19] +matrix[20][8] * vector[20] +matrix[21][8] * vector[21] +matrix[22][8] * vector[22] +matrix[23][8] * vector[23] +matrix[24][8] * vector[24] +matrix[25][8] * vector[25] +matrix[26][8] * vector[26] +matrix[27][8] * vector[27] +matrix[28][8] * vector[28] +matrix[29][8] * vector[29] +matrix[30][8] * vector[30] +matrix[31][8] * vector[31] +matrix[32][8] * vector[32] +matrix[33][8] * vector[33] +matrix[34][8] * vector[34] +matrix[35][8] * vector[35] +matrix[36][8] * vector[36] +matrix[37][8] * vector[37] +matrix[38][8] * vector[38] +matrix[39][8] * vector[39] +matrix[40][8] * vector[40] +matrix[41][8] * vector[41] +matrix[42][8] * vector[42] +matrix[43][8] * vector[43] +matrix[44][8] * vector[44] +matrix[45][8] * vector[45] +matrix[46][8] * vector[46] +matrix[47][8] * vector[47] +matrix[48][8] * vector[48] +matrix[49][8] * vector[49] +matrix[50][8] * vector[50] +matrix[51][8] * vector[51] +matrix[52][8] * vector[52] +matrix[53][8] * vector[53] +matrix[54][8] * vector[54] +matrix[55][8] * vector[55] +matrix[56][8] * vector[56] +matrix[57][8] * vector[57] +matrix[58][8] * vector[58] +matrix[59][8] * vector[59] +matrix[60][8] * vector[60] +matrix[61][8] * vector[61] +matrix[62][8] * vector[62] +matrix[63][8] * vector[63] +matrix[64][8] * vector[64] +matrix[65][8] * vector[65] +matrix[66][8] * vector[66] +matrix[67][8] * vector[67] +matrix[68][8] * vector[68] +matrix[69][8] * vector[69] +matrix[70][8] * vector[70] +matrix[71][8] * vector[71] +matrix[72][8] * vector[72] +matrix[73][8] * vector[73] +matrix[74][8] * vector[74] +matrix[75][8] * vector[75] +matrix[76][8] * vector[76] +matrix[77][8] * vector[77] +matrix[78][8] * vector[78] +matrix[79][8] * vector[79] +matrix[80][8] * vector[80] +matrix[81][8] * vector[81] +matrix[82][8] * vector[82] +matrix[83][8] * vector[83] +matrix[84][8] * vector[84] +matrix[85][8] * vector[85] +matrix[86][8] * vector[86] +matrix[87][8] * vector[87] +matrix[88][8] * vector[88] +matrix[89][8] * vector[89] +matrix[90][8] * vector[90] +matrix[91][8] * vector[91] +matrix[92][8] * vector[92] +matrix[93][8] * vector[93] +matrix[94][8] * vector[94] +matrix[95][8] * vector[95] +matrix[96][8] * vector[96] +matrix[97][8] * vector[97] +matrix[98][8] * vector[98] +matrix[99][8] * vector[99] +b[8];
assign result[9] = matrix[0][9] * vector[0] +matrix[1][9] * vector[1] +matrix[2][9] * vector[2] +matrix[3][9] * vector[3] +matrix[4][9] * vector[4] +matrix[5][9] * vector[5] +matrix[6][9] * vector[6] +matrix[7][9] * vector[7] +matrix[8][9] * vector[8] +matrix[9][9] * vector[9] +matrix[10][9] * vector[10] +matrix[11][9] * vector[11] +matrix[12][9] * vector[12] +matrix[13][9] * vector[13] +matrix[14][9] * vector[14] +matrix[15][9] * vector[15] +matrix[16][9] * vector[16] +matrix[17][9] * vector[17] +matrix[18][9] * vector[18] +matrix[19][9] * vector[19] +matrix[20][9] * vector[20] +matrix[21][9] * vector[21] +matrix[22][9] * vector[22] +matrix[23][9] * vector[23] +matrix[24][9] * vector[24] +matrix[25][9] * vector[25] +matrix[26][9] * vector[26] +matrix[27][9] * vector[27] +matrix[28][9] * vector[28] +matrix[29][9] * vector[29] +matrix[30][9] * vector[30] +matrix[31][9] * vector[31] +matrix[32][9] * vector[32] +matrix[33][9] * vector[33] +matrix[34][9] * vector[34] +matrix[35][9] * vector[35] +matrix[36][9] * vector[36] +matrix[37][9] * vector[37] +matrix[38][9] * vector[38] +matrix[39][9] * vector[39] +matrix[40][9] * vector[40] +matrix[41][9] * vector[41] +matrix[42][9] * vector[42] +matrix[43][9] * vector[43] +matrix[44][9] * vector[44] +matrix[45][9] * vector[45] +matrix[46][9] * vector[46] +matrix[47][9] * vector[47] +matrix[48][9] * vector[48] +matrix[49][9] * vector[49] +matrix[50][9] * vector[50] +matrix[51][9] * vector[51] +matrix[52][9] * vector[52] +matrix[53][9] * vector[53] +matrix[54][9] * vector[54] +matrix[55][9] * vector[55] +matrix[56][9] * vector[56] +matrix[57][9] * vector[57] +matrix[58][9] * vector[58] +matrix[59][9] * vector[59] +matrix[60][9] * vector[60] +matrix[61][9] * vector[61] +matrix[62][9] * vector[62] +matrix[63][9] * vector[63] +matrix[64][9] * vector[64] +matrix[65][9] * vector[65] +matrix[66][9] * vector[66] +matrix[67][9] * vector[67] +matrix[68][9] * vector[68] +matrix[69][9] * vector[69] +matrix[70][9] * vector[70] +matrix[71][9] * vector[71] +matrix[72][9] * vector[72] +matrix[73][9] * vector[73] +matrix[74][9] * vector[74] +matrix[75][9] * vector[75] +matrix[76][9] * vector[76] +matrix[77][9] * vector[77] +matrix[78][9] * vector[78] +matrix[79][9] * vector[79] +matrix[80][9] * vector[80] +matrix[81][9] * vector[81] +matrix[82][9] * vector[82] +matrix[83][9] * vector[83] +matrix[84][9] * vector[84] +matrix[85][9] * vector[85] +matrix[86][9] * vector[86] +matrix[87][9] * vector[87] +matrix[88][9] * vector[88] +matrix[89][9] * vector[89] +matrix[90][9] * vector[90] +matrix[91][9] * vector[91] +matrix[92][9] * vector[92] +matrix[93][9] * vector[93] +matrix[94][9] * vector[94] +matrix[95][9] * vector[95] +matrix[96][9] * vector[96] +matrix[97][9] * vector[97] +matrix[98][9] * vector[98] +matrix[99][9] * vector[99] +b[9];
assign result[10] = matrix[0][10] * vector[0] +matrix[1][10] * vector[1] +matrix[2][10] * vector[2] +matrix[3][10] * vector[3] +matrix[4][10] * vector[4] +matrix[5][10] * vector[5] +matrix[6][10] * vector[6] +matrix[7][10] * vector[7] +matrix[8][10] * vector[8] +matrix[9][10] * vector[9] +matrix[10][10] * vector[10] +matrix[11][10] * vector[11] +matrix[12][10] * vector[12] +matrix[13][10] * vector[13] +matrix[14][10] * vector[14] +matrix[15][10] * vector[15] +matrix[16][10] * vector[16] +matrix[17][10] * vector[17] +matrix[18][10] * vector[18] +matrix[19][10] * vector[19] +matrix[20][10] * vector[20] +matrix[21][10] * vector[21] +matrix[22][10] * vector[22] +matrix[23][10] * vector[23] +matrix[24][10] * vector[24] +matrix[25][10] * vector[25] +matrix[26][10] * vector[26] +matrix[27][10] * vector[27] +matrix[28][10] * vector[28] +matrix[29][10] * vector[29] +matrix[30][10] * vector[30] +matrix[31][10] * vector[31] +matrix[32][10] * vector[32] +matrix[33][10] * vector[33] +matrix[34][10] * vector[34] +matrix[35][10] * vector[35] +matrix[36][10] * vector[36] +matrix[37][10] * vector[37] +matrix[38][10] * vector[38] +matrix[39][10] * vector[39] +matrix[40][10] * vector[40] +matrix[41][10] * vector[41] +matrix[42][10] * vector[42] +matrix[43][10] * vector[43] +matrix[44][10] * vector[44] +matrix[45][10] * vector[45] +matrix[46][10] * vector[46] +matrix[47][10] * vector[47] +matrix[48][10] * vector[48] +matrix[49][10] * vector[49] +matrix[50][10] * vector[50] +matrix[51][10] * vector[51] +matrix[52][10] * vector[52] +matrix[53][10] * vector[53] +matrix[54][10] * vector[54] +matrix[55][10] * vector[55] +matrix[56][10] * vector[56] +matrix[57][10] * vector[57] +matrix[58][10] * vector[58] +matrix[59][10] * vector[59] +matrix[60][10] * vector[60] +matrix[61][10] * vector[61] +matrix[62][10] * vector[62] +matrix[63][10] * vector[63] +matrix[64][10] * vector[64] +matrix[65][10] * vector[65] +matrix[66][10] * vector[66] +matrix[67][10] * vector[67] +matrix[68][10] * vector[68] +matrix[69][10] * vector[69] +matrix[70][10] * vector[70] +matrix[71][10] * vector[71] +matrix[72][10] * vector[72] +matrix[73][10] * vector[73] +matrix[74][10] * vector[74] +matrix[75][10] * vector[75] +matrix[76][10] * vector[76] +matrix[77][10] * vector[77] +matrix[78][10] * vector[78] +matrix[79][10] * vector[79] +matrix[80][10] * vector[80] +matrix[81][10] * vector[81] +matrix[82][10] * vector[82] +matrix[83][10] * vector[83] +matrix[84][10] * vector[84] +matrix[85][10] * vector[85] +matrix[86][10] * vector[86] +matrix[87][10] * vector[87] +matrix[88][10] * vector[88] +matrix[89][10] * vector[89] +matrix[90][10] * vector[90] +matrix[91][10] * vector[91] +matrix[92][10] * vector[92] +matrix[93][10] * vector[93] +matrix[94][10] * vector[94] +matrix[95][10] * vector[95] +matrix[96][10] * vector[96] +matrix[97][10] * vector[97] +matrix[98][10] * vector[98] +matrix[99][10] * vector[99] +b[10];
assign result[11] = matrix[0][11] * vector[0] +matrix[1][11] * vector[1] +matrix[2][11] * vector[2] +matrix[3][11] * vector[3] +matrix[4][11] * vector[4] +matrix[5][11] * vector[5] +matrix[6][11] * vector[6] +matrix[7][11] * vector[7] +matrix[8][11] * vector[8] +matrix[9][11] * vector[9] +matrix[10][11] * vector[10] +matrix[11][11] * vector[11] +matrix[12][11] * vector[12] +matrix[13][11] * vector[13] +matrix[14][11] * vector[14] +matrix[15][11] * vector[15] +matrix[16][11] * vector[16] +matrix[17][11] * vector[17] +matrix[18][11] * vector[18] +matrix[19][11] * vector[19] +matrix[20][11] * vector[20] +matrix[21][11] * vector[21] +matrix[22][11] * vector[22] +matrix[23][11] * vector[23] +matrix[24][11] * vector[24] +matrix[25][11] * vector[25] +matrix[26][11] * vector[26] +matrix[27][11] * vector[27] +matrix[28][11] * vector[28] +matrix[29][11] * vector[29] +matrix[30][11] * vector[30] +matrix[31][11] * vector[31] +matrix[32][11] * vector[32] +matrix[33][11] * vector[33] +matrix[34][11] * vector[34] +matrix[35][11] * vector[35] +matrix[36][11] * vector[36] +matrix[37][11] * vector[37] +matrix[38][11] * vector[38] +matrix[39][11] * vector[39] +matrix[40][11] * vector[40] +matrix[41][11] * vector[41] +matrix[42][11] * vector[42] +matrix[43][11] * vector[43] +matrix[44][11] * vector[44] +matrix[45][11] * vector[45] +matrix[46][11] * vector[46] +matrix[47][11] * vector[47] +matrix[48][11] * vector[48] +matrix[49][11] * vector[49] +matrix[50][11] * vector[50] +matrix[51][11] * vector[51] +matrix[52][11] * vector[52] +matrix[53][11] * vector[53] +matrix[54][11] * vector[54] +matrix[55][11] * vector[55] +matrix[56][11] * vector[56] +matrix[57][11] * vector[57] +matrix[58][11] * vector[58] +matrix[59][11] * vector[59] +matrix[60][11] * vector[60] +matrix[61][11] * vector[61] +matrix[62][11] * vector[62] +matrix[63][11] * vector[63] +matrix[64][11] * vector[64] +matrix[65][11] * vector[65] +matrix[66][11] * vector[66] +matrix[67][11] * vector[67] +matrix[68][11] * vector[68] +matrix[69][11] * vector[69] +matrix[70][11] * vector[70] +matrix[71][11] * vector[71] +matrix[72][11] * vector[72] +matrix[73][11] * vector[73] +matrix[74][11] * vector[74] +matrix[75][11] * vector[75] +matrix[76][11] * vector[76] +matrix[77][11] * vector[77] +matrix[78][11] * vector[78] +matrix[79][11] * vector[79] +matrix[80][11] * vector[80] +matrix[81][11] * vector[81] +matrix[82][11] * vector[82] +matrix[83][11] * vector[83] +matrix[84][11] * vector[84] +matrix[85][11] * vector[85] +matrix[86][11] * vector[86] +matrix[87][11] * vector[87] +matrix[88][11] * vector[88] +matrix[89][11] * vector[89] +matrix[90][11] * vector[90] +matrix[91][11] * vector[91] +matrix[92][11] * vector[92] +matrix[93][11] * vector[93] +matrix[94][11] * vector[94] +matrix[95][11] * vector[95] +matrix[96][11] * vector[96] +matrix[97][11] * vector[97] +matrix[98][11] * vector[98] +matrix[99][11] * vector[99] +b[11];
assign result[12] = matrix[0][12] * vector[0] +matrix[1][12] * vector[1] +matrix[2][12] * vector[2] +matrix[3][12] * vector[3] +matrix[4][12] * vector[4] +matrix[5][12] * vector[5] +matrix[6][12] * vector[6] +matrix[7][12] * vector[7] +matrix[8][12] * vector[8] +matrix[9][12] * vector[9] +matrix[10][12] * vector[10] +matrix[11][12] * vector[11] +matrix[12][12] * vector[12] +matrix[13][12] * vector[13] +matrix[14][12] * vector[14] +matrix[15][12] * vector[15] +matrix[16][12] * vector[16] +matrix[17][12] * vector[17] +matrix[18][12] * vector[18] +matrix[19][12] * vector[19] +matrix[20][12] * vector[20] +matrix[21][12] * vector[21] +matrix[22][12] * vector[22] +matrix[23][12] * vector[23] +matrix[24][12] * vector[24] +matrix[25][12] * vector[25] +matrix[26][12] * vector[26] +matrix[27][12] * vector[27] +matrix[28][12] * vector[28] +matrix[29][12] * vector[29] +matrix[30][12] * vector[30] +matrix[31][12] * vector[31] +matrix[32][12] * vector[32] +matrix[33][12] * vector[33] +matrix[34][12] * vector[34] +matrix[35][12] * vector[35] +matrix[36][12] * vector[36] +matrix[37][12] * vector[37] +matrix[38][12] * vector[38] +matrix[39][12] * vector[39] +matrix[40][12] * vector[40] +matrix[41][12] * vector[41] +matrix[42][12] * vector[42] +matrix[43][12] * vector[43] +matrix[44][12] * vector[44] +matrix[45][12] * vector[45] +matrix[46][12] * vector[46] +matrix[47][12] * vector[47] +matrix[48][12] * vector[48] +matrix[49][12] * vector[49] +matrix[50][12] * vector[50] +matrix[51][12] * vector[51] +matrix[52][12] * vector[52] +matrix[53][12] * vector[53] +matrix[54][12] * vector[54] +matrix[55][12] * vector[55] +matrix[56][12] * vector[56] +matrix[57][12] * vector[57] +matrix[58][12] * vector[58] +matrix[59][12] * vector[59] +matrix[60][12] * vector[60] +matrix[61][12] * vector[61] +matrix[62][12] * vector[62] +matrix[63][12] * vector[63] +matrix[64][12] * vector[64] +matrix[65][12] * vector[65] +matrix[66][12] * vector[66] +matrix[67][12] * vector[67] +matrix[68][12] * vector[68] +matrix[69][12] * vector[69] +matrix[70][12] * vector[70] +matrix[71][12] * vector[71] +matrix[72][12] * vector[72] +matrix[73][12] * vector[73] +matrix[74][12] * vector[74] +matrix[75][12] * vector[75] +matrix[76][12] * vector[76] +matrix[77][12] * vector[77] +matrix[78][12] * vector[78] +matrix[79][12] * vector[79] +matrix[80][12] * vector[80] +matrix[81][12] * vector[81] +matrix[82][12] * vector[82] +matrix[83][12] * vector[83] +matrix[84][12] * vector[84] +matrix[85][12] * vector[85] +matrix[86][12] * vector[86] +matrix[87][12] * vector[87] +matrix[88][12] * vector[88] +matrix[89][12] * vector[89] +matrix[90][12] * vector[90] +matrix[91][12] * vector[91] +matrix[92][12] * vector[92] +matrix[93][12] * vector[93] +matrix[94][12] * vector[94] +matrix[95][12] * vector[95] +matrix[96][12] * vector[96] +matrix[97][12] * vector[97] +matrix[98][12] * vector[98] +matrix[99][12] * vector[99] +b[12];
assign result[13] = matrix[0][13] * vector[0] +matrix[1][13] * vector[1] +matrix[2][13] * vector[2] +matrix[3][13] * vector[3] +matrix[4][13] * vector[4] +matrix[5][13] * vector[5] +matrix[6][13] * vector[6] +matrix[7][13] * vector[7] +matrix[8][13] * vector[8] +matrix[9][13] * vector[9] +matrix[10][13] * vector[10] +matrix[11][13] * vector[11] +matrix[12][13] * vector[12] +matrix[13][13] * vector[13] +matrix[14][13] * vector[14] +matrix[15][13] * vector[15] +matrix[16][13] * vector[16] +matrix[17][13] * vector[17] +matrix[18][13] * vector[18] +matrix[19][13] * vector[19] +matrix[20][13] * vector[20] +matrix[21][13] * vector[21] +matrix[22][13] * vector[22] +matrix[23][13] * vector[23] +matrix[24][13] * vector[24] +matrix[25][13] * vector[25] +matrix[26][13] * vector[26] +matrix[27][13] * vector[27] +matrix[28][13] * vector[28] +matrix[29][13] * vector[29] +matrix[30][13] * vector[30] +matrix[31][13] * vector[31] +matrix[32][13] * vector[32] +matrix[33][13] * vector[33] +matrix[34][13] * vector[34] +matrix[35][13] * vector[35] +matrix[36][13] * vector[36] +matrix[37][13] * vector[37] +matrix[38][13] * vector[38] +matrix[39][13] * vector[39] +matrix[40][13] * vector[40] +matrix[41][13] * vector[41] +matrix[42][13] * vector[42] +matrix[43][13] * vector[43] +matrix[44][13] * vector[44] +matrix[45][13] * vector[45] +matrix[46][13] * vector[46] +matrix[47][13] * vector[47] +matrix[48][13] * vector[48] +matrix[49][13] * vector[49] +matrix[50][13] * vector[50] +matrix[51][13] * vector[51] +matrix[52][13] * vector[52] +matrix[53][13] * vector[53] +matrix[54][13] * vector[54] +matrix[55][13] * vector[55] +matrix[56][13] * vector[56] +matrix[57][13] * vector[57] +matrix[58][13] * vector[58] +matrix[59][13] * vector[59] +matrix[60][13] * vector[60] +matrix[61][13] * vector[61] +matrix[62][13] * vector[62] +matrix[63][13] * vector[63] +matrix[64][13] * vector[64] +matrix[65][13] * vector[65] +matrix[66][13] * vector[66] +matrix[67][13] * vector[67] +matrix[68][13] * vector[68] +matrix[69][13] * vector[69] +matrix[70][13] * vector[70] +matrix[71][13] * vector[71] +matrix[72][13] * vector[72] +matrix[73][13] * vector[73] +matrix[74][13] * vector[74] +matrix[75][13] * vector[75] +matrix[76][13] * vector[76] +matrix[77][13] * vector[77] +matrix[78][13] * vector[78] +matrix[79][13] * vector[79] +matrix[80][13] * vector[80] +matrix[81][13] * vector[81] +matrix[82][13] * vector[82] +matrix[83][13] * vector[83] +matrix[84][13] * vector[84] +matrix[85][13] * vector[85] +matrix[86][13] * vector[86] +matrix[87][13] * vector[87] +matrix[88][13] * vector[88] +matrix[89][13] * vector[89] +matrix[90][13] * vector[90] +matrix[91][13] * vector[91] +matrix[92][13] * vector[92] +matrix[93][13] * vector[93] +matrix[94][13] * vector[94] +matrix[95][13] * vector[95] +matrix[96][13] * vector[96] +matrix[97][13] * vector[97] +matrix[98][13] * vector[98] +matrix[99][13] * vector[99] +b[13];
assign result[14] = matrix[0][14] * vector[0] +matrix[1][14] * vector[1] +matrix[2][14] * vector[2] +matrix[3][14] * vector[3] +matrix[4][14] * vector[4] +matrix[5][14] * vector[5] +matrix[6][14] * vector[6] +matrix[7][14] * vector[7] +matrix[8][14] * vector[8] +matrix[9][14] * vector[9] +matrix[10][14] * vector[10] +matrix[11][14] * vector[11] +matrix[12][14] * vector[12] +matrix[13][14] * vector[13] +matrix[14][14] * vector[14] +matrix[15][14] * vector[15] +matrix[16][14] * vector[16] +matrix[17][14] * vector[17] +matrix[18][14] * vector[18] +matrix[19][14] * vector[19] +matrix[20][14] * vector[20] +matrix[21][14] * vector[21] +matrix[22][14] * vector[22] +matrix[23][14] * vector[23] +matrix[24][14] * vector[24] +matrix[25][14] * vector[25] +matrix[26][14] * vector[26] +matrix[27][14] * vector[27] +matrix[28][14] * vector[28] +matrix[29][14] * vector[29] +matrix[30][14] * vector[30] +matrix[31][14] * vector[31] +matrix[32][14] * vector[32] +matrix[33][14] * vector[33] +matrix[34][14] * vector[34] +matrix[35][14] * vector[35] +matrix[36][14] * vector[36] +matrix[37][14] * vector[37] +matrix[38][14] * vector[38] +matrix[39][14] * vector[39] +matrix[40][14] * vector[40] +matrix[41][14] * vector[41] +matrix[42][14] * vector[42] +matrix[43][14] * vector[43] +matrix[44][14] * vector[44] +matrix[45][14] * vector[45] +matrix[46][14] * vector[46] +matrix[47][14] * vector[47] +matrix[48][14] * vector[48] +matrix[49][14] * vector[49] +matrix[50][14] * vector[50] +matrix[51][14] * vector[51] +matrix[52][14] * vector[52] +matrix[53][14] * vector[53] +matrix[54][14] * vector[54] +matrix[55][14] * vector[55] +matrix[56][14] * vector[56] +matrix[57][14] * vector[57] +matrix[58][14] * vector[58] +matrix[59][14] * vector[59] +matrix[60][14] * vector[60] +matrix[61][14] * vector[61] +matrix[62][14] * vector[62] +matrix[63][14] * vector[63] +matrix[64][14] * vector[64] +matrix[65][14] * vector[65] +matrix[66][14] * vector[66] +matrix[67][14] * vector[67] +matrix[68][14] * vector[68] +matrix[69][14] * vector[69] +matrix[70][14] * vector[70] +matrix[71][14] * vector[71] +matrix[72][14] * vector[72] +matrix[73][14] * vector[73] +matrix[74][14] * vector[74] +matrix[75][14] * vector[75] +matrix[76][14] * vector[76] +matrix[77][14] * vector[77] +matrix[78][14] * vector[78] +matrix[79][14] * vector[79] +matrix[80][14] * vector[80] +matrix[81][14] * vector[81] +matrix[82][14] * vector[82] +matrix[83][14] * vector[83] +matrix[84][14] * vector[84] +matrix[85][14] * vector[85] +matrix[86][14] * vector[86] +matrix[87][14] * vector[87] +matrix[88][14] * vector[88] +matrix[89][14] * vector[89] +matrix[90][14] * vector[90] +matrix[91][14] * vector[91] +matrix[92][14] * vector[92] +matrix[93][14] * vector[93] +matrix[94][14] * vector[94] +matrix[95][14] * vector[95] +matrix[96][14] * vector[96] +matrix[97][14] * vector[97] +matrix[98][14] * vector[98] +matrix[99][14] * vector[99] +b[14];
assign result[15] = matrix[0][15] * vector[0] +matrix[1][15] * vector[1] +matrix[2][15] * vector[2] +matrix[3][15] * vector[3] +matrix[4][15] * vector[4] +matrix[5][15] * vector[5] +matrix[6][15] * vector[6] +matrix[7][15] * vector[7] +matrix[8][15] * vector[8] +matrix[9][15] * vector[9] +matrix[10][15] * vector[10] +matrix[11][15] * vector[11] +matrix[12][15] * vector[12] +matrix[13][15] * vector[13] +matrix[14][15] * vector[14] +matrix[15][15] * vector[15] +matrix[16][15] * vector[16] +matrix[17][15] * vector[17] +matrix[18][15] * vector[18] +matrix[19][15] * vector[19] +matrix[20][15] * vector[20] +matrix[21][15] * vector[21] +matrix[22][15] * vector[22] +matrix[23][15] * vector[23] +matrix[24][15] * vector[24] +matrix[25][15] * vector[25] +matrix[26][15] * vector[26] +matrix[27][15] * vector[27] +matrix[28][15] * vector[28] +matrix[29][15] * vector[29] +matrix[30][15] * vector[30] +matrix[31][15] * vector[31] +matrix[32][15] * vector[32] +matrix[33][15] * vector[33] +matrix[34][15] * vector[34] +matrix[35][15] * vector[35] +matrix[36][15] * vector[36] +matrix[37][15] * vector[37] +matrix[38][15] * vector[38] +matrix[39][15] * vector[39] +matrix[40][15] * vector[40] +matrix[41][15] * vector[41] +matrix[42][15] * vector[42] +matrix[43][15] * vector[43] +matrix[44][15] * vector[44] +matrix[45][15] * vector[45] +matrix[46][15] * vector[46] +matrix[47][15] * vector[47] +matrix[48][15] * vector[48] +matrix[49][15] * vector[49] +matrix[50][15] * vector[50] +matrix[51][15] * vector[51] +matrix[52][15] * vector[52] +matrix[53][15] * vector[53] +matrix[54][15] * vector[54] +matrix[55][15] * vector[55] +matrix[56][15] * vector[56] +matrix[57][15] * vector[57] +matrix[58][15] * vector[58] +matrix[59][15] * vector[59] +matrix[60][15] * vector[60] +matrix[61][15] * vector[61] +matrix[62][15] * vector[62] +matrix[63][15] * vector[63] +matrix[64][15] * vector[64] +matrix[65][15] * vector[65] +matrix[66][15] * vector[66] +matrix[67][15] * vector[67] +matrix[68][15] * vector[68] +matrix[69][15] * vector[69] +matrix[70][15] * vector[70] +matrix[71][15] * vector[71] +matrix[72][15] * vector[72] +matrix[73][15] * vector[73] +matrix[74][15] * vector[74] +matrix[75][15] * vector[75] +matrix[76][15] * vector[76] +matrix[77][15] * vector[77] +matrix[78][15] * vector[78] +matrix[79][15] * vector[79] +matrix[80][15] * vector[80] +matrix[81][15] * vector[81] +matrix[82][15] * vector[82] +matrix[83][15] * vector[83] +matrix[84][15] * vector[84] +matrix[85][15] * vector[85] +matrix[86][15] * vector[86] +matrix[87][15] * vector[87] +matrix[88][15] * vector[88] +matrix[89][15] * vector[89] +matrix[90][15] * vector[90] +matrix[91][15] * vector[91] +matrix[92][15] * vector[92] +matrix[93][15] * vector[93] +matrix[94][15] * vector[94] +matrix[95][15] * vector[95] +matrix[96][15] * vector[96] +matrix[97][15] * vector[97] +matrix[98][15] * vector[98] +matrix[99][15] * vector[99] +b[15];
assign result[16] = matrix[0][16] * vector[0] +matrix[1][16] * vector[1] +matrix[2][16] * vector[2] +matrix[3][16] * vector[3] +matrix[4][16] * vector[4] +matrix[5][16] * vector[5] +matrix[6][16] * vector[6] +matrix[7][16] * vector[7] +matrix[8][16] * vector[8] +matrix[9][16] * vector[9] +matrix[10][16] * vector[10] +matrix[11][16] * vector[11] +matrix[12][16] * vector[12] +matrix[13][16] * vector[13] +matrix[14][16] * vector[14] +matrix[15][16] * vector[15] +matrix[16][16] * vector[16] +matrix[17][16] * vector[17] +matrix[18][16] * vector[18] +matrix[19][16] * vector[19] +matrix[20][16] * vector[20] +matrix[21][16] * vector[21] +matrix[22][16] * vector[22] +matrix[23][16] * vector[23] +matrix[24][16] * vector[24] +matrix[25][16] * vector[25] +matrix[26][16] * vector[26] +matrix[27][16] * vector[27] +matrix[28][16] * vector[28] +matrix[29][16] * vector[29] +matrix[30][16] * vector[30] +matrix[31][16] * vector[31] +matrix[32][16] * vector[32] +matrix[33][16] * vector[33] +matrix[34][16] * vector[34] +matrix[35][16] * vector[35] +matrix[36][16] * vector[36] +matrix[37][16] * vector[37] +matrix[38][16] * vector[38] +matrix[39][16] * vector[39] +matrix[40][16] * vector[40] +matrix[41][16] * vector[41] +matrix[42][16] * vector[42] +matrix[43][16] * vector[43] +matrix[44][16] * vector[44] +matrix[45][16] * vector[45] +matrix[46][16] * vector[46] +matrix[47][16] * vector[47] +matrix[48][16] * vector[48] +matrix[49][16] * vector[49] +matrix[50][16] * vector[50] +matrix[51][16] * vector[51] +matrix[52][16] * vector[52] +matrix[53][16] * vector[53] +matrix[54][16] * vector[54] +matrix[55][16] * vector[55] +matrix[56][16] * vector[56] +matrix[57][16] * vector[57] +matrix[58][16] * vector[58] +matrix[59][16] * vector[59] +matrix[60][16] * vector[60] +matrix[61][16] * vector[61] +matrix[62][16] * vector[62] +matrix[63][16] * vector[63] +matrix[64][16] * vector[64] +matrix[65][16] * vector[65] +matrix[66][16] * vector[66] +matrix[67][16] * vector[67] +matrix[68][16] * vector[68] +matrix[69][16] * vector[69] +matrix[70][16] * vector[70] +matrix[71][16] * vector[71] +matrix[72][16] * vector[72] +matrix[73][16] * vector[73] +matrix[74][16] * vector[74] +matrix[75][16] * vector[75] +matrix[76][16] * vector[76] +matrix[77][16] * vector[77] +matrix[78][16] * vector[78] +matrix[79][16] * vector[79] +matrix[80][16] * vector[80] +matrix[81][16] * vector[81] +matrix[82][16] * vector[82] +matrix[83][16] * vector[83] +matrix[84][16] * vector[84] +matrix[85][16] * vector[85] +matrix[86][16] * vector[86] +matrix[87][16] * vector[87] +matrix[88][16] * vector[88] +matrix[89][16] * vector[89] +matrix[90][16] * vector[90] +matrix[91][16] * vector[91] +matrix[92][16] * vector[92] +matrix[93][16] * vector[93] +matrix[94][16] * vector[94] +matrix[95][16] * vector[95] +matrix[96][16] * vector[96] +matrix[97][16] * vector[97] +matrix[98][16] * vector[98] +matrix[99][16] * vector[99] +b[16];
assign result[17] = matrix[0][17] * vector[0] +matrix[1][17] * vector[1] +matrix[2][17] * vector[2] +matrix[3][17] * vector[3] +matrix[4][17] * vector[4] +matrix[5][17] * vector[5] +matrix[6][17] * vector[6] +matrix[7][17] * vector[7] +matrix[8][17] * vector[8] +matrix[9][17] * vector[9] +matrix[10][17] * vector[10] +matrix[11][17] * vector[11] +matrix[12][17] * vector[12] +matrix[13][17] * vector[13] +matrix[14][17] * vector[14] +matrix[15][17] * vector[15] +matrix[16][17] * vector[16] +matrix[17][17] * vector[17] +matrix[18][17] * vector[18] +matrix[19][17] * vector[19] +matrix[20][17] * vector[20] +matrix[21][17] * vector[21] +matrix[22][17] * vector[22] +matrix[23][17] * vector[23] +matrix[24][17] * vector[24] +matrix[25][17] * vector[25] +matrix[26][17] * vector[26] +matrix[27][17] * vector[27] +matrix[28][17] * vector[28] +matrix[29][17] * vector[29] +matrix[30][17] * vector[30] +matrix[31][17] * vector[31] +matrix[32][17] * vector[32] +matrix[33][17] * vector[33] +matrix[34][17] * vector[34] +matrix[35][17] * vector[35] +matrix[36][17] * vector[36] +matrix[37][17] * vector[37] +matrix[38][17] * vector[38] +matrix[39][17] * vector[39] +matrix[40][17] * vector[40] +matrix[41][17] * vector[41] +matrix[42][17] * vector[42] +matrix[43][17] * vector[43] +matrix[44][17] * vector[44] +matrix[45][17] * vector[45] +matrix[46][17] * vector[46] +matrix[47][17] * vector[47] +matrix[48][17] * vector[48] +matrix[49][17] * vector[49] +matrix[50][17] * vector[50] +matrix[51][17] * vector[51] +matrix[52][17] * vector[52] +matrix[53][17] * vector[53] +matrix[54][17] * vector[54] +matrix[55][17] * vector[55] +matrix[56][17] * vector[56] +matrix[57][17] * vector[57] +matrix[58][17] * vector[58] +matrix[59][17] * vector[59] +matrix[60][17] * vector[60] +matrix[61][17] * vector[61] +matrix[62][17] * vector[62] +matrix[63][17] * vector[63] +matrix[64][17] * vector[64] +matrix[65][17] * vector[65] +matrix[66][17] * vector[66] +matrix[67][17] * vector[67] +matrix[68][17] * vector[68] +matrix[69][17] * vector[69] +matrix[70][17] * vector[70] +matrix[71][17] * vector[71] +matrix[72][17] * vector[72] +matrix[73][17] * vector[73] +matrix[74][17] * vector[74] +matrix[75][17] * vector[75] +matrix[76][17] * vector[76] +matrix[77][17] * vector[77] +matrix[78][17] * vector[78] +matrix[79][17] * vector[79] +matrix[80][17] * vector[80] +matrix[81][17] * vector[81] +matrix[82][17] * vector[82] +matrix[83][17] * vector[83] +matrix[84][17] * vector[84] +matrix[85][17] * vector[85] +matrix[86][17] * vector[86] +matrix[87][17] * vector[87] +matrix[88][17] * vector[88] +matrix[89][17] * vector[89] +matrix[90][17] * vector[90] +matrix[91][17] * vector[91] +matrix[92][17] * vector[92] +matrix[93][17] * vector[93] +matrix[94][17] * vector[94] +matrix[95][17] * vector[95] +matrix[96][17] * vector[96] +matrix[97][17] * vector[97] +matrix[98][17] * vector[98] +matrix[99][17] * vector[99] +b[17];
assign result[18] = matrix[0][18] * vector[0] +matrix[1][18] * vector[1] +matrix[2][18] * vector[2] +matrix[3][18] * vector[3] +matrix[4][18] * vector[4] +matrix[5][18] * vector[5] +matrix[6][18] * vector[6] +matrix[7][18] * vector[7] +matrix[8][18] * vector[8] +matrix[9][18] * vector[9] +matrix[10][18] * vector[10] +matrix[11][18] * vector[11] +matrix[12][18] * vector[12] +matrix[13][18] * vector[13] +matrix[14][18] * vector[14] +matrix[15][18] * vector[15] +matrix[16][18] * vector[16] +matrix[17][18] * vector[17] +matrix[18][18] * vector[18] +matrix[19][18] * vector[19] +matrix[20][18] * vector[20] +matrix[21][18] * vector[21] +matrix[22][18] * vector[22] +matrix[23][18] * vector[23] +matrix[24][18] * vector[24] +matrix[25][18] * vector[25] +matrix[26][18] * vector[26] +matrix[27][18] * vector[27] +matrix[28][18] * vector[28] +matrix[29][18] * vector[29] +matrix[30][18] * vector[30] +matrix[31][18] * vector[31] +matrix[32][18] * vector[32] +matrix[33][18] * vector[33] +matrix[34][18] * vector[34] +matrix[35][18] * vector[35] +matrix[36][18] * vector[36] +matrix[37][18] * vector[37] +matrix[38][18] * vector[38] +matrix[39][18] * vector[39] +matrix[40][18] * vector[40] +matrix[41][18] * vector[41] +matrix[42][18] * vector[42] +matrix[43][18] * vector[43] +matrix[44][18] * vector[44] +matrix[45][18] * vector[45] +matrix[46][18] * vector[46] +matrix[47][18] * vector[47] +matrix[48][18] * vector[48] +matrix[49][18] * vector[49] +matrix[50][18] * vector[50] +matrix[51][18] * vector[51] +matrix[52][18] * vector[52] +matrix[53][18] * vector[53] +matrix[54][18] * vector[54] +matrix[55][18] * vector[55] +matrix[56][18] * vector[56] +matrix[57][18] * vector[57] +matrix[58][18] * vector[58] +matrix[59][18] * vector[59] +matrix[60][18] * vector[60] +matrix[61][18] * vector[61] +matrix[62][18] * vector[62] +matrix[63][18] * vector[63] +matrix[64][18] * vector[64] +matrix[65][18] * vector[65] +matrix[66][18] * vector[66] +matrix[67][18] * vector[67] +matrix[68][18] * vector[68] +matrix[69][18] * vector[69] +matrix[70][18] * vector[70] +matrix[71][18] * vector[71] +matrix[72][18] * vector[72] +matrix[73][18] * vector[73] +matrix[74][18] * vector[74] +matrix[75][18] * vector[75] +matrix[76][18] * vector[76] +matrix[77][18] * vector[77] +matrix[78][18] * vector[78] +matrix[79][18] * vector[79] +matrix[80][18] * vector[80] +matrix[81][18] * vector[81] +matrix[82][18] * vector[82] +matrix[83][18] * vector[83] +matrix[84][18] * vector[84] +matrix[85][18] * vector[85] +matrix[86][18] * vector[86] +matrix[87][18] * vector[87] +matrix[88][18] * vector[88] +matrix[89][18] * vector[89] +matrix[90][18] * vector[90] +matrix[91][18] * vector[91] +matrix[92][18] * vector[92] +matrix[93][18] * vector[93] +matrix[94][18] * vector[94] +matrix[95][18] * vector[95] +matrix[96][18] * vector[96] +matrix[97][18] * vector[97] +matrix[98][18] * vector[98] +matrix[99][18] * vector[99] +b[18];
assign result[19] = matrix[0][19] * vector[0] +matrix[1][19] * vector[1] +matrix[2][19] * vector[2] +matrix[3][19] * vector[3] +matrix[4][19] * vector[4] +matrix[5][19] * vector[5] +matrix[6][19] * vector[6] +matrix[7][19] * vector[7] +matrix[8][19] * vector[8] +matrix[9][19] * vector[9] +matrix[10][19] * vector[10] +matrix[11][19] * vector[11] +matrix[12][19] * vector[12] +matrix[13][19] * vector[13] +matrix[14][19] * vector[14] +matrix[15][19] * vector[15] +matrix[16][19] * vector[16] +matrix[17][19] * vector[17] +matrix[18][19] * vector[18] +matrix[19][19] * vector[19] +matrix[20][19] * vector[20] +matrix[21][19] * vector[21] +matrix[22][19] * vector[22] +matrix[23][19] * vector[23] +matrix[24][19] * vector[24] +matrix[25][19] * vector[25] +matrix[26][19] * vector[26] +matrix[27][19] * vector[27] +matrix[28][19] * vector[28] +matrix[29][19] * vector[29] +matrix[30][19] * vector[30] +matrix[31][19] * vector[31] +matrix[32][19] * vector[32] +matrix[33][19] * vector[33] +matrix[34][19] * vector[34] +matrix[35][19] * vector[35] +matrix[36][19] * vector[36] +matrix[37][19] * vector[37] +matrix[38][19] * vector[38] +matrix[39][19] * vector[39] +matrix[40][19] * vector[40] +matrix[41][19] * vector[41] +matrix[42][19] * vector[42] +matrix[43][19] * vector[43] +matrix[44][19] * vector[44] +matrix[45][19] * vector[45] +matrix[46][19] * vector[46] +matrix[47][19] * vector[47] +matrix[48][19] * vector[48] +matrix[49][19] * vector[49] +matrix[50][19] * vector[50] +matrix[51][19] * vector[51] +matrix[52][19] * vector[52] +matrix[53][19] * vector[53] +matrix[54][19] * vector[54] +matrix[55][19] * vector[55] +matrix[56][19] * vector[56] +matrix[57][19] * vector[57] +matrix[58][19] * vector[58] +matrix[59][19] * vector[59] +matrix[60][19] * vector[60] +matrix[61][19] * vector[61] +matrix[62][19] * vector[62] +matrix[63][19] * vector[63] +matrix[64][19] * vector[64] +matrix[65][19] * vector[65] +matrix[66][19] * vector[66] +matrix[67][19] * vector[67] +matrix[68][19] * vector[68] +matrix[69][19] * vector[69] +matrix[70][19] * vector[70] +matrix[71][19] * vector[71] +matrix[72][19] * vector[72] +matrix[73][19] * vector[73] +matrix[74][19] * vector[74] +matrix[75][19] * vector[75] +matrix[76][19] * vector[76] +matrix[77][19] * vector[77] +matrix[78][19] * vector[78] +matrix[79][19] * vector[79] +matrix[80][19] * vector[80] +matrix[81][19] * vector[81] +matrix[82][19] * vector[82] +matrix[83][19] * vector[83] +matrix[84][19] * vector[84] +matrix[85][19] * vector[85] +matrix[86][19] * vector[86] +matrix[87][19] * vector[87] +matrix[88][19] * vector[88] +matrix[89][19] * vector[89] +matrix[90][19] * vector[90] +matrix[91][19] * vector[91] +matrix[92][19] * vector[92] +matrix[93][19] * vector[93] +matrix[94][19] * vector[94] +matrix[95][19] * vector[95] +matrix[96][19] * vector[96] +matrix[97][19] * vector[97] +matrix[98][19] * vector[98] +matrix[99][19] * vector[99] +b[19];
assign result[20] = matrix[0][20] * vector[0] +matrix[1][20] * vector[1] +matrix[2][20] * vector[2] +matrix[3][20] * vector[3] +matrix[4][20] * vector[4] +matrix[5][20] * vector[5] +matrix[6][20] * vector[6] +matrix[7][20] * vector[7] +matrix[8][20] * vector[8] +matrix[9][20] * vector[9] +matrix[10][20] * vector[10] +matrix[11][20] * vector[11] +matrix[12][20] * vector[12] +matrix[13][20] * vector[13] +matrix[14][20] * vector[14] +matrix[15][20] * vector[15] +matrix[16][20] * vector[16] +matrix[17][20] * vector[17] +matrix[18][20] * vector[18] +matrix[19][20] * vector[19] +matrix[20][20] * vector[20] +matrix[21][20] * vector[21] +matrix[22][20] * vector[22] +matrix[23][20] * vector[23] +matrix[24][20] * vector[24] +matrix[25][20] * vector[25] +matrix[26][20] * vector[26] +matrix[27][20] * vector[27] +matrix[28][20] * vector[28] +matrix[29][20] * vector[29] +matrix[30][20] * vector[30] +matrix[31][20] * vector[31] +matrix[32][20] * vector[32] +matrix[33][20] * vector[33] +matrix[34][20] * vector[34] +matrix[35][20] * vector[35] +matrix[36][20] * vector[36] +matrix[37][20] * vector[37] +matrix[38][20] * vector[38] +matrix[39][20] * vector[39] +matrix[40][20] * vector[40] +matrix[41][20] * vector[41] +matrix[42][20] * vector[42] +matrix[43][20] * vector[43] +matrix[44][20] * vector[44] +matrix[45][20] * vector[45] +matrix[46][20] * vector[46] +matrix[47][20] * vector[47] +matrix[48][20] * vector[48] +matrix[49][20] * vector[49] +matrix[50][20] * vector[50] +matrix[51][20] * vector[51] +matrix[52][20] * vector[52] +matrix[53][20] * vector[53] +matrix[54][20] * vector[54] +matrix[55][20] * vector[55] +matrix[56][20] * vector[56] +matrix[57][20] * vector[57] +matrix[58][20] * vector[58] +matrix[59][20] * vector[59] +matrix[60][20] * vector[60] +matrix[61][20] * vector[61] +matrix[62][20] * vector[62] +matrix[63][20] * vector[63] +matrix[64][20] * vector[64] +matrix[65][20] * vector[65] +matrix[66][20] * vector[66] +matrix[67][20] * vector[67] +matrix[68][20] * vector[68] +matrix[69][20] * vector[69] +matrix[70][20] * vector[70] +matrix[71][20] * vector[71] +matrix[72][20] * vector[72] +matrix[73][20] * vector[73] +matrix[74][20] * vector[74] +matrix[75][20] * vector[75] +matrix[76][20] * vector[76] +matrix[77][20] * vector[77] +matrix[78][20] * vector[78] +matrix[79][20] * vector[79] +matrix[80][20] * vector[80] +matrix[81][20] * vector[81] +matrix[82][20] * vector[82] +matrix[83][20] * vector[83] +matrix[84][20] * vector[84] +matrix[85][20] * vector[85] +matrix[86][20] * vector[86] +matrix[87][20] * vector[87] +matrix[88][20] * vector[88] +matrix[89][20] * vector[89] +matrix[90][20] * vector[90] +matrix[91][20] * vector[91] +matrix[92][20] * vector[92] +matrix[93][20] * vector[93] +matrix[94][20] * vector[94] +matrix[95][20] * vector[95] +matrix[96][20] * vector[96] +matrix[97][20] * vector[97] +matrix[98][20] * vector[98] +matrix[99][20] * vector[99] +b[20];
assign result[21] = matrix[0][21] * vector[0] +matrix[1][21] * vector[1] +matrix[2][21] * vector[2] +matrix[3][21] * vector[3] +matrix[4][21] * vector[4] +matrix[5][21] * vector[5] +matrix[6][21] * vector[6] +matrix[7][21] * vector[7] +matrix[8][21] * vector[8] +matrix[9][21] * vector[9] +matrix[10][21] * vector[10] +matrix[11][21] * vector[11] +matrix[12][21] * vector[12] +matrix[13][21] * vector[13] +matrix[14][21] * vector[14] +matrix[15][21] * vector[15] +matrix[16][21] * vector[16] +matrix[17][21] * vector[17] +matrix[18][21] * vector[18] +matrix[19][21] * vector[19] +matrix[20][21] * vector[20] +matrix[21][21] * vector[21] +matrix[22][21] * vector[22] +matrix[23][21] * vector[23] +matrix[24][21] * vector[24] +matrix[25][21] * vector[25] +matrix[26][21] * vector[26] +matrix[27][21] * vector[27] +matrix[28][21] * vector[28] +matrix[29][21] * vector[29] +matrix[30][21] * vector[30] +matrix[31][21] * vector[31] +matrix[32][21] * vector[32] +matrix[33][21] * vector[33] +matrix[34][21] * vector[34] +matrix[35][21] * vector[35] +matrix[36][21] * vector[36] +matrix[37][21] * vector[37] +matrix[38][21] * vector[38] +matrix[39][21] * vector[39] +matrix[40][21] * vector[40] +matrix[41][21] * vector[41] +matrix[42][21] * vector[42] +matrix[43][21] * vector[43] +matrix[44][21] * vector[44] +matrix[45][21] * vector[45] +matrix[46][21] * vector[46] +matrix[47][21] * vector[47] +matrix[48][21] * vector[48] +matrix[49][21] * vector[49] +matrix[50][21] * vector[50] +matrix[51][21] * vector[51] +matrix[52][21] * vector[52] +matrix[53][21] * vector[53] +matrix[54][21] * vector[54] +matrix[55][21] * vector[55] +matrix[56][21] * vector[56] +matrix[57][21] * vector[57] +matrix[58][21] * vector[58] +matrix[59][21] * vector[59] +matrix[60][21] * vector[60] +matrix[61][21] * vector[61] +matrix[62][21] * vector[62] +matrix[63][21] * vector[63] +matrix[64][21] * vector[64] +matrix[65][21] * vector[65] +matrix[66][21] * vector[66] +matrix[67][21] * vector[67] +matrix[68][21] * vector[68] +matrix[69][21] * vector[69] +matrix[70][21] * vector[70] +matrix[71][21] * vector[71] +matrix[72][21] * vector[72] +matrix[73][21] * vector[73] +matrix[74][21] * vector[74] +matrix[75][21] * vector[75] +matrix[76][21] * vector[76] +matrix[77][21] * vector[77] +matrix[78][21] * vector[78] +matrix[79][21] * vector[79] +matrix[80][21] * vector[80] +matrix[81][21] * vector[81] +matrix[82][21] * vector[82] +matrix[83][21] * vector[83] +matrix[84][21] * vector[84] +matrix[85][21] * vector[85] +matrix[86][21] * vector[86] +matrix[87][21] * vector[87] +matrix[88][21] * vector[88] +matrix[89][21] * vector[89] +matrix[90][21] * vector[90] +matrix[91][21] * vector[91] +matrix[92][21] * vector[92] +matrix[93][21] * vector[93] +matrix[94][21] * vector[94] +matrix[95][21] * vector[95] +matrix[96][21] * vector[96] +matrix[97][21] * vector[97] +matrix[98][21] * vector[98] +matrix[99][21] * vector[99] +b[21];
assign result[22] = matrix[0][22] * vector[0] +matrix[1][22] * vector[1] +matrix[2][22] * vector[2] +matrix[3][22] * vector[3] +matrix[4][22] * vector[4] +matrix[5][22] * vector[5] +matrix[6][22] * vector[6] +matrix[7][22] * vector[7] +matrix[8][22] * vector[8] +matrix[9][22] * vector[9] +matrix[10][22] * vector[10] +matrix[11][22] * vector[11] +matrix[12][22] * vector[12] +matrix[13][22] * vector[13] +matrix[14][22] * vector[14] +matrix[15][22] * vector[15] +matrix[16][22] * vector[16] +matrix[17][22] * vector[17] +matrix[18][22] * vector[18] +matrix[19][22] * vector[19] +matrix[20][22] * vector[20] +matrix[21][22] * vector[21] +matrix[22][22] * vector[22] +matrix[23][22] * vector[23] +matrix[24][22] * vector[24] +matrix[25][22] * vector[25] +matrix[26][22] * vector[26] +matrix[27][22] * vector[27] +matrix[28][22] * vector[28] +matrix[29][22] * vector[29] +matrix[30][22] * vector[30] +matrix[31][22] * vector[31] +matrix[32][22] * vector[32] +matrix[33][22] * vector[33] +matrix[34][22] * vector[34] +matrix[35][22] * vector[35] +matrix[36][22] * vector[36] +matrix[37][22] * vector[37] +matrix[38][22] * vector[38] +matrix[39][22] * vector[39] +matrix[40][22] * vector[40] +matrix[41][22] * vector[41] +matrix[42][22] * vector[42] +matrix[43][22] * vector[43] +matrix[44][22] * vector[44] +matrix[45][22] * vector[45] +matrix[46][22] * vector[46] +matrix[47][22] * vector[47] +matrix[48][22] * vector[48] +matrix[49][22] * vector[49] +matrix[50][22] * vector[50] +matrix[51][22] * vector[51] +matrix[52][22] * vector[52] +matrix[53][22] * vector[53] +matrix[54][22] * vector[54] +matrix[55][22] * vector[55] +matrix[56][22] * vector[56] +matrix[57][22] * vector[57] +matrix[58][22] * vector[58] +matrix[59][22] * vector[59] +matrix[60][22] * vector[60] +matrix[61][22] * vector[61] +matrix[62][22] * vector[62] +matrix[63][22] * vector[63] +matrix[64][22] * vector[64] +matrix[65][22] * vector[65] +matrix[66][22] * vector[66] +matrix[67][22] * vector[67] +matrix[68][22] * vector[68] +matrix[69][22] * vector[69] +matrix[70][22] * vector[70] +matrix[71][22] * vector[71] +matrix[72][22] * vector[72] +matrix[73][22] * vector[73] +matrix[74][22] * vector[74] +matrix[75][22] * vector[75] +matrix[76][22] * vector[76] +matrix[77][22] * vector[77] +matrix[78][22] * vector[78] +matrix[79][22] * vector[79] +matrix[80][22] * vector[80] +matrix[81][22] * vector[81] +matrix[82][22] * vector[82] +matrix[83][22] * vector[83] +matrix[84][22] * vector[84] +matrix[85][22] * vector[85] +matrix[86][22] * vector[86] +matrix[87][22] * vector[87] +matrix[88][22] * vector[88] +matrix[89][22] * vector[89] +matrix[90][22] * vector[90] +matrix[91][22] * vector[91] +matrix[92][22] * vector[92] +matrix[93][22] * vector[93] +matrix[94][22] * vector[94] +matrix[95][22] * vector[95] +matrix[96][22] * vector[96] +matrix[97][22] * vector[97] +matrix[98][22] * vector[98] +matrix[99][22] * vector[99] +b[22];
assign result[23] = matrix[0][23] * vector[0] +matrix[1][23] * vector[1] +matrix[2][23] * vector[2] +matrix[3][23] * vector[3] +matrix[4][23] * vector[4] +matrix[5][23] * vector[5] +matrix[6][23] * vector[6] +matrix[7][23] * vector[7] +matrix[8][23] * vector[8] +matrix[9][23] * vector[9] +matrix[10][23] * vector[10] +matrix[11][23] * vector[11] +matrix[12][23] * vector[12] +matrix[13][23] * vector[13] +matrix[14][23] * vector[14] +matrix[15][23] * vector[15] +matrix[16][23] * vector[16] +matrix[17][23] * vector[17] +matrix[18][23] * vector[18] +matrix[19][23] * vector[19] +matrix[20][23] * vector[20] +matrix[21][23] * vector[21] +matrix[22][23] * vector[22] +matrix[23][23] * vector[23] +matrix[24][23] * vector[24] +matrix[25][23] * vector[25] +matrix[26][23] * vector[26] +matrix[27][23] * vector[27] +matrix[28][23] * vector[28] +matrix[29][23] * vector[29] +matrix[30][23] * vector[30] +matrix[31][23] * vector[31] +matrix[32][23] * vector[32] +matrix[33][23] * vector[33] +matrix[34][23] * vector[34] +matrix[35][23] * vector[35] +matrix[36][23] * vector[36] +matrix[37][23] * vector[37] +matrix[38][23] * vector[38] +matrix[39][23] * vector[39] +matrix[40][23] * vector[40] +matrix[41][23] * vector[41] +matrix[42][23] * vector[42] +matrix[43][23] * vector[43] +matrix[44][23] * vector[44] +matrix[45][23] * vector[45] +matrix[46][23] * vector[46] +matrix[47][23] * vector[47] +matrix[48][23] * vector[48] +matrix[49][23] * vector[49] +matrix[50][23] * vector[50] +matrix[51][23] * vector[51] +matrix[52][23] * vector[52] +matrix[53][23] * vector[53] +matrix[54][23] * vector[54] +matrix[55][23] * vector[55] +matrix[56][23] * vector[56] +matrix[57][23] * vector[57] +matrix[58][23] * vector[58] +matrix[59][23] * vector[59] +matrix[60][23] * vector[60] +matrix[61][23] * vector[61] +matrix[62][23] * vector[62] +matrix[63][23] * vector[63] +matrix[64][23] * vector[64] +matrix[65][23] * vector[65] +matrix[66][23] * vector[66] +matrix[67][23] * vector[67] +matrix[68][23] * vector[68] +matrix[69][23] * vector[69] +matrix[70][23] * vector[70] +matrix[71][23] * vector[71] +matrix[72][23] * vector[72] +matrix[73][23] * vector[73] +matrix[74][23] * vector[74] +matrix[75][23] * vector[75] +matrix[76][23] * vector[76] +matrix[77][23] * vector[77] +matrix[78][23] * vector[78] +matrix[79][23] * vector[79] +matrix[80][23] * vector[80] +matrix[81][23] * vector[81] +matrix[82][23] * vector[82] +matrix[83][23] * vector[83] +matrix[84][23] * vector[84] +matrix[85][23] * vector[85] +matrix[86][23] * vector[86] +matrix[87][23] * vector[87] +matrix[88][23] * vector[88] +matrix[89][23] * vector[89] +matrix[90][23] * vector[90] +matrix[91][23] * vector[91] +matrix[92][23] * vector[92] +matrix[93][23] * vector[93] +matrix[94][23] * vector[94] +matrix[95][23] * vector[95] +matrix[96][23] * vector[96] +matrix[97][23] * vector[97] +matrix[98][23] * vector[98] +matrix[99][23] * vector[99] +b[23];
assign result[24] = matrix[0][24] * vector[0] +matrix[1][24] * vector[1] +matrix[2][24] * vector[2] +matrix[3][24] * vector[3] +matrix[4][24] * vector[4] +matrix[5][24] * vector[5] +matrix[6][24] * vector[6] +matrix[7][24] * vector[7] +matrix[8][24] * vector[8] +matrix[9][24] * vector[9] +matrix[10][24] * vector[10] +matrix[11][24] * vector[11] +matrix[12][24] * vector[12] +matrix[13][24] * vector[13] +matrix[14][24] * vector[14] +matrix[15][24] * vector[15] +matrix[16][24] * vector[16] +matrix[17][24] * vector[17] +matrix[18][24] * vector[18] +matrix[19][24] * vector[19] +matrix[20][24] * vector[20] +matrix[21][24] * vector[21] +matrix[22][24] * vector[22] +matrix[23][24] * vector[23] +matrix[24][24] * vector[24] +matrix[25][24] * vector[25] +matrix[26][24] * vector[26] +matrix[27][24] * vector[27] +matrix[28][24] * vector[28] +matrix[29][24] * vector[29] +matrix[30][24] * vector[30] +matrix[31][24] * vector[31] +matrix[32][24] * vector[32] +matrix[33][24] * vector[33] +matrix[34][24] * vector[34] +matrix[35][24] * vector[35] +matrix[36][24] * vector[36] +matrix[37][24] * vector[37] +matrix[38][24] * vector[38] +matrix[39][24] * vector[39] +matrix[40][24] * vector[40] +matrix[41][24] * vector[41] +matrix[42][24] * vector[42] +matrix[43][24] * vector[43] +matrix[44][24] * vector[44] +matrix[45][24] * vector[45] +matrix[46][24] * vector[46] +matrix[47][24] * vector[47] +matrix[48][24] * vector[48] +matrix[49][24] * vector[49] +matrix[50][24] * vector[50] +matrix[51][24] * vector[51] +matrix[52][24] * vector[52] +matrix[53][24] * vector[53] +matrix[54][24] * vector[54] +matrix[55][24] * vector[55] +matrix[56][24] * vector[56] +matrix[57][24] * vector[57] +matrix[58][24] * vector[58] +matrix[59][24] * vector[59] +matrix[60][24] * vector[60] +matrix[61][24] * vector[61] +matrix[62][24] * vector[62] +matrix[63][24] * vector[63] +matrix[64][24] * vector[64] +matrix[65][24] * vector[65] +matrix[66][24] * vector[66] +matrix[67][24] * vector[67] +matrix[68][24] * vector[68] +matrix[69][24] * vector[69] +matrix[70][24] * vector[70] +matrix[71][24] * vector[71] +matrix[72][24] * vector[72] +matrix[73][24] * vector[73] +matrix[74][24] * vector[74] +matrix[75][24] * vector[75] +matrix[76][24] * vector[76] +matrix[77][24] * vector[77] +matrix[78][24] * vector[78] +matrix[79][24] * vector[79] +matrix[80][24] * vector[80] +matrix[81][24] * vector[81] +matrix[82][24] * vector[82] +matrix[83][24] * vector[83] +matrix[84][24] * vector[84] +matrix[85][24] * vector[85] +matrix[86][24] * vector[86] +matrix[87][24] * vector[87] +matrix[88][24] * vector[88] +matrix[89][24] * vector[89] +matrix[90][24] * vector[90] +matrix[91][24] * vector[91] +matrix[92][24] * vector[92] +matrix[93][24] * vector[93] +matrix[94][24] * vector[94] +matrix[95][24] * vector[95] +matrix[96][24] * vector[96] +matrix[97][24] * vector[97] +matrix[98][24] * vector[98] +matrix[99][24] * vector[99] +b[24];
assign result[25] = matrix[0][25] * vector[0] +matrix[1][25] * vector[1] +matrix[2][25] * vector[2] +matrix[3][25] * vector[3] +matrix[4][25] * vector[4] +matrix[5][25] * vector[5] +matrix[6][25] * vector[6] +matrix[7][25] * vector[7] +matrix[8][25] * vector[8] +matrix[9][25] * vector[9] +matrix[10][25] * vector[10] +matrix[11][25] * vector[11] +matrix[12][25] * vector[12] +matrix[13][25] * vector[13] +matrix[14][25] * vector[14] +matrix[15][25] * vector[15] +matrix[16][25] * vector[16] +matrix[17][25] * vector[17] +matrix[18][25] * vector[18] +matrix[19][25] * vector[19] +matrix[20][25] * vector[20] +matrix[21][25] * vector[21] +matrix[22][25] * vector[22] +matrix[23][25] * vector[23] +matrix[24][25] * vector[24] +matrix[25][25] * vector[25] +matrix[26][25] * vector[26] +matrix[27][25] * vector[27] +matrix[28][25] * vector[28] +matrix[29][25] * vector[29] +matrix[30][25] * vector[30] +matrix[31][25] * vector[31] +matrix[32][25] * vector[32] +matrix[33][25] * vector[33] +matrix[34][25] * vector[34] +matrix[35][25] * vector[35] +matrix[36][25] * vector[36] +matrix[37][25] * vector[37] +matrix[38][25] * vector[38] +matrix[39][25] * vector[39] +matrix[40][25] * vector[40] +matrix[41][25] * vector[41] +matrix[42][25] * vector[42] +matrix[43][25] * vector[43] +matrix[44][25] * vector[44] +matrix[45][25] * vector[45] +matrix[46][25] * vector[46] +matrix[47][25] * vector[47] +matrix[48][25] * vector[48] +matrix[49][25] * vector[49] +matrix[50][25] * vector[50] +matrix[51][25] * vector[51] +matrix[52][25] * vector[52] +matrix[53][25] * vector[53] +matrix[54][25] * vector[54] +matrix[55][25] * vector[55] +matrix[56][25] * vector[56] +matrix[57][25] * vector[57] +matrix[58][25] * vector[58] +matrix[59][25] * vector[59] +matrix[60][25] * vector[60] +matrix[61][25] * vector[61] +matrix[62][25] * vector[62] +matrix[63][25] * vector[63] +matrix[64][25] * vector[64] +matrix[65][25] * vector[65] +matrix[66][25] * vector[66] +matrix[67][25] * vector[67] +matrix[68][25] * vector[68] +matrix[69][25] * vector[69] +matrix[70][25] * vector[70] +matrix[71][25] * vector[71] +matrix[72][25] * vector[72] +matrix[73][25] * vector[73] +matrix[74][25] * vector[74] +matrix[75][25] * vector[75] +matrix[76][25] * vector[76] +matrix[77][25] * vector[77] +matrix[78][25] * vector[78] +matrix[79][25] * vector[79] +matrix[80][25] * vector[80] +matrix[81][25] * vector[81] +matrix[82][25] * vector[82] +matrix[83][25] * vector[83] +matrix[84][25] * vector[84] +matrix[85][25] * vector[85] +matrix[86][25] * vector[86] +matrix[87][25] * vector[87] +matrix[88][25] * vector[88] +matrix[89][25] * vector[89] +matrix[90][25] * vector[90] +matrix[91][25] * vector[91] +matrix[92][25] * vector[92] +matrix[93][25] * vector[93] +matrix[94][25] * vector[94] +matrix[95][25] * vector[95] +matrix[96][25] * vector[96] +matrix[97][25] * vector[97] +matrix[98][25] * vector[98] +matrix[99][25] * vector[99] +b[25];
assign result[26] = matrix[0][26] * vector[0] +matrix[1][26] * vector[1] +matrix[2][26] * vector[2] +matrix[3][26] * vector[3] +matrix[4][26] * vector[4] +matrix[5][26] * vector[5] +matrix[6][26] * vector[6] +matrix[7][26] * vector[7] +matrix[8][26] * vector[8] +matrix[9][26] * vector[9] +matrix[10][26] * vector[10] +matrix[11][26] * vector[11] +matrix[12][26] * vector[12] +matrix[13][26] * vector[13] +matrix[14][26] * vector[14] +matrix[15][26] * vector[15] +matrix[16][26] * vector[16] +matrix[17][26] * vector[17] +matrix[18][26] * vector[18] +matrix[19][26] * vector[19] +matrix[20][26] * vector[20] +matrix[21][26] * vector[21] +matrix[22][26] * vector[22] +matrix[23][26] * vector[23] +matrix[24][26] * vector[24] +matrix[25][26] * vector[25] +matrix[26][26] * vector[26] +matrix[27][26] * vector[27] +matrix[28][26] * vector[28] +matrix[29][26] * vector[29] +matrix[30][26] * vector[30] +matrix[31][26] * vector[31] +matrix[32][26] * vector[32] +matrix[33][26] * vector[33] +matrix[34][26] * vector[34] +matrix[35][26] * vector[35] +matrix[36][26] * vector[36] +matrix[37][26] * vector[37] +matrix[38][26] * vector[38] +matrix[39][26] * vector[39] +matrix[40][26] * vector[40] +matrix[41][26] * vector[41] +matrix[42][26] * vector[42] +matrix[43][26] * vector[43] +matrix[44][26] * vector[44] +matrix[45][26] * vector[45] +matrix[46][26] * vector[46] +matrix[47][26] * vector[47] +matrix[48][26] * vector[48] +matrix[49][26] * vector[49] +matrix[50][26] * vector[50] +matrix[51][26] * vector[51] +matrix[52][26] * vector[52] +matrix[53][26] * vector[53] +matrix[54][26] * vector[54] +matrix[55][26] * vector[55] +matrix[56][26] * vector[56] +matrix[57][26] * vector[57] +matrix[58][26] * vector[58] +matrix[59][26] * vector[59] +matrix[60][26] * vector[60] +matrix[61][26] * vector[61] +matrix[62][26] * vector[62] +matrix[63][26] * vector[63] +matrix[64][26] * vector[64] +matrix[65][26] * vector[65] +matrix[66][26] * vector[66] +matrix[67][26] * vector[67] +matrix[68][26] * vector[68] +matrix[69][26] * vector[69] +matrix[70][26] * vector[70] +matrix[71][26] * vector[71] +matrix[72][26] * vector[72] +matrix[73][26] * vector[73] +matrix[74][26] * vector[74] +matrix[75][26] * vector[75] +matrix[76][26] * vector[76] +matrix[77][26] * vector[77] +matrix[78][26] * vector[78] +matrix[79][26] * vector[79] +matrix[80][26] * vector[80] +matrix[81][26] * vector[81] +matrix[82][26] * vector[82] +matrix[83][26] * vector[83] +matrix[84][26] * vector[84] +matrix[85][26] * vector[85] +matrix[86][26] * vector[86] +matrix[87][26] * vector[87] +matrix[88][26] * vector[88] +matrix[89][26] * vector[89] +matrix[90][26] * vector[90] +matrix[91][26] * vector[91] +matrix[92][26] * vector[92] +matrix[93][26] * vector[93] +matrix[94][26] * vector[94] +matrix[95][26] * vector[95] +matrix[96][26] * vector[96] +matrix[97][26] * vector[97] +matrix[98][26] * vector[98] +matrix[99][26] * vector[99] +b[26];
assign result[27] = matrix[0][27] * vector[0] +matrix[1][27] * vector[1] +matrix[2][27] * vector[2] +matrix[3][27] * vector[3] +matrix[4][27] * vector[4] +matrix[5][27] * vector[5] +matrix[6][27] * vector[6] +matrix[7][27] * vector[7] +matrix[8][27] * vector[8] +matrix[9][27] * vector[9] +matrix[10][27] * vector[10] +matrix[11][27] * vector[11] +matrix[12][27] * vector[12] +matrix[13][27] * vector[13] +matrix[14][27] * vector[14] +matrix[15][27] * vector[15] +matrix[16][27] * vector[16] +matrix[17][27] * vector[17] +matrix[18][27] * vector[18] +matrix[19][27] * vector[19] +matrix[20][27] * vector[20] +matrix[21][27] * vector[21] +matrix[22][27] * vector[22] +matrix[23][27] * vector[23] +matrix[24][27] * vector[24] +matrix[25][27] * vector[25] +matrix[26][27] * vector[26] +matrix[27][27] * vector[27] +matrix[28][27] * vector[28] +matrix[29][27] * vector[29] +matrix[30][27] * vector[30] +matrix[31][27] * vector[31] +matrix[32][27] * vector[32] +matrix[33][27] * vector[33] +matrix[34][27] * vector[34] +matrix[35][27] * vector[35] +matrix[36][27] * vector[36] +matrix[37][27] * vector[37] +matrix[38][27] * vector[38] +matrix[39][27] * vector[39] +matrix[40][27] * vector[40] +matrix[41][27] * vector[41] +matrix[42][27] * vector[42] +matrix[43][27] * vector[43] +matrix[44][27] * vector[44] +matrix[45][27] * vector[45] +matrix[46][27] * vector[46] +matrix[47][27] * vector[47] +matrix[48][27] * vector[48] +matrix[49][27] * vector[49] +matrix[50][27] * vector[50] +matrix[51][27] * vector[51] +matrix[52][27] * vector[52] +matrix[53][27] * vector[53] +matrix[54][27] * vector[54] +matrix[55][27] * vector[55] +matrix[56][27] * vector[56] +matrix[57][27] * vector[57] +matrix[58][27] * vector[58] +matrix[59][27] * vector[59] +matrix[60][27] * vector[60] +matrix[61][27] * vector[61] +matrix[62][27] * vector[62] +matrix[63][27] * vector[63] +matrix[64][27] * vector[64] +matrix[65][27] * vector[65] +matrix[66][27] * vector[66] +matrix[67][27] * vector[67] +matrix[68][27] * vector[68] +matrix[69][27] * vector[69] +matrix[70][27] * vector[70] +matrix[71][27] * vector[71] +matrix[72][27] * vector[72] +matrix[73][27] * vector[73] +matrix[74][27] * vector[74] +matrix[75][27] * vector[75] +matrix[76][27] * vector[76] +matrix[77][27] * vector[77] +matrix[78][27] * vector[78] +matrix[79][27] * vector[79] +matrix[80][27] * vector[80] +matrix[81][27] * vector[81] +matrix[82][27] * vector[82] +matrix[83][27] * vector[83] +matrix[84][27] * vector[84] +matrix[85][27] * vector[85] +matrix[86][27] * vector[86] +matrix[87][27] * vector[87] +matrix[88][27] * vector[88] +matrix[89][27] * vector[89] +matrix[90][27] * vector[90] +matrix[91][27] * vector[91] +matrix[92][27] * vector[92] +matrix[93][27] * vector[93] +matrix[94][27] * vector[94] +matrix[95][27] * vector[95] +matrix[96][27] * vector[96] +matrix[97][27] * vector[97] +matrix[98][27] * vector[98] +matrix[99][27] * vector[99] +b[27];
assign result[28] = matrix[0][28] * vector[0] +matrix[1][28] * vector[1] +matrix[2][28] * vector[2] +matrix[3][28] * vector[3] +matrix[4][28] * vector[4] +matrix[5][28] * vector[5] +matrix[6][28] * vector[6] +matrix[7][28] * vector[7] +matrix[8][28] * vector[8] +matrix[9][28] * vector[9] +matrix[10][28] * vector[10] +matrix[11][28] * vector[11] +matrix[12][28] * vector[12] +matrix[13][28] * vector[13] +matrix[14][28] * vector[14] +matrix[15][28] * vector[15] +matrix[16][28] * vector[16] +matrix[17][28] * vector[17] +matrix[18][28] * vector[18] +matrix[19][28] * vector[19] +matrix[20][28] * vector[20] +matrix[21][28] * vector[21] +matrix[22][28] * vector[22] +matrix[23][28] * vector[23] +matrix[24][28] * vector[24] +matrix[25][28] * vector[25] +matrix[26][28] * vector[26] +matrix[27][28] * vector[27] +matrix[28][28] * vector[28] +matrix[29][28] * vector[29] +matrix[30][28] * vector[30] +matrix[31][28] * vector[31] +matrix[32][28] * vector[32] +matrix[33][28] * vector[33] +matrix[34][28] * vector[34] +matrix[35][28] * vector[35] +matrix[36][28] * vector[36] +matrix[37][28] * vector[37] +matrix[38][28] * vector[38] +matrix[39][28] * vector[39] +matrix[40][28] * vector[40] +matrix[41][28] * vector[41] +matrix[42][28] * vector[42] +matrix[43][28] * vector[43] +matrix[44][28] * vector[44] +matrix[45][28] * vector[45] +matrix[46][28] * vector[46] +matrix[47][28] * vector[47] +matrix[48][28] * vector[48] +matrix[49][28] * vector[49] +matrix[50][28] * vector[50] +matrix[51][28] * vector[51] +matrix[52][28] * vector[52] +matrix[53][28] * vector[53] +matrix[54][28] * vector[54] +matrix[55][28] * vector[55] +matrix[56][28] * vector[56] +matrix[57][28] * vector[57] +matrix[58][28] * vector[58] +matrix[59][28] * vector[59] +matrix[60][28] * vector[60] +matrix[61][28] * vector[61] +matrix[62][28] * vector[62] +matrix[63][28] * vector[63] +matrix[64][28] * vector[64] +matrix[65][28] * vector[65] +matrix[66][28] * vector[66] +matrix[67][28] * vector[67] +matrix[68][28] * vector[68] +matrix[69][28] * vector[69] +matrix[70][28] * vector[70] +matrix[71][28] * vector[71] +matrix[72][28] * vector[72] +matrix[73][28] * vector[73] +matrix[74][28] * vector[74] +matrix[75][28] * vector[75] +matrix[76][28] * vector[76] +matrix[77][28] * vector[77] +matrix[78][28] * vector[78] +matrix[79][28] * vector[79] +matrix[80][28] * vector[80] +matrix[81][28] * vector[81] +matrix[82][28] * vector[82] +matrix[83][28] * vector[83] +matrix[84][28] * vector[84] +matrix[85][28] * vector[85] +matrix[86][28] * vector[86] +matrix[87][28] * vector[87] +matrix[88][28] * vector[88] +matrix[89][28] * vector[89] +matrix[90][28] * vector[90] +matrix[91][28] * vector[91] +matrix[92][28] * vector[92] +matrix[93][28] * vector[93] +matrix[94][28] * vector[94] +matrix[95][28] * vector[95] +matrix[96][28] * vector[96] +matrix[97][28] * vector[97] +matrix[98][28] * vector[98] +matrix[99][28] * vector[99] +b[28];
assign result[29] = matrix[0][29] * vector[0] +matrix[1][29] * vector[1] +matrix[2][29] * vector[2] +matrix[3][29] * vector[3] +matrix[4][29] * vector[4] +matrix[5][29] * vector[5] +matrix[6][29] * vector[6] +matrix[7][29] * vector[7] +matrix[8][29] * vector[8] +matrix[9][29] * vector[9] +matrix[10][29] * vector[10] +matrix[11][29] * vector[11] +matrix[12][29] * vector[12] +matrix[13][29] * vector[13] +matrix[14][29] * vector[14] +matrix[15][29] * vector[15] +matrix[16][29] * vector[16] +matrix[17][29] * vector[17] +matrix[18][29] * vector[18] +matrix[19][29] * vector[19] +matrix[20][29] * vector[20] +matrix[21][29] * vector[21] +matrix[22][29] * vector[22] +matrix[23][29] * vector[23] +matrix[24][29] * vector[24] +matrix[25][29] * vector[25] +matrix[26][29] * vector[26] +matrix[27][29] * vector[27] +matrix[28][29] * vector[28] +matrix[29][29] * vector[29] +matrix[30][29] * vector[30] +matrix[31][29] * vector[31] +matrix[32][29] * vector[32] +matrix[33][29] * vector[33] +matrix[34][29] * vector[34] +matrix[35][29] * vector[35] +matrix[36][29] * vector[36] +matrix[37][29] * vector[37] +matrix[38][29] * vector[38] +matrix[39][29] * vector[39] +matrix[40][29] * vector[40] +matrix[41][29] * vector[41] +matrix[42][29] * vector[42] +matrix[43][29] * vector[43] +matrix[44][29] * vector[44] +matrix[45][29] * vector[45] +matrix[46][29] * vector[46] +matrix[47][29] * vector[47] +matrix[48][29] * vector[48] +matrix[49][29] * vector[49] +matrix[50][29] * vector[50] +matrix[51][29] * vector[51] +matrix[52][29] * vector[52] +matrix[53][29] * vector[53] +matrix[54][29] * vector[54] +matrix[55][29] * vector[55] +matrix[56][29] * vector[56] +matrix[57][29] * vector[57] +matrix[58][29] * vector[58] +matrix[59][29] * vector[59] +matrix[60][29] * vector[60] +matrix[61][29] * vector[61] +matrix[62][29] * vector[62] +matrix[63][29] * vector[63] +matrix[64][29] * vector[64] +matrix[65][29] * vector[65] +matrix[66][29] * vector[66] +matrix[67][29] * vector[67] +matrix[68][29] * vector[68] +matrix[69][29] * vector[69] +matrix[70][29] * vector[70] +matrix[71][29] * vector[71] +matrix[72][29] * vector[72] +matrix[73][29] * vector[73] +matrix[74][29] * vector[74] +matrix[75][29] * vector[75] +matrix[76][29] * vector[76] +matrix[77][29] * vector[77] +matrix[78][29] * vector[78] +matrix[79][29] * vector[79] +matrix[80][29] * vector[80] +matrix[81][29] * vector[81] +matrix[82][29] * vector[82] +matrix[83][29] * vector[83] +matrix[84][29] * vector[84] +matrix[85][29] * vector[85] +matrix[86][29] * vector[86] +matrix[87][29] * vector[87] +matrix[88][29] * vector[88] +matrix[89][29] * vector[89] +matrix[90][29] * vector[90] +matrix[91][29] * vector[91] +matrix[92][29] * vector[92] +matrix[93][29] * vector[93] +matrix[94][29] * vector[94] +matrix[95][29] * vector[95] +matrix[96][29] * vector[96] +matrix[97][29] * vector[97] +matrix[98][29] * vector[98] +matrix[99][29] * vector[99] +b[29];
assign result[30] = matrix[0][30] * vector[0] +matrix[1][30] * vector[1] +matrix[2][30] * vector[2] +matrix[3][30] * vector[3] +matrix[4][30] * vector[4] +matrix[5][30] * vector[5] +matrix[6][30] * vector[6] +matrix[7][30] * vector[7] +matrix[8][30] * vector[8] +matrix[9][30] * vector[9] +matrix[10][30] * vector[10] +matrix[11][30] * vector[11] +matrix[12][30] * vector[12] +matrix[13][30] * vector[13] +matrix[14][30] * vector[14] +matrix[15][30] * vector[15] +matrix[16][30] * vector[16] +matrix[17][30] * vector[17] +matrix[18][30] * vector[18] +matrix[19][30] * vector[19] +matrix[20][30] * vector[20] +matrix[21][30] * vector[21] +matrix[22][30] * vector[22] +matrix[23][30] * vector[23] +matrix[24][30] * vector[24] +matrix[25][30] * vector[25] +matrix[26][30] * vector[26] +matrix[27][30] * vector[27] +matrix[28][30] * vector[28] +matrix[29][30] * vector[29] +matrix[30][30] * vector[30] +matrix[31][30] * vector[31] +matrix[32][30] * vector[32] +matrix[33][30] * vector[33] +matrix[34][30] * vector[34] +matrix[35][30] * vector[35] +matrix[36][30] * vector[36] +matrix[37][30] * vector[37] +matrix[38][30] * vector[38] +matrix[39][30] * vector[39] +matrix[40][30] * vector[40] +matrix[41][30] * vector[41] +matrix[42][30] * vector[42] +matrix[43][30] * vector[43] +matrix[44][30] * vector[44] +matrix[45][30] * vector[45] +matrix[46][30] * vector[46] +matrix[47][30] * vector[47] +matrix[48][30] * vector[48] +matrix[49][30] * vector[49] +matrix[50][30] * vector[50] +matrix[51][30] * vector[51] +matrix[52][30] * vector[52] +matrix[53][30] * vector[53] +matrix[54][30] * vector[54] +matrix[55][30] * vector[55] +matrix[56][30] * vector[56] +matrix[57][30] * vector[57] +matrix[58][30] * vector[58] +matrix[59][30] * vector[59] +matrix[60][30] * vector[60] +matrix[61][30] * vector[61] +matrix[62][30] * vector[62] +matrix[63][30] * vector[63] +matrix[64][30] * vector[64] +matrix[65][30] * vector[65] +matrix[66][30] * vector[66] +matrix[67][30] * vector[67] +matrix[68][30] * vector[68] +matrix[69][30] * vector[69] +matrix[70][30] * vector[70] +matrix[71][30] * vector[71] +matrix[72][30] * vector[72] +matrix[73][30] * vector[73] +matrix[74][30] * vector[74] +matrix[75][30] * vector[75] +matrix[76][30] * vector[76] +matrix[77][30] * vector[77] +matrix[78][30] * vector[78] +matrix[79][30] * vector[79] +matrix[80][30] * vector[80] +matrix[81][30] * vector[81] +matrix[82][30] * vector[82] +matrix[83][30] * vector[83] +matrix[84][30] * vector[84] +matrix[85][30] * vector[85] +matrix[86][30] * vector[86] +matrix[87][30] * vector[87] +matrix[88][30] * vector[88] +matrix[89][30] * vector[89] +matrix[90][30] * vector[90] +matrix[91][30] * vector[91] +matrix[92][30] * vector[92] +matrix[93][30] * vector[93] +matrix[94][30] * vector[94] +matrix[95][30] * vector[95] +matrix[96][30] * vector[96] +matrix[97][30] * vector[97] +matrix[98][30] * vector[98] +matrix[99][30] * vector[99] +b[30];
assign result[31] = matrix[0][31] * vector[0] +matrix[1][31] * vector[1] +matrix[2][31] * vector[2] +matrix[3][31] * vector[3] +matrix[4][31] * vector[4] +matrix[5][31] * vector[5] +matrix[6][31] * vector[6] +matrix[7][31] * vector[7] +matrix[8][31] * vector[8] +matrix[9][31] * vector[9] +matrix[10][31] * vector[10] +matrix[11][31] * vector[11] +matrix[12][31] * vector[12] +matrix[13][31] * vector[13] +matrix[14][31] * vector[14] +matrix[15][31] * vector[15] +matrix[16][31] * vector[16] +matrix[17][31] * vector[17] +matrix[18][31] * vector[18] +matrix[19][31] * vector[19] +matrix[20][31] * vector[20] +matrix[21][31] * vector[21] +matrix[22][31] * vector[22] +matrix[23][31] * vector[23] +matrix[24][31] * vector[24] +matrix[25][31] * vector[25] +matrix[26][31] * vector[26] +matrix[27][31] * vector[27] +matrix[28][31] * vector[28] +matrix[29][31] * vector[29] +matrix[30][31] * vector[30] +matrix[31][31] * vector[31] +matrix[32][31] * vector[32] +matrix[33][31] * vector[33] +matrix[34][31] * vector[34] +matrix[35][31] * vector[35] +matrix[36][31] * vector[36] +matrix[37][31] * vector[37] +matrix[38][31] * vector[38] +matrix[39][31] * vector[39] +matrix[40][31] * vector[40] +matrix[41][31] * vector[41] +matrix[42][31] * vector[42] +matrix[43][31] * vector[43] +matrix[44][31] * vector[44] +matrix[45][31] * vector[45] +matrix[46][31] * vector[46] +matrix[47][31] * vector[47] +matrix[48][31] * vector[48] +matrix[49][31] * vector[49] +matrix[50][31] * vector[50] +matrix[51][31] * vector[51] +matrix[52][31] * vector[52] +matrix[53][31] * vector[53] +matrix[54][31] * vector[54] +matrix[55][31] * vector[55] +matrix[56][31] * vector[56] +matrix[57][31] * vector[57] +matrix[58][31] * vector[58] +matrix[59][31] * vector[59] +matrix[60][31] * vector[60] +matrix[61][31] * vector[61] +matrix[62][31] * vector[62] +matrix[63][31] * vector[63] +matrix[64][31] * vector[64] +matrix[65][31] * vector[65] +matrix[66][31] * vector[66] +matrix[67][31] * vector[67] +matrix[68][31] * vector[68] +matrix[69][31] * vector[69] +matrix[70][31] * vector[70] +matrix[71][31] * vector[71] +matrix[72][31] * vector[72] +matrix[73][31] * vector[73] +matrix[74][31] * vector[74] +matrix[75][31] * vector[75] +matrix[76][31] * vector[76] +matrix[77][31] * vector[77] +matrix[78][31] * vector[78] +matrix[79][31] * vector[79] +matrix[80][31] * vector[80] +matrix[81][31] * vector[81] +matrix[82][31] * vector[82] +matrix[83][31] * vector[83] +matrix[84][31] * vector[84] +matrix[85][31] * vector[85] +matrix[86][31] * vector[86] +matrix[87][31] * vector[87] +matrix[88][31] * vector[88] +matrix[89][31] * vector[89] +matrix[90][31] * vector[90] +matrix[91][31] * vector[91] +matrix[92][31] * vector[92] +matrix[93][31] * vector[93] +matrix[94][31] * vector[94] +matrix[95][31] * vector[95] +matrix[96][31] * vector[96] +matrix[97][31] * vector[97] +matrix[98][31] * vector[98] +matrix[99][31] * vector[99] +b[31];
assign result[32] = matrix[0][32] * vector[0] +matrix[1][32] * vector[1] +matrix[2][32] * vector[2] +matrix[3][32] * vector[3] +matrix[4][32] * vector[4] +matrix[5][32] * vector[5] +matrix[6][32] * vector[6] +matrix[7][32] * vector[7] +matrix[8][32] * vector[8] +matrix[9][32] * vector[9] +matrix[10][32] * vector[10] +matrix[11][32] * vector[11] +matrix[12][32] * vector[12] +matrix[13][32] * vector[13] +matrix[14][32] * vector[14] +matrix[15][32] * vector[15] +matrix[16][32] * vector[16] +matrix[17][32] * vector[17] +matrix[18][32] * vector[18] +matrix[19][32] * vector[19] +matrix[20][32] * vector[20] +matrix[21][32] * vector[21] +matrix[22][32] * vector[22] +matrix[23][32] * vector[23] +matrix[24][32] * vector[24] +matrix[25][32] * vector[25] +matrix[26][32] * vector[26] +matrix[27][32] * vector[27] +matrix[28][32] * vector[28] +matrix[29][32] * vector[29] +matrix[30][32] * vector[30] +matrix[31][32] * vector[31] +matrix[32][32] * vector[32] +matrix[33][32] * vector[33] +matrix[34][32] * vector[34] +matrix[35][32] * vector[35] +matrix[36][32] * vector[36] +matrix[37][32] * vector[37] +matrix[38][32] * vector[38] +matrix[39][32] * vector[39] +matrix[40][32] * vector[40] +matrix[41][32] * vector[41] +matrix[42][32] * vector[42] +matrix[43][32] * vector[43] +matrix[44][32] * vector[44] +matrix[45][32] * vector[45] +matrix[46][32] * vector[46] +matrix[47][32] * vector[47] +matrix[48][32] * vector[48] +matrix[49][32] * vector[49] +matrix[50][32] * vector[50] +matrix[51][32] * vector[51] +matrix[52][32] * vector[52] +matrix[53][32] * vector[53] +matrix[54][32] * vector[54] +matrix[55][32] * vector[55] +matrix[56][32] * vector[56] +matrix[57][32] * vector[57] +matrix[58][32] * vector[58] +matrix[59][32] * vector[59] +matrix[60][32] * vector[60] +matrix[61][32] * vector[61] +matrix[62][32] * vector[62] +matrix[63][32] * vector[63] +matrix[64][32] * vector[64] +matrix[65][32] * vector[65] +matrix[66][32] * vector[66] +matrix[67][32] * vector[67] +matrix[68][32] * vector[68] +matrix[69][32] * vector[69] +matrix[70][32] * vector[70] +matrix[71][32] * vector[71] +matrix[72][32] * vector[72] +matrix[73][32] * vector[73] +matrix[74][32] * vector[74] +matrix[75][32] * vector[75] +matrix[76][32] * vector[76] +matrix[77][32] * vector[77] +matrix[78][32] * vector[78] +matrix[79][32] * vector[79] +matrix[80][32] * vector[80] +matrix[81][32] * vector[81] +matrix[82][32] * vector[82] +matrix[83][32] * vector[83] +matrix[84][32] * vector[84] +matrix[85][32] * vector[85] +matrix[86][32] * vector[86] +matrix[87][32] * vector[87] +matrix[88][32] * vector[88] +matrix[89][32] * vector[89] +matrix[90][32] * vector[90] +matrix[91][32] * vector[91] +matrix[92][32] * vector[92] +matrix[93][32] * vector[93] +matrix[94][32] * vector[94] +matrix[95][32] * vector[95] +matrix[96][32] * vector[96] +matrix[97][32] * vector[97] +matrix[98][32] * vector[98] +matrix[99][32] * vector[99] +b[32];
assign result[33] = matrix[0][33] * vector[0] +matrix[1][33] * vector[1] +matrix[2][33] * vector[2] +matrix[3][33] * vector[3] +matrix[4][33] * vector[4] +matrix[5][33] * vector[5] +matrix[6][33] * vector[6] +matrix[7][33] * vector[7] +matrix[8][33] * vector[8] +matrix[9][33] * vector[9] +matrix[10][33] * vector[10] +matrix[11][33] * vector[11] +matrix[12][33] * vector[12] +matrix[13][33] * vector[13] +matrix[14][33] * vector[14] +matrix[15][33] * vector[15] +matrix[16][33] * vector[16] +matrix[17][33] * vector[17] +matrix[18][33] * vector[18] +matrix[19][33] * vector[19] +matrix[20][33] * vector[20] +matrix[21][33] * vector[21] +matrix[22][33] * vector[22] +matrix[23][33] * vector[23] +matrix[24][33] * vector[24] +matrix[25][33] * vector[25] +matrix[26][33] * vector[26] +matrix[27][33] * vector[27] +matrix[28][33] * vector[28] +matrix[29][33] * vector[29] +matrix[30][33] * vector[30] +matrix[31][33] * vector[31] +matrix[32][33] * vector[32] +matrix[33][33] * vector[33] +matrix[34][33] * vector[34] +matrix[35][33] * vector[35] +matrix[36][33] * vector[36] +matrix[37][33] * vector[37] +matrix[38][33] * vector[38] +matrix[39][33] * vector[39] +matrix[40][33] * vector[40] +matrix[41][33] * vector[41] +matrix[42][33] * vector[42] +matrix[43][33] * vector[43] +matrix[44][33] * vector[44] +matrix[45][33] * vector[45] +matrix[46][33] * vector[46] +matrix[47][33] * vector[47] +matrix[48][33] * vector[48] +matrix[49][33] * vector[49] +matrix[50][33] * vector[50] +matrix[51][33] * vector[51] +matrix[52][33] * vector[52] +matrix[53][33] * vector[53] +matrix[54][33] * vector[54] +matrix[55][33] * vector[55] +matrix[56][33] * vector[56] +matrix[57][33] * vector[57] +matrix[58][33] * vector[58] +matrix[59][33] * vector[59] +matrix[60][33] * vector[60] +matrix[61][33] * vector[61] +matrix[62][33] * vector[62] +matrix[63][33] * vector[63] +matrix[64][33] * vector[64] +matrix[65][33] * vector[65] +matrix[66][33] * vector[66] +matrix[67][33] * vector[67] +matrix[68][33] * vector[68] +matrix[69][33] * vector[69] +matrix[70][33] * vector[70] +matrix[71][33] * vector[71] +matrix[72][33] * vector[72] +matrix[73][33] * vector[73] +matrix[74][33] * vector[74] +matrix[75][33] * vector[75] +matrix[76][33] * vector[76] +matrix[77][33] * vector[77] +matrix[78][33] * vector[78] +matrix[79][33] * vector[79] +matrix[80][33] * vector[80] +matrix[81][33] * vector[81] +matrix[82][33] * vector[82] +matrix[83][33] * vector[83] +matrix[84][33] * vector[84] +matrix[85][33] * vector[85] +matrix[86][33] * vector[86] +matrix[87][33] * vector[87] +matrix[88][33] * vector[88] +matrix[89][33] * vector[89] +matrix[90][33] * vector[90] +matrix[91][33] * vector[91] +matrix[92][33] * vector[92] +matrix[93][33] * vector[93] +matrix[94][33] * vector[94] +matrix[95][33] * vector[95] +matrix[96][33] * vector[96] +matrix[97][33] * vector[97] +matrix[98][33] * vector[98] +matrix[99][33] * vector[99] +b[33];
assign result[34] = matrix[0][34] * vector[0] +matrix[1][34] * vector[1] +matrix[2][34] * vector[2] +matrix[3][34] * vector[3] +matrix[4][34] * vector[4] +matrix[5][34] * vector[5] +matrix[6][34] * vector[6] +matrix[7][34] * vector[7] +matrix[8][34] * vector[8] +matrix[9][34] * vector[9] +matrix[10][34] * vector[10] +matrix[11][34] * vector[11] +matrix[12][34] * vector[12] +matrix[13][34] * vector[13] +matrix[14][34] * vector[14] +matrix[15][34] * vector[15] +matrix[16][34] * vector[16] +matrix[17][34] * vector[17] +matrix[18][34] * vector[18] +matrix[19][34] * vector[19] +matrix[20][34] * vector[20] +matrix[21][34] * vector[21] +matrix[22][34] * vector[22] +matrix[23][34] * vector[23] +matrix[24][34] * vector[24] +matrix[25][34] * vector[25] +matrix[26][34] * vector[26] +matrix[27][34] * vector[27] +matrix[28][34] * vector[28] +matrix[29][34] * vector[29] +matrix[30][34] * vector[30] +matrix[31][34] * vector[31] +matrix[32][34] * vector[32] +matrix[33][34] * vector[33] +matrix[34][34] * vector[34] +matrix[35][34] * vector[35] +matrix[36][34] * vector[36] +matrix[37][34] * vector[37] +matrix[38][34] * vector[38] +matrix[39][34] * vector[39] +matrix[40][34] * vector[40] +matrix[41][34] * vector[41] +matrix[42][34] * vector[42] +matrix[43][34] * vector[43] +matrix[44][34] * vector[44] +matrix[45][34] * vector[45] +matrix[46][34] * vector[46] +matrix[47][34] * vector[47] +matrix[48][34] * vector[48] +matrix[49][34] * vector[49] +matrix[50][34] * vector[50] +matrix[51][34] * vector[51] +matrix[52][34] * vector[52] +matrix[53][34] * vector[53] +matrix[54][34] * vector[54] +matrix[55][34] * vector[55] +matrix[56][34] * vector[56] +matrix[57][34] * vector[57] +matrix[58][34] * vector[58] +matrix[59][34] * vector[59] +matrix[60][34] * vector[60] +matrix[61][34] * vector[61] +matrix[62][34] * vector[62] +matrix[63][34] * vector[63] +matrix[64][34] * vector[64] +matrix[65][34] * vector[65] +matrix[66][34] * vector[66] +matrix[67][34] * vector[67] +matrix[68][34] * vector[68] +matrix[69][34] * vector[69] +matrix[70][34] * vector[70] +matrix[71][34] * vector[71] +matrix[72][34] * vector[72] +matrix[73][34] * vector[73] +matrix[74][34] * vector[74] +matrix[75][34] * vector[75] +matrix[76][34] * vector[76] +matrix[77][34] * vector[77] +matrix[78][34] * vector[78] +matrix[79][34] * vector[79] +matrix[80][34] * vector[80] +matrix[81][34] * vector[81] +matrix[82][34] * vector[82] +matrix[83][34] * vector[83] +matrix[84][34] * vector[84] +matrix[85][34] * vector[85] +matrix[86][34] * vector[86] +matrix[87][34] * vector[87] +matrix[88][34] * vector[88] +matrix[89][34] * vector[89] +matrix[90][34] * vector[90] +matrix[91][34] * vector[91] +matrix[92][34] * vector[92] +matrix[93][34] * vector[93] +matrix[94][34] * vector[94] +matrix[95][34] * vector[95] +matrix[96][34] * vector[96] +matrix[97][34] * vector[97] +matrix[98][34] * vector[98] +matrix[99][34] * vector[99] +b[34];
assign result[35] = matrix[0][35] * vector[0] +matrix[1][35] * vector[1] +matrix[2][35] * vector[2] +matrix[3][35] * vector[3] +matrix[4][35] * vector[4] +matrix[5][35] * vector[5] +matrix[6][35] * vector[6] +matrix[7][35] * vector[7] +matrix[8][35] * vector[8] +matrix[9][35] * vector[9] +matrix[10][35] * vector[10] +matrix[11][35] * vector[11] +matrix[12][35] * vector[12] +matrix[13][35] * vector[13] +matrix[14][35] * vector[14] +matrix[15][35] * vector[15] +matrix[16][35] * vector[16] +matrix[17][35] * vector[17] +matrix[18][35] * vector[18] +matrix[19][35] * vector[19] +matrix[20][35] * vector[20] +matrix[21][35] * vector[21] +matrix[22][35] * vector[22] +matrix[23][35] * vector[23] +matrix[24][35] * vector[24] +matrix[25][35] * vector[25] +matrix[26][35] * vector[26] +matrix[27][35] * vector[27] +matrix[28][35] * vector[28] +matrix[29][35] * vector[29] +matrix[30][35] * vector[30] +matrix[31][35] * vector[31] +matrix[32][35] * vector[32] +matrix[33][35] * vector[33] +matrix[34][35] * vector[34] +matrix[35][35] * vector[35] +matrix[36][35] * vector[36] +matrix[37][35] * vector[37] +matrix[38][35] * vector[38] +matrix[39][35] * vector[39] +matrix[40][35] * vector[40] +matrix[41][35] * vector[41] +matrix[42][35] * vector[42] +matrix[43][35] * vector[43] +matrix[44][35] * vector[44] +matrix[45][35] * vector[45] +matrix[46][35] * vector[46] +matrix[47][35] * vector[47] +matrix[48][35] * vector[48] +matrix[49][35] * vector[49] +matrix[50][35] * vector[50] +matrix[51][35] * vector[51] +matrix[52][35] * vector[52] +matrix[53][35] * vector[53] +matrix[54][35] * vector[54] +matrix[55][35] * vector[55] +matrix[56][35] * vector[56] +matrix[57][35] * vector[57] +matrix[58][35] * vector[58] +matrix[59][35] * vector[59] +matrix[60][35] * vector[60] +matrix[61][35] * vector[61] +matrix[62][35] * vector[62] +matrix[63][35] * vector[63] +matrix[64][35] * vector[64] +matrix[65][35] * vector[65] +matrix[66][35] * vector[66] +matrix[67][35] * vector[67] +matrix[68][35] * vector[68] +matrix[69][35] * vector[69] +matrix[70][35] * vector[70] +matrix[71][35] * vector[71] +matrix[72][35] * vector[72] +matrix[73][35] * vector[73] +matrix[74][35] * vector[74] +matrix[75][35] * vector[75] +matrix[76][35] * vector[76] +matrix[77][35] * vector[77] +matrix[78][35] * vector[78] +matrix[79][35] * vector[79] +matrix[80][35] * vector[80] +matrix[81][35] * vector[81] +matrix[82][35] * vector[82] +matrix[83][35] * vector[83] +matrix[84][35] * vector[84] +matrix[85][35] * vector[85] +matrix[86][35] * vector[86] +matrix[87][35] * vector[87] +matrix[88][35] * vector[88] +matrix[89][35] * vector[89] +matrix[90][35] * vector[90] +matrix[91][35] * vector[91] +matrix[92][35] * vector[92] +matrix[93][35] * vector[93] +matrix[94][35] * vector[94] +matrix[95][35] * vector[95] +matrix[96][35] * vector[96] +matrix[97][35] * vector[97] +matrix[98][35] * vector[98] +matrix[99][35] * vector[99] +b[35];
assign result[36] = matrix[0][36] * vector[0] +matrix[1][36] * vector[1] +matrix[2][36] * vector[2] +matrix[3][36] * vector[3] +matrix[4][36] * vector[4] +matrix[5][36] * vector[5] +matrix[6][36] * vector[6] +matrix[7][36] * vector[7] +matrix[8][36] * vector[8] +matrix[9][36] * vector[9] +matrix[10][36] * vector[10] +matrix[11][36] * vector[11] +matrix[12][36] * vector[12] +matrix[13][36] * vector[13] +matrix[14][36] * vector[14] +matrix[15][36] * vector[15] +matrix[16][36] * vector[16] +matrix[17][36] * vector[17] +matrix[18][36] * vector[18] +matrix[19][36] * vector[19] +matrix[20][36] * vector[20] +matrix[21][36] * vector[21] +matrix[22][36] * vector[22] +matrix[23][36] * vector[23] +matrix[24][36] * vector[24] +matrix[25][36] * vector[25] +matrix[26][36] * vector[26] +matrix[27][36] * vector[27] +matrix[28][36] * vector[28] +matrix[29][36] * vector[29] +matrix[30][36] * vector[30] +matrix[31][36] * vector[31] +matrix[32][36] * vector[32] +matrix[33][36] * vector[33] +matrix[34][36] * vector[34] +matrix[35][36] * vector[35] +matrix[36][36] * vector[36] +matrix[37][36] * vector[37] +matrix[38][36] * vector[38] +matrix[39][36] * vector[39] +matrix[40][36] * vector[40] +matrix[41][36] * vector[41] +matrix[42][36] * vector[42] +matrix[43][36] * vector[43] +matrix[44][36] * vector[44] +matrix[45][36] * vector[45] +matrix[46][36] * vector[46] +matrix[47][36] * vector[47] +matrix[48][36] * vector[48] +matrix[49][36] * vector[49] +matrix[50][36] * vector[50] +matrix[51][36] * vector[51] +matrix[52][36] * vector[52] +matrix[53][36] * vector[53] +matrix[54][36] * vector[54] +matrix[55][36] * vector[55] +matrix[56][36] * vector[56] +matrix[57][36] * vector[57] +matrix[58][36] * vector[58] +matrix[59][36] * vector[59] +matrix[60][36] * vector[60] +matrix[61][36] * vector[61] +matrix[62][36] * vector[62] +matrix[63][36] * vector[63] +matrix[64][36] * vector[64] +matrix[65][36] * vector[65] +matrix[66][36] * vector[66] +matrix[67][36] * vector[67] +matrix[68][36] * vector[68] +matrix[69][36] * vector[69] +matrix[70][36] * vector[70] +matrix[71][36] * vector[71] +matrix[72][36] * vector[72] +matrix[73][36] * vector[73] +matrix[74][36] * vector[74] +matrix[75][36] * vector[75] +matrix[76][36] * vector[76] +matrix[77][36] * vector[77] +matrix[78][36] * vector[78] +matrix[79][36] * vector[79] +matrix[80][36] * vector[80] +matrix[81][36] * vector[81] +matrix[82][36] * vector[82] +matrix[83][36] * vector[83] +matrix[84][36] * vector[84] +matrix[85][36] * vector[85] +matrix[86][36] * vector[86] +matrix[87][36] * vector[87] +matrix[88][36] * vector[88] +matrix[89][36] * vector[89] +matrix[90][36] * vector[90] +matrix[91][36] * vector[91] +matrix[92][36] * vector[92] +matrix[93][36] * vector[93] +matrix[94][36] * vector[94] +matrix[95][36] * vector[95] +matrix[96][36] * vector[96] +matrix[97][36] * vector[97] +matrix[98][36] * vector[98] +matrix[99][36] * vector[99] +b[36];
assign result[37] = matrix[0][37] * vector[0] +matrix[1][37] * vector[1] +matrix[2][37] * vector[2] +matrix[3][37] * vector[3] +matrix[4][37] * vector[4] +matrix[5][37] * vector[5] +matrix[6][37] * vector[6] +matrix[7][37] * vector[7] +matrix[8][37] * vector[8] +matrix[9][37] * vector[9] +matrix[10][37] * vector[10] +matrix[11][37] * vector[11] +matrix[12][37] * vector[12] +matrix[13][37] * vector[13] +matrix[14][37] * vector[14] +matrix[15][37] * vector[15] +matrix[16][37] * vector[16] +matrix[17][37] * vector[17] +matrix[18][37] * vector[18] +matrix[19][37] * vector[19] +matrix[20][37] * vector[20] +matrix[21][37] * vector[21] +matrix[22][37] * vector[22] +matrix[23][37] * vector[23] +matrix[24][37] * vector[24] +matrix[25][37] * vector[25] +matrix[26][37] * vector[26] +matrix[27][37] * vector[27] +matrix[28][37] * vector[28] +matrix[29][37] * vector[29] +matrix[30][37] * vector[30] +matrix[31][37] * vector[31] +matrix[32][37] * vector[32] +matrix[33][37] * vector[33] +matrix[34][37] * vector[34] +matrix[35][37] * vector[35] +matrix[36][37] * vector[36] +matrix[37][37] * vector[37] +matrix[38][37] * vector[38] +matrix[39][37] * vector[39] +matrix[40][37] * vector[40] +matrix[41][37] * vector[41] +matrix[42][37] * vector[42] +matrix[43][37] * vector[43] +matrix[44][37] * vector[44] +matrix[45][37] * vector[45] +matrix[46][37] * vector[46] +matrix[47][37] * vector[47] +matrix[48][37] * vector[48] +matrix[49][37] * vector[49] +matrix[50][37] * vector[50] +matrix[51][37] * vector[51] +matrix[52][37] * vector[52] +matrix[53][37] * vector[53] +matrix[54][37] * vector[54] +matrix[55][37] * vector[55] +matrix[56][37] * vector[56] +matrix[57][37] * vector[57] +matrix[58][37] * vector[58] +matrix[59][37] * vector[59] +matrix[60][37] * vector[60] +matrix[61][37] * vector[61] +matrix[62][37] * vector[62] +matrix[63][37] * vector[63] +matrix[64][37] * vector[64] +matrix[65][37] * vector[65] +matrix[66][37] * vector[66] +matrix[67][37] * vector[67] +matrix[68][37] * vector[68] +matrix[69][37] * vector[69] +matrix[70][37] * vector[70] +matrix[71][37] * vector[71] +matrix[72][37] * vector[72] +matrix[73][37] * vector[73] +matrix[74][37] * vector[74] +matrix[75][37] * vector[75] +matrix[76][37] * vector[76] +matrix[77][37] * vector[77] +matrix[78][37] * vector[78] +matrix[79][37] * vector[79] +matrix[80][37] * vector[80] +matrix[81][37] * vector[81] +matrix[82][37] * vector[82] +matrix[83][37] * vector[83] +matrix[84][37] * vector[84] +matrix[85][37] * vector[85] +matrix[86][37] * vector[86] +matrix[87][37] * vector[87] +matrix[88][37] * vector[88] +matrix[89][37] * vector[89] +matrix[90][37] * vector[90] +matrix[91][37] * vector[91] +matrix[92][37] * vector[92] +matrix[93][37] * vector[93] +matrix[94][37] * vector[94] +matrix[95][37] * vector[95] +matrix[96][37] * vector[96] +matrix[97][37] * vector[97] +matrix[98][37] * vector[98] +matrix[99][37] * vector[99] +b[37];
assign result[38] = matrix[0][38] * vector[0] +matrix[1][38] * vector[1] +matrix[2][38] * vector[2] +matrix[3][38] * vector[3] +matrix[4][38] * vector[4] +matrix[5][38] * vector[5] +matrix[6][38] * vector[6] +matrix[7][38] * vector[7] +matrix[8][38] * vector[8] +matrix[9][38] * vector[9] +matrix[10][38] * vector[10] +matrix[11][38] * vector[11] +matrix[12][38] * vector[12] +matrix[13][38] * vector[13] +matrix[14][38] * vector[14] +matrix[15][38] * vector[15] +matrix[16][38] * vector[16] +matrix[17][38] * vector[17] +matrix[18][38] * vector[18] +matrix[19][38] * vector[19] +matrix[20][38] * vector[20] +matrix[21][38] * vector[21] +matrix[22][38] * vector[22] +matrix[23][38] * vector[23] +matrix[24][38] * vector[24] +matrix[25][38] * vector[25] +matrix[26][38] * vector[26] +matrix[27][38] * vector[27] +matrix[28][38] * vector[28] +matrix[29][38] * vector[29] +matrix[30][38] * vector[30] +matrix[31][38] * vector[31] +matrix[32][38] * vector[32] +matrix[33][38] * vector[33] +matrix[34][38] * vector[34] +matrix[35][38] * vector[35] +matrix[36][38] * vector[36] +matrix[37][38] * vector[37] +matrix[38][38] * vector[38] +matrix[39][38] * vector[39] +matrix[40][38] * vector[40] +matrix[41][38] * vector[41] +matrix[42][38] * vector[42] +matrix[43][38] * vector[43] +matrix[44][38] * vector[44] +matrix[45][38] * vector[45] +matrix[46][38] * vector[46] +matrix[47][38] * vector[47] +matrix[48][38] * vector[48] +matrix[49][38] * vector[49] +matrix[50][38] * vector[50] +matrix[51][38] * vector[51] +matrix[52][38] * vector[52] +matrix[53][38] * vector[53] +matrix[54][38] * vector[54] +matrix[55][38] * vector[55] +matrix[56][38] * vector[56] +matrix[57][38] * vector[57] +matrix[58][38] * vector[58] +matrix[59][38] * vector[59] +matrix[60][38] * vector[60] +matrix[61][38] * vector[61] +matrix[62][38] * vector[62] +matrix[63][38] * vector[63] +matrix[64][38] * vector[64] +matrix[65][38] * vector[65] +matrix[66][38] * vector[66] +matrix[67][38] * vector[67] +matrix[68][38] * vector[68] +matrix[69][38] * vector[69] +matrix[70][38] * vector[70] +matrix[71][38] * vector[71] +matrix[72][38] * vector[72] +matrix[73][38] * vector[73] +matrix[74][38] * vector[74] +matrix[75][38] * vector[75] +matrix[76][38] * vector[76] +matrix[77][38] * vector[77] +matrix[78][38] * vector[78] +matrix[79][38] * vector[79] +matrix[80][38] * vector[80] +matrix[81][38] * vector[81] +matrix[82][38] * vector[82] +matrix[83][38] * vector[83] +matrix[84][38] * vector[84] +matrix[85][38] * vector[85] +matrix[86][38] * vector[86] +matrix[87][38] * vector[87] +matrix[88][38] * vector[88] +matrix[89][38] * vector[89] +matrix[90][38] * vector[90] +matrix[91][38] * vector[91] +matrix[92][38] * vector[92] +matrix[93][38] * vector[93] +matrix[94][38] * vector[94] +matrix[95][38] * vector[95] +matrix[96][38] * vector[96] +matrix[97][38] * vector[97] +matrix[98][38] * vector[98] +matrix[99][38] * vector[99] +b[38];
assign result[39] = matrix[0][39] * vector[0] +matrix[1][39] * vector[1] +matrix[2][39] * vector[2] +matrix[3][39] * vector[3] +matrix[4][39] * vector[4] +matrix[5][39] * vector[5] +matrix[6][39] * vector[6] +matrix[7][39] * vector[7] +matrix[8][39] * vector[8] +matrix[9][39] * vector[9] +matrix[10][39] * vector[10] +matrix[11][39] * vector[11] +matrix[12][39] * vector[12] +matrix[13][39] * vector[13] +matrix[14][39] * vector[14] +matrix[15][39] * vector[15] +matrix[16][39] * vector[16] +matrix[17][39] * vector[17] +matrix[18][39] * vector[18] +matrix[19][39] * vector[19] +matrix[20][39] * vector[20] +matrix[21][39] * vector[21] +matrix[22][39] * vector[22] +matrix[23][39] * vector[23] +matrix[24][39] * vector[24] +matrix[25][39] * vector[25] +matrix[26][39] * vector[26] +matrix[27][39] * vector[27] +matrix[28][39] * vector[28] +matrix[29][39] * vector[29] +matrix[30][39] * vector[30] +matrix[31][39] * vector[31] +matrix[32][39] * vector[32] +matrix[33][39] * vector[33] +matrix[34][39] * vector[34] +matrix[35][39] * vector[35] +matrix[36][39] * vector[36] +matrix[37][39] * vector[37] +matrix[38][39] * vector[38] +matrix[39][39] * vector[39] +matrix[40][39] * vector[40] +matrix[41][39] * vector[41] +matrix[42][39] * vector[42] +matrix[43][39] * vector[43] +matrix[44][39] * vector[44] +matrix[45][39] * vector[45] +matrix[46][39] * vector[46] +matrix[47][39] * vector[47] +matrix[48][39] * vector[48] +matrix[49][39] * vector[49] +matrix[50][39] * vector[50] +matrix[51][39] * vector[51] +matrix[52][39] * vector[52] +matrix[53][39] * vector[53] +matrix[54][39] * vector[54] +matrix[55][39] * vector[55] +matrix[56][39] * vector[56] +matrix[57][39] * vector[57] +matrix[58][39] * vector[58] +matrix[59][39] * vector[59] +matrix[60][39] * vector[60] +matrix[61][39] * vector[61] +matrix[62][39] * vector[62] +matrix[63][39] * vector[63] +matrix[64][39] * vector[64] +matrix[65][39] * vector[65] +matrix[66][39] * vector[66] +matrix[67][39] * vector[67] +matrix[68][39] * vector[68] +matrix[69][39] * vector[69] +matrix[70][39] * vector[70] +matrix[71][39] * vector[71] +matrix[72][39] * vector[72] +matrix[73][39] * vector[73] +matrix[74][39] * vector[74] +matrix[75][39] * vector[75] +matrix[76][39] * vector[76] +matrix[77][39] * vector[77] +matrix[78][39] * vector[78] +matrix[79][39] * vector[79] +matrix[80][39] * vector[80] +matrix[81][39] * vector[81] +matrix[82][39] * vector[82] +matrix[83][39] * vector[83] +matrix[84][39] * vector[84] +matrix[85][39] * vector[85] +matrix[86][39] * vector[86] +matrix[87][39] * vector[87] +matrix[88][39] * vector[88] +matrix[89][39] * vector[89] +matrix[90][39] * vector[90] +matrix[91][39] * vector[91] +matrix[92][39] * vector[92] +matrix[93][39] * vector[93] +matrix[94][39] * vector[94] +matrix[95][39] * vector[95] +matrix[96][39] * vector[96] +matrix[97][39] * vector[97] +matrix[98][39] * vector[98] +matrix[99][39] * vector[99] +b[39];
assign result[40] = matrix[0][40] * vector[0] +matrix[1][40] * vector[1] +matrix[2][40] * vector[2] +matrix[3][40] * vector[3] +matrix[4][40] * vector[4] +matrix[5][40] * vector[5] +matrix[6][40] * vector[6] +matrix[7][40] * vector[7] +matrix[8][40] * vector[8] +matrix[9][40] * vector[9] +matrix[10][40] * vector[10] +matrix[11][40] * vector[11] +matrix[12][40] * vector[12] +matrix[13][40] * vector[13] +matrix[14][40] * vector[14] +matrix[15][40] * vector[15] +matrix[16][40] * vector[16] +matrix[17][40] * vector[17] +matrix[18][40] * vector[18] +matrix[19][40] * vector[19] +matrix[20][40] * vector[20] +matrix[21][40] * vector[21] +matrix[22][40] * vector[22] +matrix[23][40] * vector[23] +matrix[24][40] * vector[24] +matrix[25][40] * vector[25] +matrix[26][40] * vector[26] +matrix[27][40] * vector[27] +matrix[28][40] * vector[28] +matrix[29][40] * vector[29] +matrix[30][40] * vector[30] +matrix[31][40] * vector[31] +matrix[32][40] * vector[32] +matrix[33][40] * vector[33] +matrix[34][40] * vector[34] +matrix[35][40] * vector[35] +matrix[36][40] * vector[36] +matrix[37][40] * vector[37] +matrix[38][40] * vector[38] +matrix[39][40] * vector[39] +matrix[40][40] * vector[40] +matrix[41][40] * vector[41] +matrix[42][40] * vector[42] +matrix[43][40] * vector[43] +matrix[44][40] * vector[44] +matrix[45][40] * vector[45] +matrix[46][40] * vector[46] +matrix[47][40] * vector[47] +matrix[48][40] * vector[48] +matrix[49][40] * vector[49] +matrix[50][40] * vector[50] +matrix[51][40] * vector[51] +matrix[52][40] * vector[52] +matrix[53][40] * vector[53] +matrix[54][40] * vector[54] +matrix[55][40] * vector[55] +matrix[56][40] * vector[56] +matrix[57][40] * vector[57] +matrix[58][40] * vector[58] +matrix[59][40] * vector[59] +matrix[60][40] * vector[60] +matrix[61][40] * vector[61] +matrix[62][40] * vector[62] +matrix[63][40] * vector[63] +matrix[64][40] * vector[64] +matrix[65][40] * vector[65] +matrix[66][40] * vector[66] +matrix[67][40] * vector[67] +matrix[68][40] * vector[68] +matrix[69][40] * vector[69] +matrix[70][40] * vector[70] +matrix[71][40] * vector[71] +matrix[72][40] * vector[72] +matrix[73][40] * vector[73] +matrix[74][40] * vector[74] +matrix[75][40] * vector[75] +matrix[76][40] * vector[76] +matrix[77][40] * vector[77] +matrix[78][40] * vector[78] +matrix[79][40] * vector[79] +matrix[80][40] * vector[80] +matrix[81][40] * vector[81] +matrix[82][40] * vector[82] +matrix[83][40] * vector[83] +matrix[84][40] * vector[84] +matrix[85][40] * vector[85] +matrix[86][40] * vector[86] +matrix[87][40] * vector[87] +matrix[88][40] * vector[88] +matrix[89][40] * vector[89] +matrix[90][40] * vector[90] +matrix[91][40] * vector[91] +matrix[92][40] * vector[92] +matrix[93][40] * vector[93] +matrix[94][40] * vector[94] +matrix[95][40] * vector[95] +matrix[96][40] * vector[96] +matrix[97][40] * vector[97] +matrix[98][40] * vector[98] +matrix[99][40] * vector[99] +b[40];
assign result[41] = matrix[0][41] * vector[0] +matrix[1][41] * vector[1] +matrix[2][41] * vector[2] +matrix[3][41] * vector[3] +matrix[4][41] * vector[4] +matrix[5][41] * vector[5] +matrix[6][41] * vector[6] +matrix[7][41] * vector[7] +matrix[8][41] * vector[8] +matrix[9][41] * vector[9] +matrix[10][41] * vector[10] +matrix[11][41] * vector[11] +matrix[12][41] * vector[12] +matrix[13][41] * vector[13] +matrix[14][41] * vector[14] +matrix[15][41] * vector[15] +matrix[16][41] * vector[16] +matrix[17][41] * vector[17] +matrix[18][41] * vector[18] +matrix[19][41] * vector[19] +matrix[20][41] * vector[20] +matrix[21][41] * vector[21] +matrix[22][41] * vector[22] +matrix[23][41] * vector[23] +matrix[24][41] * vector[24] +matrix[25][41] * vector[25] +matrix[26][41] * vector[26] +matrix[27][41] * vector[27] +matrix[28][41] * vector[28] +matrix[29][41] * vector[29] +matrix[30][41] * vector[30] +matrix[31][41] * vector[31] +matrix[32][41] * vector[32] +matrix[33][41] * vector[33] +matrix[34][41] * vector[34] +matrix[35][41] * vector[35] +matrix[36][41] * vector[36] +matrix[37][41] * vector[37] +matrix[38][41] * vector[38] +matrix[39][41] * vector[39] +matrix[40][41] * vector[40] +matrix[41][41] * vector[41] +matrix[42][41] * vector[42] +matrix[43][41] * vector[43] +matrix[44][41] * vector[44] +matrix[45][41] * vector[45] +matrix[46][41] * vector[46] +matrix[47][41] * vector[47] +matrix[48][41] * vector[48] +matrix[49][41] * vector[49] +matrix[50][41] * vector[50] +matrix[51][41] * vector[51] +matrix[52][41] * vector[52] +matrix[53][41] * vector[53] +matrix[54][41] * vector[54] +matrix[55][41] * vector[55] +matrix[56][41] * vector[56] +matrix[57][41] * vector[57] +matrix[58][41] * vector[58] +matrix[59][41] * vector[59] +matrix[60][41] * vector[60] +matrix[61][41] * vector[61] +matrix[62][41] * vector[62] +matrix[63][41] * vector[63] +matrix[64][41] * vector[64] +matrix[65][41] * vector[65] +matrix[66][41] * vector[66] +matrix[67][41] * vector[67] +matrix[68][41] * vector[68] +matrix[69][41] * vector[69] +matrix[70][41] * vector[70] +matrix[71][41] * vector[71] +matrix[72][41] * vector[72] +matrix[73][41] * vector[73] +matrix[74][41] * vector[74] +matrix[75][41] * vector[75] +matrix[76][41] * vector[76] +matrix[77][41] * vector[77] +matrix[78][41] * vector[78] +matrix[79][41] * vector[79] +matrix[80][41] * vector[80] +matrix[81][41] * vector[81] +matrix[82][41] * vector[82] +matrix[83][41] * vector[83] +matrix[84][41] * vector[84] +matrix[85][41] * vector[85] +matrix[86][41] * vector[86] +matrix[87][41] * vector[87] +matrix[88][41] * vector[88] +matrix[89][41] * vector[89] +matrix[90][41] * vector[90] +matrix[91][41] * vector[91] +matrix[92][41] * vector[92] +matrix[93][41] * vector[93] +matrix[94][41] * vector[94] +matrix[95][41] * vector[95] +matrix[96][41] * vector[96] +matrix[97][41] * vector[97] +matrix[98][41] * vector[98] +matrix[99][41] * vector[99] +b[41];
assign result[42] = matrix[0][42] * vector[0] +matrix[1][42] * vector[1] +matrix[2][42] * vector[2] +matrix[3][42] * vector[3] +matrix[4][42] * vector[4] +matrix[5][42] * vector[5] +matrix[6][42] * vector[6] +matrix[7][42] * vector[7] +matrix[8][42] * vector[8] +matrix[9][42] * vector[9] +matrix[10][42] * vector[10] +matrix[11][42] * vector[11] +matrix[12][42] * vector[12] +matrix[13][42] * vector[13] +matrix[14][42] * vector[14] +matrix[15][42] * vector[15] +matrix[16][42] * vector[16] +matrix[17][42] * vector[17] +matrix[18][42] * vector[18] +matrix[19][42] * vector[19] +matrix[20][42] * vector[20] +matrix[21][42] * vector[21] +matrix[22][42] * vector[22] +matrix[23][42] * vector[23] +matrix[24][42] * vector[24] +matrix[25][42] * vector[25] +matrix[26][42] * vector[26] +matrix[27][42] * vector[27] +matrix[28][42] * vector[28] +matrix[29][42] * vector[29] +matrix[30][42] * vector[30] +matrix[31][42] * vector[31] +matrix[32][42] * vector[32] +matrix[33][42] * vector[33] +matrix[34][42] * vector[34] +matrix[35][42] * vector[35] +matrix[36][42] * vector[36] +matrix[37][42] * vector[37] +matrix[38][42] * vector[38] +matrix[39][42] * vector[39] +matrix[40][42] * vector[40] +matrix[41][42] * vector[41] +matrix[42][42] * vector[42] +matrix[43][42] * vector[43] +matrix[44][42] * vector[44] +matrix[45][42] * vector[45] +matrix[46][42] * vector[46] +matrix[47][42] * vector[47] +matrix[48][42] * vector[48] +matrix[49][42] * vector[49] +matrix[50][42] * vector[50] +matrix[51][42] * vector[51] +matrix[52][42] * vector[52] +matrix[53][42] * vector[53] +matrix[54][42] * vector[54] +matrix[55][42] * vector[55] +matrix[56][42] * vector[56] +matrix[57][42] * vector[57] +matrix[58][42] * vector[58] +matrix[59][42] * vector[59] +matrix[60][42] * vector[60] +matrix[61][42] * vector[61] +matrix[62][42] * vector[62] +matrix[63][42] * vector[63] +matrix[64][42] * vector[64] +matrix[65][42] * vector[65] +matrix[66][42] * vector[66] +matrix[67][42] * vector[67] +matrix[68][42] * vector[68] +matrix[69][42] * vector[69] +matrix[70][42] * vector[70] +matrix[71][42] * vector[71] +matrix[72][42] * vector[72] +matrix[73][42] * vector[73] +matrix[74][42] * vector[74] +matrix[75][42] * vector[75] +matrix[76][42] * vector[76] +matrix[77][42] * vector[77] +matrix[78][42] * vector[78] +matrix[79][42] * vector[79] +matrix[80][42] * vector[80] +matrix[81][42] * vector[81] +matrix[82][42] * vector[82] +matrix[83][42] * vector[83] +matrix[84][42] * vector[84] +matrix[85][42] * vector[85] +matrix[86][42] * vector[86] +matrix[87][42] * vector[87] +matrix[88][42] * vector[88] +matrix[89][42] * vector[89] +matrix[90][42] * vector[90] +matrix[91][42] * vector[91] +matrix[92][42] * vector[92] +matrix[93][42] * vector[93] +matrix[94][42] * vector[94] +matrix[95][42] * vector[95] +matrix[96][42] * vector[96] +matrix[97][42] * vector[97] +matrix[98][42] * vector[98] +matrix[99][42] * vector[99] +b[42];
assign result[43] = matrix[0][43] * vector[0] +matrix[1][43] * vector[1] +matrix[2][43] * vector[2] +matrix[3][43] * vector[3] +matrix[4][43] * vector[4] +matrix[5][43] * vector[5] +matrix[6][43] * vector[6] +matrix[7][43] * vector[7] +matrix[8][43] * vector[8] +matrix[9][43] * vector[9] +matrix[10][43] * vector[10] +matrix[11][43] * vector[11] +matrix[12][43] * vector[12] +matrix[13][43] * vector[13] +matrix[14][43] * vector[14] +matrix[15][43] * vector[15] +matrix[16][43] * vector[16] +matrix[17][43] * vector[17] +matrix[18][43] * vector[18] +matrix[19][43] * vector[19] +matrix[20][43] * vector[20] +matrix[21][43] * vector[21] +matrix[22][43] * vector[22] +matrix[23][43] * vector[23] +matrix[24][43] * vector[24] +matrix[25][43] * vector[25] +matrix[26][43] * vector[26] +matrix[27][43] * vector[27] +matrix[28][43] * vector[28] +matrix[29][43] * vector[29] +matrix[30][43] * vector[30] +matrix[31][43] * vector[31] +matrix[32][43] * vector[32] +matrix[33][43] * vector[33] +matrix[34][43] * vector[34] +matrix[35][43] * vector[35] +matrix[36][43] * vector[36] +matrix[37][43] * vector[37] +matrix[38][43] * vector[38] +matrix[39][43] * vector[39] +matrix[40][43] * vector[40] +matrix[41][43] * vector[41] +matrix[42][43] * vector[42] +matrix[43][43] * vector[43] +matrix[44][43] * vector[44] +matrix[45][43] * vector[45] +matrix[46][43] * vector[46] +matrix[47][43] * vector[47] +matrix[48][43] * vector[48] +matrix[49][43] * vector[49] +matrix[50][43] * vector[50] +matrix[51][43] * vector[51] +matrix[52][43] * vector[52] +matrix[53][43] * vector[53] +matrix[54][43] * vector[54] +matrix[55][43] * vector[55] +matrix[56][43] * vector[56] +matrix[57][43] * vector[57] +matrix[58][43] * vector[58] +matrix[59][43] * vector[59] +matrix[60][43] * vector[60] +matrix[61][43] * vector[61] +matrix[62][43] * vector[62] +matrix[63][43] * vector[63] +matrix[64][43] * vector[64] +matrix[65][43] * vector[65] +matrix[66][43] * vector[66] +matrix[67][43] * vector[67] +matrix[68][43] * vector[68] +matrix[69][43] * vector[69] +matrix[70][43] * vector[70] +matrix[71][43] * vector[71] +matrix[72][43] * vector[72] +matrix[73][43] * vector[73] +matrix[74][43] * vector[74] +matrix[75][43] * vector[75] +matrix[76][43] * vector[76] +matrix[77][43] * vector[77] +matrix[78][43] * vector[78] +matrix[79][43] * vector[79] +matrix[80][43] * vector[80] +matrix[81][43] * vector[81] +matrix[82][43] * vector[82] +matrix[83][43] * vector[83] +matrix[84][43] * vector[84] +matrix[85][43] * vector[85] +matrix[86][43] * vector[86] +matrix[87][43] * vector[87] +matrix[88][43] * vector[88] +matrix[89][43] * vector[89] +matrix[90][43] * vector[90] +matrix[91][43] * vector[91] +matrix[92][43] * vector[92] +matrix[93][43] * vector[93] +matrix[94][43] * vector[94] +matrix[95][43] * vector[95] +matrix[96][43] * vector[96] +matrix[97][43] * vector[97] +matrix[98][43] * vector[98] +matrix[99][43] * vector[99] +b[43];
assign result[44] = matrix[0][44] * vector[0] +matrix[1][44] * vector[1] +matrix[2][44] * vector[2] +matrix[3][44] * vector[3] +matrix[4][44] * vector[4] +matrix[5][44] * vector[5] +matrix[6][44] * vector[6] +matrix[7][44] * vector[7] +matrix[8][44] * vector[8] +matrix[9][44] * vector[9] +matrix[10][44] * vector[10] +matrix[11][44] * vector[11] +matrix[12][44] * vector[12] +matrix[13][44] * vector[13] +matrix[14][44] * vector[14] +matrix[15][44] * vector[15] +matrix[16][44] * vector[16] +matrix[17][44] * vector[17] +matrix[18][44] * vector[18] +matrix[19][44] * vector[19] +matrix[20][44] * vector[20] +matrix[21][44] * vector[21] +matrix[22][44] * vector[22] +matrix[23][44] * vector[23] +matrix[24][44] * vector[24] +matrix[25][44] * vector[25] +matrix[26][44] * vector[26] +matrix[27][44] * vector[27] +matrix[28][44] * vector[28] +matrix[29][44] * vector[29] +matrix[30][44] * vector[30] +matrix[31][44] * vector[31] +matrix[32][44] * vector[32] +matrix[33][44] * vector[33] +matrix[34][44] * vector[34] +matrix[35][44] * vector[35] +matrix[36][44] * vector[36] +matrix[37][44] * vector[37] +matrix[38][44] * vector[38] +matrix[39][44] * vector[39] +matrix[40][44] * vector[40] +matrix[41][44] * vector[41] +matrix[42][44] * vector[42] +matrix[43][44] * vector[43] +matrix[44][44] * vector[44] +matrix[45][44] * vector[45] +matrix[46][44] * vector[46] +matrix[47][44] * vector[47] +matrix[48][44] * vector[48] +matrix[49][44] * vector[49] +matrix[50][44] * vector[50] +matrix[51][44] * vector[51] +matrix[52][44] * vector[52] +matrix[53][44] * vector[53] +matrix[54][44] * vector[54] +matrix[55][44] * vector[55] +matrix[56][44] * vector[56] +matrix[57][44] * vector[57] +matrix[58][44] * vector[58] +matrix[59][44] * vector[59] +matrix[60][44] * vector[60] +matrix[61][44] * vector[61] +matrix[62][44] * vector[62] +matrix[63][44] * vector[63] +matrix[64][44] * vector[64] +matrix[65][44] * vector[65] +matrix[66][44] * vector[66] +matrix[67][44] * vector[67] +matrix[68][44] * vector[68] +matrix[69][44] * vector[69] +matrix[70][44] * vector[70] +matrix[71][44] * vector[71] +matrix[72][44] * vector[72] +matrix[73][44] * vector[73] +matrix[74][44] * vector[74] +matrix[75][44] * vector[75] +matrix[76][44] * vector[76] +matrix[77][44] * vector[77] +matrix[78][44] * vector[78] +matrix[79][44] * vector[79] +matrix[80][44] * vector[80] +matrix[81][44] * vector[81] +matrix[82][44] * vector[82] +matrix[83][44] * vector[83] +matrix[84][44] * vector[84] +matrix[85][44] * vector[85] +matrix[86][44] * vector[86] +matrix[87][44] * vector[87] +matrix[88][44] * vector[88] +matrix[89][44] * vector[89] +matrix[90][44] * vector[90] +matrix[91][44] * vector[91] +matrix[92][44] * vector[92] +matrix[93][44] * vector[93] +matrix[94][44] * vector[94] +matrix[95][44] * vector[95] +matrix[96][44] * vector[96] +matrix[97][44] * vector[97] +matrix[98][44] * vector[98] +matrix[99][44] * vector[99] +b[44];
assign result[45] = matrix[0][45] * vector[0] +matrix[1][45] * vector[1] +matrix[2][45] * vector[2] +matrix[3][45] * vector[3] +matrix[4][45] * vector[4] +matrix[5][45] * vector[5] +matrix[6][45] * vector[6] +matrix[7][45] * vector[7] +matrix[8][45] * vector[8] +matrix[9][45] * vector[9] +matrix[10][45] * vector[10] +matrix[11][45] * vector[11] +matrix[12][45] * vector[12] +matrix[13][45] * vector[13] +matrix[14][45] * vector[14] +matrix[15][45] * vector[15] +matrix[16][45] * vector[16] +matrix[17][45] * vector[17] +matrix[18][45] * vector[18] +matrix[19][45] * vector[19] +matrix[20][45] * vector[20] +matrix[21][45] * vector[21] +matrix[22][45] * vector[22] +matrix[23][45] * vector[23] +matrix[24][45] * vector[24] +matrix[25][45] * vector[25] +matrix[26][45] * vector[26] +matrix[27][45] * vector[27] +matrix[28][45] * vector[28] +matrix[29][45] * vector[29] +matrix[30][45] * vector[30] +matrix[31][45] * vector[31] +matrix[32][45] * vector[32] +matrix[33][45] * vector[33] +matrix[34][45] * vector[34] +matrix[35][45] * vector[35] +matrix[36][45] * vector[36] +matrix[37][45] * vector[37] +matrix[38][45] * vector[38] +matrix[39][45] * vector[39] +matrix[40][45] * vector[40] +matrix[41][45] * vector[41] +matrix[42][45] * vector[42] +matrix[43][45] * vector[43] +matrix[44][45] * vector[44] +matrix[45][45] * vector[45] +matrix[46][45] * vector[46] +matrix[47][45] * vector[47] +matrix[48][45] * vector[48] +matrix[49][45] * vector[49] +matrix[50][45] * vector[50] +matrix[51][45] * vector[51] +matrix[52][45] * vector[52] +matrix[53][45] * vector[53] +matrix[54][45] * vector[54] +matrix[55][45] * vector[55] +matrix[56][45] * vector[56] +matrix[57][45] * vector[57] +matrix[58][45] * vector[58] +matrix[59][45] * vector[59] +matrix[60][45] * vector[60] +matrix[61][45] * vector[61] +matrix[62][45] * vector[62] +matrix[63][45] * vector[63] +matrix[64][45] * vector[64] +matrix[65][45] * vector[65] +matrix[66][45] * vector[66] +matrix[67][45] * vector[67] +matrix[68][45] * vector[68] +matrix[69][45] * vector[69] +matrix[70][45] * vector[70] +matrix[71][45] * vector[71] +matrix[72][45] * vector[72] +matrix[73][45] * vector[73] +matrix[74][45] * vector[74] +matrix[75][45] * vector[75] +matrix[76][45] * vector[76] +matrix[77][45] * vector[77] +matrix[78][45] * vector[78] +matrix[79][45] * vector[79] +matrix[80][45] * vector[80] +matrix[81][45] * vector[81] +matrix[82][45] * vector[82] +matrix[83][45] * vector[83] +matrix[84][45] * vector[84] +matrix[85][45] * vector[85] +matrix[86][45] * vector[86] +matrix[87][45] * vector[87] +matrix[88][45] * vector[88] +matrix[89][45] * vector[89] +matrix[90][45] * vector[90] +matrix[91][45] * vector[91] +matrix[92][45] * vector[92] +matrix[93][45] * vector[93] +matrix[94][45] * vector[94] +matrix[95][45] * vector[95] +matrix[96][45] * vector[96] +matrix[97][45] * vector[97] +matrix[98][45] * vector[98] +matrix[99][45] * vector[99] +b[45];
assign result[46] = matrix[0][46] * vector[0] +matrix[1][46] * vector[1] +matrix[2][46] * vector[2] +matrix[3][46] * vector[3] +matrix[4][46] * vector[4] +matrix[5][46] * vector[5] +matrix[6][46] * vector[6] +matrix[7][46] * vector[7] +matrix[8][46] * vector[8] +matrix[9][46] * vector[9] +matrix[10][46] * vector[10] +matrix[11][46] * vector[11] +matrix[12][46] * vector[12] +matrix[13][46] * vector[13] +matrix[14][46] * vector[14] +matrix[15][46] * vector[15] +matrix[16][46] * vector[16] +matrix[17][46] * vector[17] +matrix[18][46] * vector[18] +matrix[19][46] * vector[19] +matrix[20][46] * vector[20] +matrix[21][46] * vector[21] +matrix[22][46] * vector[22] +matrix[23][46] * vector[23] +matrix[24][46] * vector[24] +matrix[25][46] * vector[25] +matrix[26][46] * vector[26] +matrix[27][46] * vector[27] +matrix[28][46] * vector[28] +matrix[29][46] * vector[29] +matrix[30][46] * vector[30] +matrix[31][46] * vector[31] +matrix[32][46] * vector[32] +matrix[33][46] * vector[33] +matrix[34][46] * vector[34] +matrix[35][46] * vector[35] +matrix[36][46] * vector[36] +matrix[37][46] * vector[37] +matrix[38][46] * vector[38] +matrix[39][46] * vector[39] +matrix[40][46] * vector[40] +matrix[41][46] * vector[41] +matrix[42][46] * vector[42] +matrix[43][46] * vector[43] +matrix[44][46] * vector[44] +matrix[45][46] * vector[45] +matrix[46][46] * vector[46] +matrix[47][46] * vector[47] +matrix[48][46] * vector[48] +matrix[49][46] * vector[49] +matrix[50][46] * vector[50] +matrix[51][46] * vector[51] +matrix[52][46] * vector[52] +matrix[53][46] * vector[53] +matrix[54][46] * vector[54] +matrix[55][46] * vector[55] +matrix[56][46] * vector[56] +matrix[57][46] * vector[57] +matrix[58][46] * vector[58] +matrix[59][46] * vector[59] +matrix[60][46] * vector[60] +matrix[61][46] * vector[61] +matrix[62][46] * vector[62] +matrix[63][46] * vector[63] +matrix[64][46] * vector[64] +matrix[65][46] * vector[65] +matrix[66][46] * vector[66] +matrix[67][46] * vector[67] +matrix[68][46] * vector[68] +matrix[69][46] * vector[69] +matrix[70][46] * vector[70] +matrix[71][46] * vector[71] +matrix[72][46] * vector[72] +matrix[73][46] * vector[73] +matrix[74][46] * vector[74] +matrix[75][46] * vector[75] +matrix[76][46] * vector[76] +matrix[77][46] * vector[77] +matrix[78][46] * vector[78] +matrix[79][46] * vector[79] +matrix[80][46] * vector[80] +matrix[81][46] * vector[81] +matrix[82][46] * vector[82] +matrix[83][46] * vector[83] +matrix[84][46] * vector[84] +matrix[85][46] * vector[85] +matrix[86][46] * vector[86] +matrix[87][46] * vector[87] +matrix[88][46] * vector[88] +matrix[89][46] * vector[89] +matrix[90][46] * vector[90] +matrix[91][46] * vector[91] +matrix[92][46] * vector[92] +matrix[93][46] * vector[93] +matrix[94][46] * vector[94] +matrix[95][46] * vector[95] +matrix[96][46] * vector[96] +matrix[97][46] * vector[97] +matrix[98][46] * vector[98] +matrix[99][46] * vector[99] +b[46];
assign result[47] = matrix[0][47] * vector[0] +matrix[1][47] * vector[1] +matrix[2][47] * vector[2] +matrix[3][47] * vector[3] +matrix[4][47] * vector[4] +matrix[5][47] * vector[5] +matrix[6][47] * vector[6] +matrix[7][47] * vector[7] +matrix[8][47] * vector[8] +matrix[9][47] * vector[9] +matrix[10][47] * vector[10] +matrix[11][47] * vector[11] +matrix[12][47] * vector[12] +matrix[13][47] * vector[13] +matrix[14][47] * vector[14] +matrix[15][47] * vector[15] +matrix[16][47] * vector[16] +matrix[17][47] * vector[17] +matrix[18][47] * vector[18] +matrix[19][47] * vector[19] +matrix[20][47] * vector[20] +matrix[21][47] * vector[21] +matrix[22][47] * vector[22] +matrix[23][47] * vector[23] +matrix[24][47] * vector[24] +matrix[25][47] * vector[25] +matrix[26][47] * vector[26] +matrix[27][47] * vector[27] +matrix[28][47] * vector[28] +matrix[29][47] * vector[29] +matrix[30][47] * vector[30] +matrix[31][47] * vector[31] +matrix[32][47] * vector[32] +matrix[33][47] * vector[33] +matrix[34][47] * vector[34] +matrix[35][47] * vector[35] +matrix[36][47] * vector[36] +matrix[37][47] * vector[37] +matrix[38][47] * vector[38] +matrix[39][47] * vector[39] +matrix[40][47] * vector[40] +matrix[41][47] * vector[41] +matrix[42][47] * vector[42] +matrix[43][47] * vector[43] +matrix[44][47] * vector[44] +matrix[45][47] * vector[45] +matrix[46][47] * vector[46] +matrix[47][47] * vector[47] +matrix[48][47] * vector[48] +matrix[49][47] * vector[49] +matrix[50][47] * vector[50] +matrix[51][47] * vector[51] +matrix[52][47] * vector[52] +matrix[53][47] * vector[53] +matrix[54][47] * vector[54] +matrix[55][47] * vector[55] +matrix[56][47] * vector[56] +matrix[57][47] * vector[57] +matrix[58][47] * vector[58] +matrix[59][47] * vector[59] +matrix[60][47] * vector[60] +matrix[61][47] * vector[61] +matrix[62][47] * vector[62] +matrix[63][47] * vector[63] +matrix[64][47] * vector[64] +matrix[65][47] * vector[65] +matrix[66][47] * vector[66] +matrix[67][47] * vector[67] +matrix[68][47] * vector[68] +matrix[69][47] * vector[69] +matrix[70][47] * vector[70] +matrix[71][47] * vector[71] +matrix[72][47] * vector[72] +matrix[73][47] * vector[73] +matrix[74][47] * vector[74] +matrix[75][47] * vector[75] +matrix[76][47] * vector[76] +matrix[77][47] * vector[77] +matrix[78][47] * vector[78] +matrix[79][47] * vector[79] +matrix[80][47] * vector[80] +matrix[81][47] * vector[81] +matrix[82][47] * vector[82] +matrix[83][47] * vector[83] +matrix[84][47] * vector[84] +matrix[85][47] * vector[85] +matrix[86][47] * vector[86] +matrix[87][47] * vector[87] +matrix[88][47] * vector[88] +matrix[89][47] * vector[89] +matrix[90][47] * vector[90] +matrix[91][47] * vector[91] +matrix[92][47] * vector[92] +matrix[93][47] * vector[93] +matrix[94][47] * vector[94] +matrix[95][47] * vector[95] +matrix[96][47] * vector[96] +matrix[97][47] * vector[97] +matrix[98][47] * vector[98] +matrix[99][47] * vector[99] +b[47];
assign result[48] = matrix[0][48] * vector[0] +matrix[1][48] * vector[1] +matrix[2][48] * vector[2] +matrix[3][48] * vector[3] +matrix[4][48] * vector[4] +matrix[5][48] * vector[5] +matrix[6][48] * vector[6] +matrix[7][48] * vector[7] +matrix[8][48] * vector[8] +matrix[9][48] * vector[9] +matrix[10][48] * vector[10] +matrix[11][48] * vector[11] +matrix[12][48] * vector[12] +matrix[13][48] * vector[13] +matrix[14][48] * vector[14] +matrix[15][48] * vector[15] +matrix[16][48] * vector[16] +matrix[17][48] * vector[17] +matrix[18][48] * vector[18] +matrix[19][48] * vector[19] +matrix[20][48] * vector[20] +matrix[21][48] * vector[21] +matrix[22][48] * vector[22] +matrix[23][48] * vector[23] +matrix[24][48] * vector[24] +matrix[25][48] * vector[25] +matrix[26][48] * vector[26] +matrix[27][48] * vector[27] +matrix[28][48] * vector[28] +matrix[29][48] * vector[29] +matrix[30][48] * vector[30] +matrix[31][48] * vector[31] +matrix[32][48] * vector[32] +matrix[33][48] * vector[33] +matrix[34][48] * vector[34] +matrix[35][48] * vector[35] +matrix[36][48] * vector[36] +matrix[37][48] * vector[37] +matrix[38][48] * vector[38] +matrix[39][48] * vector[39] +matrix[40][48] * vector[40] +matrix[41][48] * vector[41] +matrix[42][48] * vector[42] +matrix[43][48] * vector[43] +matrix[44][48] * vector[44] +matrix[45][48] * vector[45] +matrix[46][48] * vector[46] +matrix[47][48] * vector[47] +matrix[48][48] * vector[48] +matrix[49][48] * vector[49] +matrix[50][48] * vector[50] +matrix[51][48] * vector[51] +matrix[52][48] * vector[52] +matrix[53][48] * vector[53] +matrix[54][48] * vector[54] +matrix[55][48] * vector[55] +matrix[56][48] * vector[56] +matrix[57][48] * vector[57] +matrix[58][48] * vector[58] +matrix[59][48] * vector[59] +matrix[60][48] * vector[60] +matrix[61][48] * vector[61] +matrix[62][48] * vector[62] +matrix[63][48] * vector[63] +matrix[64][48] * vector[64] +matrix[65][48] * vector[65] +matrix[66][48] * vector[66] +matrix[67][48] * vector[67] +matrix[68][48] * vector[68] +matrix[69][48] * vector[69] +matrix[70][48] * vector[70] +matrix[71][48] * vector[71] +matrix[72][48] * vector[72] +matrix[73][48] * vector[73] +matrix[74][48] * vector[74] +matrix[75][48] * vector[75] +matrix[76][48] * vector[76] +matrix[77][48] * vector[77] +matrix[78][48] * vector[78] +matrix[79][48] * vector[79] +matrix[80][48] * vector[80] +matrix[81][48] * vector[81] +matrix[82][48] * vector[82] +matrix[83][48] * vector[83] +matrix[84][48] * vector[84] +matrix[85][48] * vector[85] +matrix[86][48] * vector[86] +matrix[87][48] * vector[87] +matrix[88][48] * vector[88] +matrix[89][48] * vector[89] +matrix[90][48] * vector[90] +matrix[91][48] * vector[91] +matrix[92][48] * vector[92] +matrix[93][48] * vector[93] +matrix[94][48] * vector[94] +matrix[95][48] * vector[95] +matrix[96][48] * vector[96] +matrix[97][48] * vector[97] +matrix[98][48] * vector[98] +matrix[99][48] * vector[99] +b[48];
assign result[49] = matrix[0][49] * vector[0] +matrix[1][49] * vector[1] +matrix[2][49] * vector[2] +matrix[3][49] * vector[3] +matrix[4][49] * vector[4] +matrix[5][49] * vector[5] +matrix[6][49] * vector[6] +matrix[7][49] * vector[7] +matrix[8][49] * vector[8] +matrix[9][49] * vector[9] +matrix[10][49] * vector[10] +matrix[11][49] * vector[11] +matrix[12][49] * vector[12] +matrix[13][49] * vector[13] +matrix[14][49] * vector[14] +matrix[15][49] * vector[15] +matrix[16][49] * vector[16] +matrix[17][49] * vector[17] +matrix[18][49] * vector[18] +matrix[19][49] * vector[19] +matrix[20][49] * vector[20] +matrix[21][49] * vector[21] +matrix[22][49] * vector[22] +matrix[23][49] * vector[23] +matrix[24][49] * vector[24] +matrix[25][49] * vector[25] +matrix[26][49] * vector[26] +matrix[27][49] * vector[27] +matrix[28][49] * vector[28] +matrix[29][49] * vector[29] +matrix[30][49] * vector[30] +matrix[31][49] * vector[31] +matrix[32][49] * vector[32] +matrix[33][49] * vector[33] +matrix[34][49] * vector[34] +matrix[35][49] * vector[35] +matrix[36][49] * vector[36] +matrix[37][49] * vector[37] +matrix[38][49] * vector[38] +matrix[39][49] * vector[39] +matrix[40][49] * vector[40] +matrix[41][49] * vector[41] +matrix[42][49] * vector[42] +matrix[43][49] * vector[43] +matrix[44][49] * vector[44] +matrix[45][49] * vector[45] +matrix[46][49] * vector[46] +matrix[47][49] * vector[47] +matrix[48][49] * vector[48] +matrix[49][49] * vector[49] +matrix[50][49] * vector[50] +matrix[51][49] * vector[51] +matrix[52][49] * vector[52] +matrix[53][49] * vector[53] +matrix[54][49] * vector[54] +matrix[55][49] * vector[55] +matrix[56][49] * vector[56] +matrix[57][49] * vector[57] +matrix[58][49] * vector[58] +matrix[59][49] * vector[59] +matrix[60][49] * vector[60] +matrix[61][49] * vector[61] +matrix[62][49] * vector[62] +matrix[63][49] * vector[63] +matrix[64][49] * vector[64] +matrix[65][49] * vector[65] +matrix[66][49] * vector[66] +matrix[67][49] * vector[67] +matrix[68][49] * vector[68] +matrix[69][49] * vector[69] +matrix[70][49] * vector[70] +matrix[71][49] * vector[71] +matrix[72][49] * vector[72] +matrix[73][49] * vector[73] +matrix[74][49] * vector[74] +matrix[75][49] * vector[75] +matrix[76][49] * vector[76] +matrix[77][49] * vector[77] +matrix[78][49] * vector[78] +matrix[79][49] * vector[79] +matrix[80][49] * vector[80] +matrix[81][49] * vector[81] +matrix[82][49] * vector[82] +matrix[83][49] * vector[83] +matrix[84][49] * vector[84] +matrix[85][49] * vector[85] +matrix[86][49] * vector[86] +matrix[87][49] * vector[87] +matrix[88][49] * vector[88] +matrix[89][49] * vector[89] +matrix[90][49] * vector[90] +matrix[91][49] * vector[91] +matrix[92][49] * vector[92] +matrix[93][49] * vector[93] +matrix[94][49] * vector[94] +matrix[95][49] * vector[95] +matrix[96][49] * vector[96] +matrix[97][49] * vector[97] +matrix[98][49] * vector[98] +matrix[99][49] * vector[99] +b[49];
assign result[50] = matrix[0][50] * vector[0] +matrix[1][50] * vector[1] +matrix[2][50] * vector[2] +matrix[3][50] * vector[3] +matrix[4][50] * vector[4] +matrix[5][50] * vector[5] +matrix[6][50] * vector[6] +matrix[7][50] * vector[7] +matrix[8][50] * vector[8] +matrix[9][50] * vector[9] +matrix[10][50] * vector[10] +matrix[11][50] * vector[11] +matrix[12][50] * vector[12] +matrix[13][50] * vector[13] +matrix[14][50] * vector[14] +matrix[15][50] * vector[15] +matrix[16][50] * vector[16] +matrix[17][50] * vector[17] +matrix[18][50] * vector[18] +matrix[19][50] * vector[19] +matrix[20][50] * vector[20] +matrix[21][50] * vector[21] +matrix[22][50] * vector[22] +matrix[23][50] * vector[23] +matrix[24][50] * vector[24] +matrix[25][50] * vector[25] +matrix[26][50] * vector[26] +matrix[27][50] * vector[27] +matrix[28][50] * vector[28] +matrix[29][50] * vector[29] +matrix[30][50] * vector[30] +matrix[31][50] * vector[31] +matrix[32][50] * vector[32] +matrix[33][50] * vector[33] +matrix[34][50] * vector[34] +matrix[35][50] * vector[35] +matrix[36][50] * vector[36] +matrix[37][50] * vector[37] +matrix[38][50] * vector[38] +matrix[39][50] * vector[39] +matrix[40][50] * vector[40] +matrix[41][50] * vector[41] +matrix[42][50] * vector[42] +matrix[43][50] * vector[43] +matrix[44][50] * vector[44] +matrix[45][50] * vector[45] +matrix[46][50] * vector[46] +matrix[47][50] * vector[47] +matrix[48][50] * vector[48] +matrix[49][50] * vector[49] +matrix[50][50] * vector[50] +matrix[51][50] * vector[51] +matrix[52][50] * vector[52] +matrix[53][50] * vector[53] +matrix[54][50] * vector[54] +matrix[55][50] * vector[55] +matrix[56][50] * vector[56] +matrix[57][50] * vector[57] +matrix[58][50] * vector[58] +matrix[59][50] * vector[59] +matrix[60][50] * vector[60] +matrix[61][50] * vector[61] +matrix[62][50] * vector[62] +matrix[63][50] * vector[63] +matrix[64][50] * vector[64] +matrix[65][50] * vector[65] +matrix[66][50] * vector[66] +matrix[67][50] * vector[67] +matrix[68][50] * vector[68] +matrix[69][50] * vector[69] +matrix[70][50] * vector[70] +matrix[71][50] * vector[71] +matrix[72][50] * vector[72] +matrix[73][50] * vector[73] +matrix[74][50] * vector[74] +matrix[75][50] * vector[75] +matrix[76][50] * vector[76] +matrix[77][50] * vector[77] +matrix[78][50] * vector[78] +matrix[79][50] * vector[79] +matrix[80][50] * vector[80] +matrix[81][50] * vector[81] +matrix[82][50] * vector[82] +matrix[83][50] * vector[83] +matrix[84][50] * vector[84] +matrix[85][50] * vector[85] +matrix[86][50] * vector[86] +matrix[87][50] * vector[87] +matrix[88][50] * vector[88] +matrix[89][50] * vector[89] +matrix[90][50] * vector[90] +matrix[91][50] * vector[91] +matrix[92][50] * vector[92] +matrix[93][50] * vector[93] +matrix[94][50] * vector[94] +matrix[95][50] * vector[95] +matrix[96][50] * vector[96] +matrix[97][50] * vector[97] +matrix[98][50] * vector[98] +matrix[99][50] * vector[99] +b[50];
assign result[51] = matrix[0][51] * vector[0] +matrix[1][51] * vector[1] +matrix[2][51] * vector[2] +matrix[3][51] * vector[3] +matrix[4][51] * vector[4] +matrix[5][51] * vector[5] +matrix[6][51] * vector[6] +matrix[7][51] * vector[7] +matrix[8][51] * vector[8] +matrix[9][51] * vector[9] +matrix[10][51] * vector[10] +matrix[11][51] * vector[11] +matrix[12][51] * vector[12] +matrix[13][51] * vector[13] +matrix[14][51] * vector[14] +matrix[15][51] * vector[15] +matrix[16][51] * vector[16] +matrix[17][51] * vector[17] +matrix[18][51] * vector[18] +matrix[19][51] * vector[19] +matrix[20][51] * vector[20] +matrix[21][51] * vector[21] +matrix[22][51] * vector[22] +matrix[23][51] * vector[23] +matrix[24][51] * vector[24] +matrix[25][51] * vector[25] +matrix[26][51] * vector[26] +matrix[27][51] * vector[27] +matrix[28][51] * vector[28] +matrix[29][51] * vector[29] +matrix[30][51] * vector[30] +matrix[31][51] * vector[31] +matrix[32][51] * vector[32] +matrix[33][51] * vector[33] +matrix[34][51] * vector[34] +matrix[35][51] * vector[35] +matrix[36][51] * vector[36] +matrix[37][51] * vector[37] +matrix[38][51] * vector[38] +matrix[39][51] * vector[39] +matrix[40][51] * vector[40] +matrix[41][51] * vector[41] +matrix[42][51] * vector[42] +matrix[43][51] * vector[43] +matrix[44][51] * vector[44] +matrix[45][51] * vector[45] +matrix[46][51] * vector[46] +matrix[47][51] * vector[47] +matrix[48][51] * vector[48] +matrix[49][51] * vector[49] +matrix[50][51] * vector[50] +matrix[51][51] * vector[51] +matrix[52][51] * vector[52] +matrix[53][51] * vector[53] +matrix[54][51] * vector[54] +matrix[55][51] * vector[55] +matrix[56][51] * vector[56] +matrix[57][51] * vector[57] +matrix[58][51] * vector[58] +matrix[59][51] * vector[59] +matrix[60][51] * vector[60] +matrix[61][51] * vector[61] +matrix[62][51] * vector[62] +matrix[63][51] * vector[63] +matrix[64][51] * vector[64] +matrix[65][51] * vector[65] +matrix[66][51] * vector[66] +matrix[67][51] * vector[67] +matrix[68][51] * vector[68] +matrix[69][51] * vector[69] +matrix[70][51] * vector[70] +matrix[71][51] * vector[71] +matrix[72][51] * vector[72] +matrix[73][51] * vector[73] +matrix[74][51] * vector[74] +matrix[75][51] * vector[75] +matrix[76][51] * vector[76] +matrix[77][51] * vector[77] +matrix[78][51] * vector[78] +matrix[79][51] * vector[79] +matrix[80][51] * vector[80] +matrix[81][51] * vector[81] +matrix[82][51] * vector[82] +matrix[83][51] * vector[83] +matrix[84][51] * vector[84] +matrix[85][51] * vector[85] +matrix[86][51] * vector[86] +matrix[87][51] * vector[87] +matrix[88][51] * vector[88] +matrix[89][51] * vector[89] +matrix[90][51] * vector[90] +matrix[91][51] * vector[91] +matrix[92][51] * vector[92] +matrix[93][51] * vector[93] +matrix[94][51] * vector[94] +matrix[95][51] * vector[95] +matrix[96][51] * vector[96] +matrix[97][51] * vector[97] +matrix[98][51] * vector[98] +matrix[99][51] * vector[99] +b[51];
assign result[52] = matrix[0][52] * vector[0] +matrix[1][52] * vector[1] +matrix[2][52] * vector[2] +matrix[3][52] * vector[3] +matrix[4][52] * vector[4] +matrix[5][52] * vector[5] +matrix[6][52] * vector[6] +matrix[7][52] * vector[7] +matrix[8][52] * vector[8] +matrix[9][52] * vector[9] +matrix[10][52] * vector[10] +matrix[11][52] * vector[11] +matrix[12][52] * vector[12] +matrix[13][52] * vector[13] +matrix[14][52] * vector[14] +matrix[15][52] * vector[15] +matrix[16][52] * vector[16] +matrix[17][52] * vector[17] +matrix[18][52] * vector[18] +matrix[19][52] * vector[19] +matrix[20][52] * vector[20] +matrix[21][52] * vector[21] +matrix[22][52] * vector[22] +matrix[23][52] * vector[23] +matrix[24][52] * vector[24] +matrix[25][52] * vector[25] +matrix[26][52] * vector[26] +matrix[27][52] * vector[27] +matrix[28][52] * vector[28] +matrix[29][52] * vector[29] +matrix[30][52] * vector[30] +matrix[31][52] * vector[31] +matrix[32][52] * vector[32] +matrix[33][52] * vector[33] +matrix[34][52] * vector[34] +matrix[35][52] * vector[35] +matrix[36][52] * vector[36] +matrix[37][52] * vector[37] +matrix[38][52] * vector[38] +matrix[39][52] * vector[39] +matrix[40][52] * vector[40] +matrix[41][52] * vector[41] +matrix[42][52] * vector[42] +matrix[43][52] * vector[43] +matrix[44][52] * vector[44] +matrix[45][52] * vector[45] +matrix[46][52] * vector[46] +matrix[47][52] * vector[47] +matrix[48][52] * vector[48] +matrix[49][52] * vector[49] +matrix[50][52] * vector[50] +matrix[51][52] * vector[51] +matrix[52][52] * vector[52] +matrix[53][52] * vector[53] +matrix[54][52] * vector[54] +matrix[55][52] * vector[55] +matrix[56][52] * vector[56] +matrix[57][52] * vector[57] +matrix[58][52] * vector[58] +matrix[59][52] * vector[59] +matrix[60][52] * vector[60] +matrix[61][52] * vector[61] +matrix[62][52] * vector[62] +matrix[63][52] * vector[63] +matrix[64][52] * vector[64] +matrix[65][52] * vector[65] +matrix[66][52] * vector[66] +matrix[67][52] * vector[67] +matrix[68][52] * vector[68] +matrix[69][52] * vector[69] +matrix[70][52] * vector[70] +matrix[71][52] * vector[71] +matrix[72][52] * vector[72] +matrix[73][52] * vector[73] +matrix[74][52] * vector[74] +matrix[75][52] * vector[75] +matrix[76][52] * vector[76] +matrix[77][52] * vector[77] +matrix[78][52] * vector[78] +matrix[79][52] * vector[79] +matrix[80][52] * vector[80] +matrix[81][52] * vector[81] +matrix[82][52] * vector[82] +matrix[83][52] * vector[83] +matrix[84][52] * vector[84] +matrix[85][52] * vector[85] +matrix[86][52] * vector[86] +matrix[87][52] * vector[87] +matrix[88][52] * vector[88] +matrix[89][52] * vector[89] +matrix[90][52] * vector[90] +matrix[91][52] * vector[91] +matrix[92][52] * vector[92] +matrix[93][52] * vector[93] +matrix[94][52] * vector[94] +matrix[95][52] * vector[95] +matrix[96][52] * vector[96] +matrix[97][52] * vector[97] +matrix[98][52] * vector[98] +matrix[99][52] * vector[99] +b[52];
assign result[53] = matrix[0][53] * vector[0] +matrix[1][53] * vector[1] +matrix[2][53] * vector[2] +matrix[3][53] * vector[3] +matrix[4][53] * vector[4] +matrix[5][53] * vector[5] +matrix[6][53] * vector[6] +matrix[7][53] * vector[7] +matrix[8][53] * vector[8] +matrix[9][53] * vector[9] +matrix[10][53] * vector[10] +matrix[11][53] * vector[11] +matrix[12][53] * vector[12] +matrix[13][53] * vector[13] +matrix[14][53] * vector[14] +matrix[15][53] * vector[15] +matrix[16][53] * vector[16] +matrix[17][53] * vector[17] +matrix[18][53] * vector[18] +matrix[19][53] * vector[19] +matrix[20][53] * vector[20] +matrix[21][53] * vector[21] +matrix[22][53] * vector[22] +matrix[23][53] * vector[23] +matrix[24][53] * vector[24] +matrix[25][53] * vector[25] +matrix[26][53] * vector[26] +matrix[27][53] * vector[27] +matrix[28][53] * vector[28] +matrix[29][53] * vector[29] +matrix[30][53] * vector[30] +matrix[31][53] * vector[31] +matrix[32][53] * vector[32] +matrix[33][53] * vector[33] +matrix[34][53] * vector[34] +matrix[35][53] * vector[35] +matrix[36][53] * vector[36] +matrix[37][53] * vector[37] +matrix[38][53] * vector[38] +matrix[39][53] * vector[39] +matrix[40][53] * vector[40] +matrix[41][53] * vector[41] +matrix[42][53] * vector[42] +matrix[43][53] * vector[43] +matrix[44][53] * vector[44] +matrix[45][53] * vector[45] +matrix[46][53] * vector[46] +matrix[47][53] * vector[47] +matrix[48][53] * vector[48] +matrix[49][53] * vector[49] +matrix[50][53] * vector[50] +matrix[51][53] * vector[51] +matrix[52][53] * vector[52] +matrix[53][53] * vector[53] +matrix[54][53] * vector[54] +matrix[55][53] * vector[55] +matrix[56][53] * vector[56] +matrix[57][53] * vector[57] +matrix[58][53] * vector[58] +matrix[59][53] * vector[59] +matrix[60][53] * vector[60] +matrix[61][53] * vector[61] +matrix[62][53] * vector[62] +matrix[63][53] * vector[63] +matrix[64][53] * vector[64] +matrix[65][53] * vector[65] +matrix[66][53] * vector[66] +matrix[67][53] * vector[67] +matrix[68][53] * vector[68] +matrix[69][53] * vector[69] +matrix[70][53] * vector[70] +matrix[71][53] * vector[71] +matrix[72][53] * vector[72] +matrix[73][53] * vector[73] +matrix[74][53] * vector[74] +matrix[75][53] * vector[75] +matrix[76][53] * vector[76] +matrix[77][53] * vector[77] +matrix[78][53] * vector[78] +matrix[79][53] * vector[79] +matrix[80][53] * vector[80] +matrix[81][53] * vector[81] +matrix[82][53] * vector[82] +matrix[83][53] * vector[83] +matrix[84][53] * vector[84] +matrix[85][53] * vector[85] +matrix[86][53] * vector[86] +matrix[87][53] * vector[87] +matrix[88][53] * vector[88] +matrix[89][53] * vector[89] +matrix[90][53] * vector[90] +matrix[91][53] * vector[91] +matrix[92][53] * vector[92] +matrix[93][53] * vector[93] +matrix[94][53] * vector[94] +matrix[95][53] * vector[95] +matrix[96][53] * vector[96] +matrix[97][53] * vector[97] +matrix[98][53] * vector[98] +matrix[99][53] * vector[99] +b[53];
assign result[54] = matrix[0][54] * vector[0] +matrix[1][54] * vector[1] +matrix[2][54] * vector[2] +matrix[3][54] * vector[3] +matrix[4][54] * vector[4] +matrix[5][54] * vector[5] +matrix[6][54] * vector[6] +matrix[7][54] * vector[7] +matrix[8][54] * vector[8] +matrix[9][54] * vector[9] +matrix[10][54] * vector[10] +matrix[11][54] * vector[11] +matrix[12][54] * vector[12] +matrix[13][54] * vector[13] +matrix[14][54] * vector[14] +matrix[15][54] * vector[15] +matrix[16][54] * vector[16] +matrix[17][54] * vector[17] +matrix[18][54] * vector[18] +matrix[19][54] * vector[19] +matrix[20][54] * vector[20] +matrix[21][54] * vector[21] +matrix[22][54] * vector[22] +matrix[23][54] * vector[23] +matrix[24][54] * vector[24] +matrix[25][54] * vector[25] +matrix[26][54] * vector[26] +matrix[27][54] * vector[27] +matrix[28][54] * vector[28] +matrix[29][54] * vector[29] +matrix[30][54] * vector[30] +matrix[31][54] * vector[31] +matrix[32][54] * vector[32] +matrix[33][54] * vector[33] +matrix[34][54] * vector[34] +matrix[35][54] * vector[35] +matrix[36][54] * vector[36] +matrix[37][54] * vector[37] +matrix[38][54] * vector[38] +matrix[39][54] * vector[39] +matrix[40][54] * vector[40] +matrix[41][54] * vector[41] +matrix[42][54] * vector[42] +matrix[43][54] * vector[43] +matrix[44][54] * vector[44] +matrix[45][54] * vector[45] +matrix[46][54] * vector[46] +matrix[47][54] * vector[47] +matrix[48][54] * vector[48] +matrix[49][54] * vector[49] +matrix[50][54] * vector[50] +matrix[51][54] * vector[51] +matrix[52][54] * vector[52] +matrix[53][54] * vector[53] +matrix[54][54] * vector[54] +matrix[55][54] * vector[55] +matrix[56][54] * vector[56] +matrix[57][54] * vector[57] +matrix[58][54] * vector[58] +matrix[59][54] * vector[59] +matrix[60][54] * vector[60] +matrix[61][54] * vector[61] +matrix[62][54] * vector[62] +matrix[63][54] * vector[63] +matrix[64][54] * vector[64] +matrix[65][54] * vector[65] +matrix[66][54] * vector[66] +matrix[67][54] * vector[67] +matrix[68][54] * vector[68] +matrix[69][54] * vector[69] +matrix[70][54] * vector[70] +matrix[71][54] * vector[71] +matrix[72][54] * vector[72] +matrix[73][54] * vector[73] +matrix[74][54] * vector[74] +matrix[75][54] * vector[75] +matrix[76][54] * vector[76] +matrix[77][54] * vector[77] +matrix[78][54] * vector[78] +matrix[79][54] * vector[79] +matrix[80][54] * vector[80] +matrix[81][54] * vector[81] +matrix[82][54] * vector[82] +matrix[83][54] * vector[83] +matrix[84][54] * vector[84] +matrix[85][54] * vector[85] +matrix[86][54] * vector[86] +matrix[87][54] * vector[87] +matrix[88][54] * vector[88] +matrix[89][54] * vector[89] +matrix[90][54] * vector[90] +matrix[91][54] * vector[91] +matrix[92][54] * vector[92] +matrix[93][54] * vector[93] +matrix[94][54] * vector[94] +matrix[95][54] * vector[95] +matrix[96][54] * vector[96] +matrix[97][54] * vector[97] +matrix[98][54] * vector[98] +matrix[99][54] * vector[99] +b[54];
assign result[55] = matrix[0][55] * vector[0] +matrix[1][55] * vector[1] +matrix[2][55] * vector[2] +matrix[3][55] * vector[3] +matrix[4][55] * vector[4] +matrix[5][55] * vector[5] +matrix[6][55] * vector[6] +matrix[7][55] * vector[7] +matrix[8][55] * vector[8] +matrix[9][55] * vector[9] +matrix[10][55] * vector[10] +matrix[11][55] * vector[11] +matrix[12][55] * vector[12] +matrix[13][55] * vector[13] +matrix[14][55] * vector[14] +matrix[15][55] * vector[15] +matrix[16][55] * vector[16] +matrix[17][55] * vector[17] +matrix[18][55] * vector[18] +matrix[19][55] * vector[19] +matrix[20][55] * vector[20] +matrix[21][55] * vector[21] +matrix[22][55] * vector[22] +matrix[23][55] * vector[23] +matrix[24][55] * vector[24] +matrix[25][55] * vector[25] +matrix[26][55] * vector[26] +matrix[27][55] * vector[27] +matrix[28][55] * vector[28] +matrix[29][55] * vector[29] +matrix[30][55] * vector[30] +matrix[31][55] * vector[31] +matrix[32][55] * vector[32] +matrix[33][55] * vector[33] +matrix[34][55] * vector[34] +matrix[35][55] * vector[35] +matrix[36][55] * vector[36] +matrix[37][55] * vector[37] +matrix[38][55] * vector[38] +matrix[39][55] * vector[39] +matrix[40][55] * vector[40] +matrix[41][55] * vector[41] +matrix[42][55] * vector[42] +matrix[43][55] * vector[43] +matrix[44][55] * vector[44] +matrix[45][55] * vector[45] +matrix[46][55] * vector[46] +matrix[47][55] * vector[47] +matrix[48][55] * vector[48] +matrix[49][55] * vector[49] +matrix[50][55] * vector[50] +matrix[51][55] * vector[51] +matrix[52][55] * vector[52] +matrix[53][55] * vector[53] +matrix[54][55] * vector[54] +matrix[55][55] * vector[55] +matrix[56][55] * vector[56] +matrix[57][55] * vector[57] +matrix[58][55] * vector[58] +matrix[59][55] * vector[59] +matrix[60][55] * vector[60] +matrix[61][55] * vector[61] +matrix[62][55] * vector[62] +matrix[63][55] * vector[63] +matrix[64][55] * vector[64] +matrix[65][55] * vector[65] +matrix[66][55] * vector[66] +matrix[67][55] * vector[67] +matrix[68][55] * vector[68] +matrix[69][55] * vector[69] +matrix[70][55] * vector[70] +matrix[71][55] * vector[71] +matrix[72][55] * vector[72] +matrix[73][55] * vector[73] +matrix[74][55] * vector[74] +matrix[75][55] * vector[75] +matrix[76][55] * vector[76] +matrix[77][55] * vector[77] +matrix[78][55] * vector[78] +matrix[79][55] * vector[79] +matrix[80][55] * vector[80] +matrix[81][55] * vector[81] +matrix[82][55] * vector[82] +matrix[83][55] * vector[83] +matrix[84][55] * vector[84] +matrix[85][55] * vector[85] +matrix[86][55] * vector[86] +matrix[87][55] * vector[87] +matrix[88][55] * vector[88] +matrix[89][55] * vector[89] +matrix[90][55] * vector[90] +matrix[91][55] * vector[91] +matrix[92][55] * vector[92] +matrix[93][55] * vector[93] +matrix[94][55] * vector[94] +matrix[95][55] * vector[95] +matrix[96][55] * vector[96] +matrix[97][55] * vector[97] +matrix[98][55] * vector[98] +matrix[99][55] * vector[99] +b[55];
assign result[56] = matrix[0][56] * vector[0] +matrix[1][56] * vector[1] +matrix[2][56] * vector[2] +matrix[3][56] * vector[3] +matrix[4][56] * vector[4] +matrix[5][56] * vector[5] +matrix[6][56] * vector[6] +matrix[7][56] * vector[7] +matrix[8][56] * vector[8] +matrix[9][56] * vector[9] +matrix[10][56] * vector[10] +matrix[11][56] * vector[11] +matrix[12][56] * vector[12] +matrix[13][56] * vector[13] +matrix[14][56] * vector[14] +matrix[15][56] * vector[15] +matrix[16][56] * vector[16] +matrix[17][56] * vector[17] +matrix[18][56] * vector[18] +matrix[19][56] * vector[19] +matrix[20][56] * vector[20] +matrix[21][56] * vector[21] +matrix[22][56] * vector[22] +matrix[23][56] * vector[23] +matrix[24][56] * vector[24] +matrix[25][56] * vector[25] +matrix[26][56] * vector[26] +matrix[27][56] * vector[27] +matrix[28][56] * vector[28] +matrix[29][56] * vector[29] +matrix[30][56] * vector[30] +matrix[31][56] * vector[31] +matrix[32][56] * vector[32] +matrix[33][56] * vector[33] +matrix[34][56] * vector[34] +matrix[35][56] * vector[35] +matrix[36][56] * vector[36] +matrix[37][56] * vector[37] +matrix[38][56] * vector[38] +matrix[39][56] * vector[39] +matrix[40][56] * vector[40] +matrix[41][56] * vector[41] +matrix[42][56] * vector[42] +matrix[43][56] * vector[43] +matrix[44][56] * vector[44] +matrix[45][56] * vector[45] +matrix[46][56] * vector[46] +matrix[47][56] * vector[47] +matrix[48][56] * vector[48] +matrix[49][56] * vector[49] +matrix[50][56] * vector[50] +matrix[51][56] * vector[51] +matrix[52][56] * vector[52] +matrix[53][56] * vector[53] +matrix[54][56] * vector[54] +matrix[55][56] * vector[55] +matrix[56][56] * vector[56] +matrix[57][56] * vector[57] +matrix[58][56] * vector[58] +matrix[59][56] * vector[59] +matrix[60][56] * vector[60] +matrix[61][56] * vector[61] +matrix[62][56] * vector[62] +matrix[63][56] * vector[63] +matrix[64][56] * vector[64] +matrix[65][56] * vector[65] +matrix[66][56] * vector[66] +matrix[67][56] * vector[67] +matrix[68][56] * vector[68] +matrix[69][56] * vector[69] +matrix[70][56] * vector[70] +matrix[71][56] * vector[71] +matrix[72][56] * vector[72] +matrix[73][56] * vector[73] +matrix[74][56] * vector[74] +matrix[75][56] * vector[75] +matrix[76][56] * vector[76] +matrix[77][56] * vector[77] +matrix[78][56] * vector[78] +matrix[79][56] * vector[79] +matrix[80][56] * vector[80] +matrix[81][56] * vector[81] +matrix[82][56] * vector[82] +matrix[83][56] * vector[83] +matrix[84][56] * vector[84] +matrix[85][56] * vector[85] +matrix[86][56] * vector[86] +matrix[87][56] * vector[87] +matrix[88][56] * vector[88] +matrix[89][56] * vector[89] +matrix[90][56] * vector[90] +matrix[91][56] * vector[91] +matrix[92][56] * vector[92] +matrix[93][56] * vector[93] +matrix[94][56] * vector[94] +matrix[95][56] * vector[95] +matrix[96][56] * vector[96] +matrix[97][56] * vector[97] +matrix[98][56] * vector[98] +matrix[99][56] * vector[99] +b[56];
assign result[57] = matrix[0][57] * vector[0] +matrix[1][57] * vector[1] +matrix[2][57] * vector[2] +matrix[3][57] * vector[3] +matrix[4][57] * vector[4] +matrix[5][57] * vector[5] +matrix[6][57] * vector[6] +matrix[7][57] * vector[7] +matrix[8][57] * vector[8] +matrix[9][57] * vector[9] +matrix[10][57] * vector[10] +matrix[11][57] * vector[11] +matrix[12][57] * vector[12] +matrix[13][57] * vector[13] +matrix[14][57] * vector[14] +matrix[15][57] * vector[15] +matrix[16][57] * vector[16] +matrix[17][57] * vector[17] +matrix[18][57] * vector[18] +matrix[19][57] * vector[19] +matrix[20][57] * vector[20] +matrix[21][57] * vector[21] +matrix[22][57] * vector[22] +matrix[23][57] * vector[23] +matrix[24][57] * vector[24] +matrix[25][57] * vector[25] +matrix[26][57] * vector[26] +matrix[27][57] * vector[27] +matrix[28][57] * vector[28] +matrix[29][57] * vector[29] +matrix[30][57] * vector[30] +matrix[31][57] * vector[31] +matrix[32][57] * vector[32] +matrix[33][57] * vector[33] +matrix[34][57] * vector[34] +matrix[35][57] * vector[35] +matrix[36][57] * vector[36] +matrix[37][57] * vector[37] +matrix[38][57] * vector[38] +matrix[39][57] * vector[39] +matrix[40][57] * vector[40] +matrix[41][57] * vector[41] +matrix[42][57] * vector[42] +matrix[43][57] * vector[43] +matrix[44][57] * vector[44] +matrix[45][57] * vector[45] +matrix[46][57] * vector[46] +matrix[47][57] * vector[47] +matrix[48][57] * vector[48] +matrix[49][57] * vector[49] +matrix[50][57] * vector[50] +matrix[51][57] * vector[51] +matrix[52][57] * vector[52] +matrix[53][57] * vector[53] +matrix[54][57] * vector[54] +matrix[55][57] * vector[55] +matrix[56][57] * vector[56] +matrix[57][57] * vector[57] +matrix[58][57] * vector[58] +matrix[59][57] * vector[59] +matrix[60][57] * vector[60] +matrix[61][57] * vector[61] +matrix[62][57] * vector[62] +matrix[63][57] * vector[63] +matrix[64][57] * vector[64] +matrix[65][57] * vector[65] +matrix[66][57] * vector[66] +matrix[67][57] * vector[67] +matrix[68][57] * vector[68] +matrix[69][57] * vector[69] +matrix[70][57] * vector[70] +matrix[71][57] * vector[71] +matrix[72][57] * vector[72] +matrix[73][57] * vector[73] +matrix[74][57] * vector[74] +matrix[75][57] * vector[75] +matrix[76][57] * vector[76] +matrix[77][57] * vector[77] +matrix[78][57] * vector[78] +matrix[79][57] * vector[79] +matrix[80][57] * vector[80] +matrix[81][57] * vector[81] +matrix[82][57] * vector[82] +matrix[83][57] * vector[83] +matrix[84][57] * vector[84] +matrix[85][57] * vector[85] +matrix[86][57] * vector[86] +matrix[87][57] * vector[87] +matrix[88][57] * vector[88] +matrix[89][57] * vector[89] +matrix[90][57] * vector[90] +matrix[91][57] * vector[91] +matrix[92][57] * vector[92] +matrix[93][57] * vector[93] +matrix[94][57] * vector[94] +matrix[95][57] * vector[95] +matrix[96][57] * vector[96] +matrix[97][57] * vector[97] +matrix[98][57] * vector[98] +matrix[99][57] * vector[99] +b[57];
assign result[58] = matrix[0][58] * vector[0] +matrix[1][58] * vector[1] +matrix[2][58] * vector[2] +matrix[3][58] * vector[3] +matrix[4][58] * vector[4] +matrix[5][58] * vector[5] +matrix[6][58] * vector[6] +matrix[7][58] * vector[7] +matrix[8][58] * vector[8] +matrix[9][58] * vector[9] +matrix[10][58] * vector[10] +matrix[11][58] * vector[11] +matrix[12][58] * vector[12] +matrix[13][58] * vector[13] +matrix[14][58] * vector[14] +matrix[15][58] * vector[15] +matrix[16][58] * vector[16] +matrix[17][58] * vector[17] +matrix[18][58] * vector[18] +matrix[19][58] * vector[19] +matrix[20][58] * vector[20] +matrix[21][58] * vector[21] +matrix[22][58] * vector[22] +matrix[23][58] * vector[23] +matrix[24][58] * vector[24] +matrix[25][58] * vector[25] +matrix[26][58] * vector[26] +matrix[27][58] * vector[27] +matrix[28][58] * vector[28] +matrix[29][58] * vector[29] +matrix[30][58] * vector[30] +matrix[31][58] * vector[31] +matrix[32][58] * vector[32] +matrix[33][58] * vector[33] +matrix[34][58] * vector[34] +matrix[35][58] * vector[35] +matrix[36][58] * vector[36] +matrix[37][58] * vector[37] +matrix[38][58] * vector[38] +matrix[39][58] * vector[39] +matrix[40][58] * vector[40] +matrix[41][58] * vector[41] +matrix[42][58] * vector[42] +matrix[43][58] * vector[43] +matrix[44][58] * vector[44] +matrix[45][58] * vector[45] +matrix[46][58] * vector[46] +matrix[47][58] * vector[47] +matrix[48][58] * vector[48] +matrix[49][58] * vector[49] +matrix[50][58] * vector[50] +matrix[51][58] * vector[51] +matrix[52][58] * vector[52] +matrix[53][58] * vector[53] +matrix[54][58] * vector[54] +matrix[55][58] * vector[55] +matrix[56][58] * vector[56] +matrix[57][58] * vector[57] +matrix[58][58] * vector[58] +matrix[59][58] * vector[59] +matrix[60][58] * vector[60] +matrix[61][58] * vector[61] +matrix[62][58] * vector[62] +matrix[63][58] * vector[63] +matrix[64][58] * vector[64] +matrix[65][58] * vector[65] +matrix[66][58] * vector[66] +matrix[67][58] * vector[67] +matrix[68][58] * vector[68] +matrix[69][58] * vector[69] +matrix[70][58] * vector[70] +matrix[71][58] * vector[71] +matrix[72][58] * vector[72] +matrix[73][58] * vector[73] +matrix[74][58] * vector[74] +matrix[75][58] * vector[75] +matrix[76][58] * vector[76] +matrix[77][58] * vector[77] +matrix[78][58] * vector[78] +matrix[79][58] * vector[79] +matrix[80][58] * vector[80] +matrix[81][58] * vector[81] +matrix[82][58] * vector[82] +matrix[83][58] * vector[83] +matrix[84][58] * vector[84] +matrix[85][58] * vector[85] +matrix[86][58] * vector[86] +matrix[87][58] * vector[87] +matrix[88][58] * vector[88] +matrix[89][58] * vector[89] +matrix[90][58] * vector[90] +matrix[91][58] * vector[91] +matrix[92][58] * vector[92] +matrix[93][58] * vector[93] +matrix[94][58] * vector[94] +matrix[95][58] * vector[95] +matrix[96][58] * vector[96] +matrix[97][58] * vector[97] +matrix[98][58] * vector[98] +matrix[99][58] * vector[99] +b[58];
assign result[59] = matrix[0][59] * vector[0] +matrix[1][59] * vector[1] +matrix[2][59] * vector[2] +matrix[3][59] * vector[3] +matrix[4][59] * vector[4] +matrix[5][59] * vector[5] +matrix[6][59] * vector[6] +matrix[7][59] * vector[7] +matrix[8][59] * vector[8] +matrix[9][59] * vector[9] +matrix[10][59] * vector[10] +matrix[11][59] * vector[11] +matrix[12][59] * vector[12] +matrix[13][59] * vector[13] +matrix[14][59] * vector[14] +matrix[15][59] * vector[15] +matrix[16][59] * vector[16] +matrix[17][59] * vector[17] +matrix[18][59] * vector[18] +matrix[19][59] * vector[19] +matrix[20][59] * vector[20] +matrix[21][59] * vector[21] +matrix[22][59] * vector[22] +matrix[23][59] * vector[23] +matrix[24][59] * vector[24] +matrix[25][59] * vector[25] +matrix[26][59] * vector[26] +matrix[27][59] * vector[27] +matrix[28][59] * vector[28] +matrix[29][59] * vector[29] +matrix[30][59] * vector[30] +matrix[31][59] * vector[31] +matrix[32][59] * vector[32] +matrix[33][59] * vector[33] +matrix[34][59] * vector[34] +matrix[35][59] * vector[35] +matrix[36][59] * vector[36] +matrix[37][59] * vector[37] +matrix[38][59] * vector[38] +matrix[39][59] * vector[39] +matrix[40][59] * vector[40] +matrix[41][59] * vector[41] +matrix[42][59] * vector[42] +matrix[43][59] * vector[43] +matrix[44][59] * vector[44] +matrix[45][59] * vector[45] +matrix[46][59] * vector[46] +matrix[47][59] * vector[47] +matrix[48][59] * vector[48] +matrix[49][59] * vector[49] +matrix[50][59] * vector[50] +matrix[51][59] * vector[51] +matrix[52][59] * vector[52] +matrix[53][59] * vector[53] +matrix[54][59] * vector[54] +matrix[55][59] * vector[55] +matrix[56][59] * vector[56] +matrix[57][59] * vector[57] +matrix[58][59] * vector[58] +matrix[59][59] * vector[59] +matrix[60][59] * vector[60] +matrix[61][59] * vector[61] +matrix[62][59] * vector[62] +matrix[63][59] * vector[63] +matrix[64][59] * vector[64] +matrix[65][59] * vector[65] +matrix[66][59] * vector[66] +matrix[67][59] * vector[67] +matrix[68][59] * vector[68] +matrix[69][59] * vector[69] +matrix[70][59] * vector[70] +matrix[71][59] * vector[71] +matrix[72][59] * vector[72] +matrix[73][59] * vector[73] +matrix[74][59] * vector[74] +matrix[75][59] * vector[75] +matrix[76][59] * vector[76] +matrix[77][59] * vector[77] +matrix[78][59] * vector[78] +matrix[79][59] * vector[79] +matrix[80][59] * vector[80] +matrix[81][59] * vector[81] +matrix[82][59] * vector[82] +matrix[83][59] * vector[83] +matrix[84][59] * vector[84] +matrix[85][59] * vector[85] +matrix[86][59] * vector[86] +matrix[87][59] * vector[87] +matrix[88][59] * vector[88] +matrix[89][59] * vector[89] +matrix[90][59] * vector[90] +matrix[91][59] * vector[91] +matrix[92][59] * vector[92] +matrix[93][59] * vector[93] +matrix[94][59] * vector[94] +matrix[95][59] * vector[95] +matrix[96][59] * vector[96] +matrix[97][59] * vector[97] +matrix[98][59] * vector[98] +matrix[99][59] * vector[99] +b[59];
assign result[60] = matrix[0][60] * vector[0] +matrix[1][60] * vector[1] +matrix[2][60] * vector[2] +matrix[3][60] * vector[3] +matrix[4][60] * vector[4] +matrix[5][60] * vector[5] +matrix[6][60] * vector[6] +matrix[7][60] * vector[7] +matrix[8][60] * vector[8] +matrix[9][60] * vector[9] +matrix[10][60] * vector[10] +matrix[11][60] * vector[11] +matrix[12][60] * vector[12] +matrix[13][60] * vector[13] +matrix[14][60] * vector[14] +matrix[15][60] * vector[15] +matrix[16][60] * vector[16] +matrix[17][60] * vector[17] +matrix[18][60] * vector[18] +matrix[19][60] * vector[19] +matrix[20][60] * vector[20] +matrix[21][60] * vector[21] +matrix[22][60] * vector[22] +matrix[23][60] * vector[23] +matrix[24][60] * vector[24] +matrix[25][60] * vector[25] +matrix[26][60] * vector[26] +matrix[27][60] * vector[27] +matrix[28][60] * vector[28] +matrix[29][60] * vector[29] +matrix[30][60] * vector[30] +matrix[31][60] * vector[31] +matrix[32][60] * vector[32] +matrix[33][60] * vector[33] +matrix[34][60] * vector[34] +matrix[35][60] * vector[35] +matrix[36][60] * vector[36] +matrix[37][60] * vector[37] +matrix[38][60] * vector[38] +matrix[39][60] * vector[39] +matrix[40][60] * vector[40] +matrix[41][60] * vector[41] +matrix[42][60] * vector[42] +matrix[43][60] * vector[43] +matrix[44][60] * vector[44] +matrix[45][60] * vector[45] +matrix[46][60] * vector[46] +matrix[47][60] * vector[47] +matrix[48][60] * vector[48] +matrix[49][60] * vector[49] +matrix[50][60] * vector[50] +matrix[51][60] * vector[51] +matrix[52][60] * vector[52] +matrix[53][60] * vector[53] +matrix[54][60] * vector[54] +matrix[55][60] * vector[55] +matrix[56][60] * vector[56] +matrix[57][60] * vector[57] +matrix[58][60] * vector[58] +matrix[59][60] * vector[59] +matrix[60][60] * vector[60] +matrix[61][60] * vector[61] +matrix[62][60] * vector[62] +matrix[63][60] * vector[63] +matrix[64][60] * vector[64] +matrix[65][60] * vector[65] +matrix[66][60] * vector[66] +matrix[67][60] * vector[67] +matrix[68][60] * vector[68] +matrix[69][60] * vector[69] +matrix[70][60] * vector[70] +matrix[71][60] * vector[71] +matrix[72][60] * vector[72] +matrix[73][60] * vector[73] +matrix[74][60] * vector[74] +matrix[75][60] * vector[75] +matrix[76][60] * vector[76] +matrix[77][60] * vector[77] +matrix[78][60] * vector[78] +matrix[79][60] * vector[79] +matrix[80][60] * vector[80] +matrix[81][60] * vector[81] +matrix[82][60] * vector[82] +matrix[83][60] * vector[83] +matrix[84][60] * vector[84] +matrix[85][60] * vector[85] +matrix[86][60] * vector[86] +matrix[87][60] * vector[87] +matrix[88][60] * vector[88] +matrix[89][60] * vector[89] +matrix[90][60] * vector[90] +matrix[91][60] * vector[91] +matrix[92][60] * vector[92] +matrix[93][60] * vector[93] +matrix[94][60] * vector[94] +matrix[95][60] * vector[95] +matrix[96][60] * vector[96] +matrix[97][60] * vector[97] +matrix[98][60] * vector[98] +matrix[99][60] * vector[99] +b[60];
assign result[61] = matrix[0][61] * vector[0] +matrix[1][61] * vector[1] +matrix[2][61] * vector[2] +matrix[3][61] * vector[3] +matrix[4][61] * vector[4] +matrix[5][61] * vector[5] +matrix[6][61] * vector[6] +matrix[7][61] * vector[7] +matrix[8][61] * vector[8] +matrix[9][61] * vector[9] +matrix[10][61] * vector[10] +matrix[11][61] * vector[11] +matrix[12][61] * vector[12] +matrix[13][61] * vector[13] +matrix[14][61] * vector[14] +matrix[15][61] * vector[15] +matrix[16][61] * vector[16] +matrix[17][61] * vector[17] +matrix[18][61] * vector[18] +matrix[19][61] * vector[19] +matrix[20][61] * vector[20] +matrix[21][61] * vector[21] +matrix[22][61] * vector[22] +matrix[23][61] * vector[23] +matrix[24][61] * vector[24] +matrix[25][61] * vector[25] +matrix[26][61] * vector[26] +matrix[27][61] * vector[27] +matrix[28][61] * vector[28] +matrix[29][61] * vector[29] +matrix[30][61] * vector[30] +matrix[31][61] * vector[31] +matrix[32][61] * vector[32] +matrix[33][61] * vector[33] +matrix[34][61] * vector[34] +matrix[35][61] * vector[35] +matrix[36][61] * vector[36] +matrix[37][61] * vector[37] +matrix[38][61] * vector[38] +matrix[39][61] * vector[39] +matrix[40][61] * vector[40] +matrix[41][61] * vector[41] +matrix[42][61] * vector[42] +matrix[43][61] * vector[43] +matrix[44][61] * vector[44] +matrix[45][61] * vector[45] +matrix[46][61] * vector[46] +matrix[47][61] * vector[47] +matrix[48][61] * vector[48] +matrix[49][61] * vector[49] +matrix[50][61] * vector[50] +matrix[51][61] * vector[51] +matrix[52][61] * vector[52] +matrix[53][61] * vector[53] +matrix[54][61] * vector[54] +matrix[55][61] * vector[55] +matrix[56][61] * vector[56] +matrix[57][61] * vector[57] +matrix[58][61] * vector[58] +matrix[59][61] * vector[59] +matrix[60][61] * vector[60] +matrix[61][61] * vector[61] +matrix[62][61] * vector[62] +matrix[63][61] * vector[63] +matrix[64][61] * vector[64] +matrix[65][61] * vector[65] +matrix[66][61] * vector[66] +matrix[67][61] * vector[67] +matrix[68][61] * vector[68] +matrix[69][61] * vector[69] +matrix[70][61] * vector[70] +matrix[71][61] * vector[71] +matrix[72][61] * vector[72] +matrix[73][61] * vector[73] +matrix[74][61] * vector[74] +matrix[75][61] * vector[75] +matrix[76][61] * vector[76] +matrix[77][61] * vector[77] +matrix[78][61] * vector[78] +matrix[79][61] * vector[79] +matrix[80][61] * vector[80] +matrix[81][61] * vector[81] +matrix[82][61] * vector[82] +matrix[83][61] * vector[83] +matrix[84][61] * vector[84] +matrix[85][61] * vector[85] +matrix[86][61] * vector[86] +matrix[87][61] * vector[87] +matrix[88][61] * vector[88] +matrix[89][61] * vector[89] +matrix[90][61] * vector[90] +matrix[91][61] * vector[91] +matrix[92][61] * vector[92] +matrix[93][61] * vector[93] +matrix[94][61] * vector[94] +matrix[95][61] * vector[95] +matrix[96][61] * vector[96] +matrix[97][61] * vector[97] +matrix[98][61] * vector[98] +matrix[99][61] * vector[99] +b[61];
assign result[62] = matrix[0][62] * vector[0] +matrix[1][62] * vector[1] +matrix[2][62] * vector[2] +matrix[3][62] * vector[3] +matrix[4][62] * vector[4] +matrix[5][62] * vector[5] +matrix[6][62] * vector[6] +matrix[7][62] * vector[7] +matrix[8][62] * vector[8] +matrix[9][62] * vector[9] +matrix[10][62] * vector[10] +matrix[11][62] * vector[11] +matrix[12][62] * vector[12] +matrix[13][62] * vector[13] +matrix[14][62] * vector[14] +matrix[15][62] * vector[15] +matrix[16][62] * vector[16] +matrix[17][62] * vector[17] +matrix[18][62] * vector[18] +matrix[19][62] * vector[19] +matrix[20][62] * vector[20] +matrix[21][62] * vector[21] +matrix[22][62] * vector[22] +matrix[23][62] * vector[23] +matrix[24][62] * vector[24] +matrix[25][62] * vector[25] +matrix[26][62] * vector[26] +matrix[27][62] * vector[27] +matrix[28][62] * vector[28] +matrix[29][62] * vector[29] +matrix[30][62] * vector[30] +matrix[31][62] * vector[31] +matrix[32][62] * vector[32] +matrix[33][62] * vector[33] +matrix[34][62] * vector[34] +matrix[35][62] * vector[35] +matrix[36][62] * vector[36] +matrix[37][62] * vector[37] +matrix[38][62] * vector[38] +matrix[39][62] * vector[39] +matrix[40][62] * vector[40] +matrix[41][62] * vector[41] +matrix[42][62] * vector[42] +matrix[43][62] * vector[43] +matrix[44][62] * vector[44] +matrix[45][62] * vector[45] +matrix[46][62] * vector[46] +matrix[47][62] * vector[47] +matrix[48][62] * vector[48] +matrix[49][62] * vector[49] +matrix[50][62] * vector[50] +matrix[51][62] * vector[51] +matrix[52][62] * vector[52] +matrix[53][62] * vector[53] +matrix[54][62] * vector[54] +matrix[55][62] * vector[55] +matrix[56][62] * vector[56] +matrix[57][62] * vector[57] +matrix[58][62] * vector[58] +matrix[59][62] * vector[59] +matrix[60][62] * vector[60] +matrix[61][62] * vector[61] +matrix[62][62] * vector[62] +matrix[63][62] * vector[63] +matrix[64][62] * vector[64] +matrix[65][62] * vector[65] +matrix[66][62] * vector[66] +matrix[67][62] * vector[67] +matrix[68][62] * vector[68] +matrix[69][62] * vector[69] +matrix[70][62] * vector[70] +matrix[71][62] * vector[71] +matrix[72][62] * vector[72] +matrix[73][62] * vector[73] +matrix[74][62] * vector[74] +matrix[75][62] * vector[75] +matrix[76][62] * vector[76] +matrix[77][62] * vector[77] +matrix[78][62] * vector[78] +matrix[79][62] * vector[79] +matrix[80][62] * vector[80] +matrix[81][62] * vector[81] +matrix[82][62] * vector[82] +matrix[83][62] * vector[83] +matrix[84][62] * vector[84] +matrix[85][62] * vector[85] +matrix[86][62] * vector[86] +matrix[87][62] * vector[87] +matrix[88][62] * vector[88] +matrix[89][62] * vector[89] +matrix[90][62] * vector[90] +matrix[91][62] * vector[91] +matrix[92][62] * vector[92] +matrix[93][62] * vector[93] +matrix[94][62] * vector[94] +matrix[95][62] * vector[95] +matrix[96][62] * vector[96] +matrix[97][62] * vector[97] +matrix[98][62] * vector[98] +matrix[99][62] * vector[99] +b[62];
assign result[63] = matrix[0][63] * vector[0] +matrix[1][63] * vector[1] +matrix[2][63] * vector[2] +matrix[3][63] * vector[3] +matrix[4][63] * vector[4] +matrix[5][63] * vector[5] +matrix[6][63] * vector[6] +matrix[7][63] * vector[7] +matrix[8][63] * vector[8] +matrix[9][63] * vector[9] +matrix[10][63] * vector[10] +matrix[11][63] * vector[11] +matrix[12][63] * vector[12] +matrix[13][63] * vector[13] +matrix[14][63] * vector[14] +matrix[15][63] * vector[15] +matrix[16][63] * vector[16] +matrix[17][63] * vector[17] +matrix[18][63] * vector[18] +matrix[19][63] * vector[19] +matrix[20][63] * vector[20] +matrix[21][63] * vector[21] +matrix[22][63] * vector[22] +matrix[23][63] * vector[23] +matrix[24][63] * vector[24] +matrix[25][63] * vector[25] +matrix[26][63] * vector[26] +matrix[27][63] * vector[27] +matrix[28][63] * vector[28] +matrix[29][63] * vector[29] +matrix[30][63] * vector[30] +matrix[31][63] * vector[31] +matrix[32][63] * vector[32] +matrix[33][63] * vector[33] +matrix[34][63] * vector[34] +matrix[35][63] * vector[35] +matrix[36][63] * vector[36] +matrix[37][63] * vector[37] +matrix[38][63] * vector[38] +matrix[39][63] * vector[39] +matrix[40][63] * vector[40] +matrix[41][63] * vector[41] +matrix[42][63] * vector[42] +matrix[43][63] * vector[43] +matrix[44][63] * vector[44] +matrix[45][63] * vector[45] +matrix[46][63] * vector[46] +matrix[47][63] * vector[47] +matrix[48][63] * vector[48] +matrix[49][63] * vector[49] +matrix[50][63] * vector[50] +matrix[51][63] * vector[51] +matrix[52][63] * vector[52] +matrix[53][63] * vector[53] +matrix[54][63] * vector[54] +matrix[55][63] * vector[55] +matrix[56][63] * vector[56] +matrix[57][63] * vector[57] +matrix[58][63] * vector[58] +matrix[59][63] * vector[59] +matrix[60][63] * vector[60] +matrix[61][63] * vector[61] +matrix[62][63] * vector[62] +matrix[63][63] * vector[63] +matrix[64][63] * vector[64] +matrix[65][63] * vector[65] +matrix[66][63] * vector[66] +matrix[67][63] * vector[67] +matrix[68][63] * vector[68] +matrix[69][63] * vector[69] +matrix[70][63] * vector[70] +matrix[71][63] * vector[71] +matrix[72][63] * vector[72] +matrix[73][63] * vector[73] +matrix[74][63] * vector[74] +matrix[75][63] * vector[75] +matrix[76][63] * vector[76] +matrix[77][63] * vector[77] +matrix[78][63] * vector[78] +matrix[79][63] * vector[79] +matrix[80][63] * vector[80] +matrix[81][63] * vector[81] +matrix[82][63] * vector[82] +matrix[83][63] * vector[83] +matrix[84][63] * vector[84] +matrix[85][63] * vector[85] +matrix[86][63] * vector[86] +matrix[87][63] * vector[87] +matrix[88][63] * vector[88] +matrix[89][63] * vector[89] +matrix[90][63] * vector[90] +matrix[91][63] * vector[91] +matrix[92][63] * vector[92] +matrix[93][63] * vector[93] +matrix[94][63] * vector[94] +matrix[95][63] * vector[95] +matrix[96][63] * vector[96] +matrix[97][63] * vector[97] +matrix[98][63] * vector[98] +matrix[99][63] * vector[99] +b[63];
assign result[64] = matrix[0][64] * vector[0] +matrix[1][64] * vector[1] +matrix[2][64] * vector[2] +matrix[3][64] * vector[3] +matrix[4][64] * vector[4] +matrix[5][64] * vector[5] +matrix[6][64] * vector[6] +matrix[7][64] * vector[7] +matrix[8][64] * vector[8] +matrix[9][64] * vector[9] +matrix[10][64] * vector[10] +matrix[11][64] * vector[11] +matrix[12][64] * vector[12] +matrix[13][64] * vector[13] +matrix[14][64] * vector[14] +matrix[15][64] * vector[15] +matrix[16][64] * vector[16] +matrix[17][64] * vector[17] +matrix[18][64] * vector[18] +matrix[19][64] * vector[19] +matrix[20][64] * vector[20] +matrix[21][64] * vector[21] +matrix[22][64] * vector[22] +matrix[23][64] * vector[23] +matrix[24][64] * vector[24] +matrix[25][64] * vector[25] +matrix[26][64] * vector[26] +matrix[27][64] * vector[27] +matrix[28][64] * vector[28] +matrix[29][64] * vector[29] +matrix[30][64] * vector[30] +matrix[31][64] * vector[31] +matrix[32][64] * vector[32] +matrix[33][64] * vector[33] +matrix[34][64] * vector[34] +matrix[35][64] * vector[35] +matrix[36][64] * vector[36] +matrix[37][64] * vector[37] +matrix[38][64] * vector[38] +matrix[39][64] * vector[39] +matrix[40][64] * vector[40] +matrix[41][64] * vector[41] +matrix[42][64] * vector[42] +matrix[43][64] * vector[43] +matrix[44][64] * vector[44] +matrix[45][64] * vector[45] +matrix[46][64] * vector[46] +matrix[47][64] * vector[47] +matrix[48][64] * vector[48] +matrix[49][64] * vector[49] +matrix[50][64] * vector[50] +matrix[51][64] * vector[51] +matrix[52][64] * vector[52] +matrix[53][64] * vector[53] +matrix[54][64] * vector[54] +matrix[55][64] * vector[55] +matrix[56][64] * vector[56] +matrix[57][64] * vector[57] +matrix[58][64] * vector[58] +matrix[59][64] * vector[59] +matrix[60][64] * vector[60] +matrix[61][64] * vector[61] +matrix[62][64] * vector[62] +matrix[63][64] * vector[63] +matrix[64][64] * vector[64] +matrix[65][64] * vector[65] +matrix[66][64] * vector[66] +matrix[67][64] * vector[67] +matrix[68][64] * vector[68] +matrix[69][64] * vector[69] +matrix[70][64] * vector[70] +matrix[71][64] * vector[71] +matrix[72][64] * vector[72] +matrix[73][64] * vector[73] +matrix[74][64] * vector[74] +matrix[75][64] * vector[75] +matrix[76][64] * vector[76] +matrix[77][64] * vector[77] +matrix[78][64] * vector[78] +matrix[79][64] * vector[79] +matrix[80][64] * vector[80] +matrix[81][64] * vector[81] +matrix[82][64] * vector[82] +matrix[83][64] * vector[83] +matrix[84][64] * vector[84] +matrix[85][64] * vector[85] +matrix[86][64] * vector[86] +matrix[87][64] * vector[87] +matrix[88][64] * vector[88] +matrix[89][64] * vector[89] +matrix[90][64] * vector[90] +matrix[91][64] * vector[91] +matrix[92][64] * vector[92] +matrix[93][64] * vector[93] +matrix[94][64] * vector[94] +matrix[95][64] * vector[95] +matrix[96][64] * vector[96] +matrix[97][64] * vector[97] +matrix[98][64] * vector[98] +matrix[99][64] * vector[99] +b[64];
assign result[65] = matrix[0][65] * vector[0] +matrix[1][65] * vector[1] +matrix[2][65] * vector[2] +matrix[3][65] * vector[3] +matrix[4][65] * vector[4] +matrix[5][65] * vector[5] +matrix[6][65] * vector[6] +matrix[7][65] * vector[7] +matrix[8][65] * vector[8] +matrix[9][65] * vector[9] +matrix[10][65] * vector[10] +matrix[11][65] * vector[11] +matrix[12][65] * vector[12] +matrix[13][65] * vector[13] +matrix[14][65] * vector[14] +matrix[15][65] * vector[15] +matrix[16][65] * vector[16] +matrix[17][65] * vector[17] +matrix[18][65] * vector[18] +matrix[19][65] * vector[19] +matrix[20][65] * vector[20] +matrix[21][65] * vector[21] +matrix[22][65] * vector[22] +matrix[23][65] * vector[23] +matrix[24][65] * vector[24] +matrix[25][65] * vector[25] +matrix[26][65] * vector[26] +matrix[27][65] * vector[27] +matrix[28][65] * vector[28] +matrix[29][65] * vector[29] +matrix[30][65] * vector[30] +matrix[31][65] * vector[31] +matrix[32][65] * vector[32] +matrix[33][65] * vector[33] +matrix[34][65] * vector[34] +matrix[35][65] * vector[35] +matrix[36][65] * vector[36] +matrix[37][65] * vector[37] +matrix[38][65] * vector[38] +matrix[39][65] * vector[39] +matrix[40][65] * vector[40] +matrix[41][65] * vector[41] +matrix[42][65] * vector[42] +matrix[43][65] * vector[43] +matrix[44][65] * vector[44] +matrix[45][65] * vector[45] +matrix[46][65] * vector[46] +matrix[47][65] * vector[47] +matrix[48][65] * vector[48] +matrix[49][65] * vector[49] +matrix[50][65] * vector[50] +matrix[51][65] * vector[51] +matrix[52][65] * vector[52] +matrix[53][65] * vector[53] +matrix[54][65] * vector[54] +matrix[55][65] * vector[55] +matrix[56][65] * vector[56] +matrix[57][65] * vector[57] +matrix[58][65] * vector[58] +matrix[59][65] * vector[59] +matrix[60][65] * vector[60] +matrix[61][65] * vector[61] +matrix[62][65] * vector[62] +matrix[63][65] * vector[63] +matrix[64][65] * vector[64] +matrix[65][65] * vector[65] +matrix[66][65] * vector[66] +matrix[67][65] * vector[67] +matrix[68][65] * vector[68] +matrix[69][65] * vector[69] +matrix[70][65] * vector[70] +matrix[71][65] * vector[71] +matrix[72][65] * vector[72] +matrix[73][65] * vector[73] +matrix[74][65] * vector[74] +matrix[75][65] * vector[75] +matrix[76][65] * vector[76] +matrix[77][65] * vector[77] +matrix[78][65] * vector[78] +matrix[79][65] * vector[79] +matrix[80][65] * vector[80] +matrix[81][65] * vector[81] +matrix[82][65] * vector[82] +matrix[83][65] * vector[83] +matrix[84][65] * vector[84] +matrix[85][65] * vector[85] +matrix[86][65] * vector[86] +matrix[87][65] * vector[87] +matrix[88][65] * vector[88] +matrix[89][65] * vector[89] +matrix[90][65] * vector[90] +matrix[91][65] * vector[91] +matrix[92][65] * vector[92] +matrix[93][65] * vector[93] +matrix[94][65] * vector[94] +matrix[95][65] * vector[95] +matrix[96][65] * vector[96] +matrix[97][65] * vector[97] +matrix[98][65] * vector[98] +matrix[99][65] * vector[99] +b[65];
assign result[66] = matrix[0][66] * vector[0] +matrix[1][66] * vector[1] +matrix[2][66] * vector[2] +matrix[3][66] * vector[3] +matrix[4][66] * vector[4] +matrix[5][66] * vector[5] +matrix[6][66] * vector[6] +matrix[7][66] * vector[7] +matrix[8][66] * vector[8] +matrix[9][66] * vector[9] +matrix[10][66] * vector[10] +matrix[11][66] * vector[11] +matrix[12][66] * vector[12] +matrix[13][66] * vector[13] +matrix[14][66] * vector[14] +matrix[15][66] * vector[15] +matrix[16][66] * vector[16] +matrix[17][66] * vector[17] +matrix[18][66] * vector[18] +matrix[19][66] * vector[19] +matrix[20][66] * vector[20] +matrix[21][66] * vector[21] +matrix[22][66] * vector[22] +matrix[23][66] * vector[23] +matrix[24][66] * vector[24] +matrix[25][66] * vector[25] +matrix[26][66] * vector[26] +matrix[27][66] * vector[27] +matrix[28][66] * vector[28] +matrix[29][66] * vector[29] +matrix[30][66] * vector[30] +matrix[31][66] * vector[31] +matrix[32][66] * vector[32] +matrix[33][66] * vector[33] +matrix[34][66] * vector[34] +matrix[35][66] * vector[35] +matrix[36][66] * vector[36] +matrix[37][66] * vector[37] +matrix[38][66] * vector[38] +matrix[39][66] * vector[39] +matrix[40][66] * vector[40] +matrix[41][66] * vector[41] +matrix[42][66] * vector[42] +matrix[43][66] * vector[43] +matrix[44][66] * vector[44] +matrix[45][66] * vector[45] +matrix[46][66] * vector[46] +matrix[47][66] * vector[47] +matrix[48][66] * vector[48] +matrix[49][66] * vector[49] +matrix[50][66] * vector[50] +matrix[51][66] * vector[51] +matrix[52][66] * vector[52] +matrix[53][66] * vector[53] +matrix[54][66] * vector[54] +matrix[55][66] * vector[55] +matrix[56][66] * vector[56] +matrix[57][66] * vector[57] +matrix[58][66] * vector[58] +matrix[59][66] * vector[59] +matrix[60][66] * vector[60] +matrix[61][66] * vector[61] +matrix[62][66] * vector[62] +matrix[63][66] * vector[63] +matrix[64][66] * vector[64] +matrix[65][66] * vector[65] +matrix[66][66] * vector[66] +matrix[67][66] * vector[67] +matrix[68][66] * vector[68] +matrix[69][66] * vector[69] +matrix[70][66] * vector[70] +matrix[71][66] * vector[71] +matrix[72][66] * vector[72] +matrix[73][66] * vector[73] +matrix[74][66] * vector[74] +matrix[75][66] * vector[75] +matrix[76][66] * vector[76] +matrix[77][66] * vector[77] +matrix[78][66] * vector[78] +matrix[79][66] * vector[79] +matrix[80][66] * vector[80] +matrix[81][66] * vector[81] +matrix[82][66] * vector[82] +matrix[83][66] * vector[83] +matrix[84][66] * vector[84] +matrix[85][66] * vector[85] +matrix[86][66] * vector[86] +matrix[87][66] * vector[87] +matrix[88][66] * vector[88] +matrix[89][66] * vector[89] +matrix[90][66] * vector[90] +matrix[91][66] * vector[91] +matrix[92][66] * vector[92] +matrix[93][66] * vector[93] +matrix[94][66] * vector[94] +matrix[95][66] * vector[95] +matrix[96][66] * vector[96] +matrix[97][66] * vector[97] +matrix[98][66] * vector[98] +matrix[99][66] * vector[99] +b[66];
assign result[67] = matrix[0][67] * vector[0] +matrix[1][67] * vector[1] +matrix[2][67] * vector[2] +matrix[3][67] * vector[3] +matrix[4][67] * vector[4] +matrix[5][67] * vector[5] +matrix[6][67] * vector[6] +matrix[7][67] * vector[7] +matrix[8][67] * vector[8] +matrix[9][67] * vector[9] +matrix[10][67] * vector[10] +matrix[11][67] * vector[11] +matrix[12][67] * vector[12] +matrix[13][67] * vector[13] +matrix[14][67] * vector[14] +matrix[15][67] * vector[15] +matrix[16][67] * vector[16] +matrix[17][67] * vector[17] +matrix[18][67] * vector[18] +matrix[19][67] * vector[19] +matrix[20][67] * vector[20] +matrix[21][67] * vector[21] +matrix[22][67] * vector[22] +matrix[23][67] * vector[23] +matrix[24][67] * vector[24] +matrix[25][67] * vector[25] +matrix[26][67] * vector[26] +matrix[27][67] * vector[27] +matrix[28][67] * vector[28] +matrix[29][67] * vector[29] +matrix[30][67] * vector[30] +matrix[31][67] * vector[31] +matrix[32][67] * vector[32] +matrix[33][67] * vector[33] +matrix[34][67] * vector[34] +matrix[35][67] * vector[35] +matrix[36][67] * vector[36] +matrix[37][67] * vector[37] +matrix[38][67] * vector[38] +matrix[39][67] * vector[39] +matrix[40][67] * vector[40] +matrix[41][67] * vector[41] +matrix[42][67] * vector[42] +matrix[43][67] * vector[43] +matrix[44][67] * vector[44] +matrix[45][67] * vector[45] +matrix[46][67] * vector[46] +matrix[47][67] * vector[47] +matrix[48][67] * vector[48] +matrix[49][67] * vector[49] +matrix[50][67] * vector[50] +matrix[51][67] * vector[51] +matrix[52][67] * vector[52] +matrix[53][67] * vector[53] +matrix[54][67] * vector[54] +matrix[55][67] * vector[55] +matrix[56][67] * vector[56] +matrix[57][67] * vector[57] +matrix[58][67] * vector[58] +matrix[59][67] * vector[59] +matrix[60][67] * vector[60] +matrix[61][67] * vector[61] +matrix[62][67] * vector[62] +matrix[63][67] * vector[63] +matrix[64][67] * vector[64] +matrix[65][67] * vector[65] +matrix[66][67] * vector[66] +matrix[67][67] * vector[67] +matrix[68][67] * vector[68] +matrix[69][67] * vector[69] +matrix[70][67] * vector[70] +matrix[71][67] * vector[71] +matrix[72][67] * vector[72] +matrix[73][67] * vector[73] +matrix[74][67] * vector[74] +matrix[75][67] * vector[75] +matrix[76][67] * vector[76] +matrix[77][67] * vector[77] +matrix[78][67] * vector[78] +matrix[79][67] * vector[79] +matrix[80][67] * vector[80] +matrix[81][67] * vector[81] +matrix[82][67] * vector[82] +matrix[83][67] * vector[83] +matrix[84][67] * vector[84] +matrix[85][67] * vector[85] +matrix[86][67] * vector[86] +matrix[87][67] * vector[87] +matrix[88][67] * vector[88] +matrix[89][67] * vector[89] +matrix[90][67] * vector[90] +matrix[91][67] * vector[91] +matrix[92][67] * vector[92] +matrix[93][67] * vector[93] +matrix[94][67] * vector[94] +matrix[95][67] * vector[95] +matrix[96][67] * vector[96] +matrix[97][67] * vector[97] +matrix[98][67] * vector[98] +matrix[99][67] * vector[99] +b[67];
assign result[68] = matrix[0][68] * vector[0] +matrix[1][68] * vector[1] +matrix[2][68] * vector[2] +matrix[3][68] * vector[3] +matrix[4][68] * vector[4] +matrix[5][68] * vector[5] +matrix[6][68] * vector[6] +matrix[7][68] * vector[7] +matrix[8][68] * vector[8] +matrix[9][68] * vector[9] +matrix[10][68] * vector[10] +matrix[11][68] * vector[11] +matrix[12][68] * vector[12] +matrix[13][68] * vector[13] +matrix[14][68] * vector[14] +matrix[15][68] * vector[15] +matrix[16][68] * vector[16] +matrix[17][68] * vector[17] +matrix[18][68] * vector[18] +matrix[19][68] * vector[19] +matrix[20][68] * vector[20] +matrix[21][68] * vector[21] +matrix[22][68] * vector[22] +matrix[23][68] * vector[23] +matrix[24][68] * vector[24] +matrix[25][68] * vector[25] +matrix[26][68] * vector[26] +matrix[27][68] * vector[27] +matrix[28][68] * vector[28] +matrix[29][68] * vector[29] +matrix[30][68] * vector[30] +matrix[31][68] * vector[31] +matrix[32][68] * vector[32] +matrix[33][68] * vector[33] +matrix[34][68] * vector[34] +matrix[35][68] * vector[35] +matrix[36][68] * vector[36] +matrix[37][68] * vector[37] +matrix[38][68] * vector[38] +matrix[39][68] * vector[39] +matrix[40][68] * vector[40] +matrix[41][68] * vector[41] +matrix[42][68] * vector[42] +matrix[43][68] * vector[43] +matrix[44][68] * vector[44] +matrix[45][68] * vector[45] +matrix[46][68] * vector[46] +matrix[47][68] * vector[47] +matrix[48][68] * vector[48] +matrix[49][68] * vector[49] +matrix[50][68] * vector[50] +matrix[51][68] * vector[51] +matrix[52][68] * vector[52] +matrix[53][68] * vector[53] +matrix[54][68] * vector[54] +matrix[55][68] * vector[55] +matrix[56][68] * vector[56] +matrix[57][68] * vector[57] +matrix[58][68] * vector[58] +matrix[59][68] * vector[59] +matrix[60][68] * vector[60] +matrix[61][68] * vector[61] +matrix[62][68] * vector[62] +matrix[63][68] * vector[63] +matrix[64][68] * vector[64] +matrix[65][68] * vector[65] +matrix[66][68] * vector[66] +matrix[67][68] * vector[67] +matrix[68][68] * vector[68] +matrix[69][68] * vector[69] +matrix[70][68] * vector[70] +matrix[71][68] * vector[71] +matrix[72][68] * vector[72] +matrix[73][68] * vector[73] +matrix[74][68] * vector[74] +matrix[75][68] * vector[75] +matrix[76][68] * vector[76] +matrix[77][68] * vector[77] +matrix[78][68] * vector[78] +matrix[79][68] * vector[79] +matrix[80][68] * vector[80] +matrix[81][68] * vector[81] +matrix[82][68] * vector[82] +matrix[83][68] * vector[83] +matrix[84][68] * vector[84] +matrix[85][68] * vector[85] +matrix[86][68] * vector[86] +matrix[87][68] * vector[87] +matrix[88][68] * vector[88] +matrix[89][68] * vector[89] +matrix[90][68] * vector[90] +matrix[91][68] * vector[91] +matrix[92][68] * vector[92] +matrix[93][68] * vector[93] +matrix[94][68] * vector[94] +matrix[95][68] * vector[95] +matrix[96][68] * vector[96] +matrix[97][68] * vector[97] +matrix[98][68] * vector[98] +matrix[99][68] * vector[99] +b[68];
assign result[69] = matrix[0][69] * vector[0] +matrix[1][69] * vector[1] +matrix[2][69] * vector[2] +matrix[3][69] * vector[3] +matrix[4][69] * vector[4] +matrix[5][69] * vector[5] +matrix[6][69] * vector[6] +matrix[7][69] * vector[7] +matrix[8][69] * vector[8] +matrix[9][69] * vector[9] +matrix[10][69] * vector[10] +matrix[11][69] * vector[11] +matrix[12][69] * vector[12] +matrix[13][69] * vector[13] +matrix[14][69] * vector[14] +matrix[15][69] * vector[15] +matrix[16][69] * vector[16] +matrix[17][69] * vector[17] +matrix[18][69] * vector[18] +matrix[19][69] * vector[19] +matrix[20][69] * vector[20] +matrix[21][69] * vector[21] +matrix[22][69] * vector[22] +matrix[23][69] * vector[23] +matrix[24][69] * vector[24] +matrix[25][69] * vector[25] +matrix[26][69] * vector[26] +matrix[27][69] * vector[27] +matrix[28][69] * vector[28] +matrix[29][69] * vector[29] +matrix[30][69] * vector[30] +matrix[31][69] * vector[31] +matrix[32][69] * vector[32] +matrix[33][69] * vector[33] +matrix[34][69] * vector[34] +matrix[35][69] * vector[35] +matrix[36][69] * vector[36] +matrix[37][69] * vector[37] +matrix[38][69] * vector[38] +matrix[39][69] * vector[39] +matrix[40][69] * vector[40] +matrix[41][69] * vector[41] +matrix[42][69] * vector[42] +matrix[43][69] * vector[43] +matrix[44][69] * vector[44] +matrix[45][69] * vector[45] +matrix[46][69] * vector[46] +matrix[47][69] * vector[47] +matrix[48][69] * vector[48] +matrix[49][69] * vector[49] +matrix[50][69] * vector[50] +matrix[51][69] * vector[51] +matrix[52][69] * vector[52] +matrix[53][69] * vector[53] +matrix[54][69] * vector[54] +matrix[55][69] * vector[55] +matrix[56][69] * vector[56] +matrix[57][69] * vector[57] +matrix[58][69] * vector[58] +matrix[59][69] * vector[59] +matrix[60][69] * vector[60] +matrix[61][69] * vector[61] +matrix[62][69] * vector[62] +matrix[63][69] * vector[63] +matrix[64][69] * vector[64] +matrix[65][69] * vector[65] +matrix[66][69] * vector[66] +matrix[67][69] * vector[67] +matrix[68][69] * vector[68] +matrix[69][69] * vector[69] +matrix[70][69] * vector[70] +matrix[71][69] * vector[71] +matrix[72][69] * vector[72] +matrix[73][69] * vector[73] +matrix[74][69] * vector[74] +matrix[75][69] * vector[75] +matrix[76][69] * vector[76] +matrix[77][69] * vector[77] +matrix[78][69] * vector[78] +matrix[79][69] * vector[79] +matrix[80][69] * vector[80] +matrix[81][69] * vector[81] +matrix[82][69] * vector[82] +matrix[83][69] * vector[83] +matrix[84][69] * vector[84] +matrix[85][69] * vector[85] +matrix[86][69] * vector[86] +matrix[87][69] * vector[87] +matrix[88][69] * vector[88] +matrix[89][69] * vector[89] +matrix[90][69] * vector[90] +matrix[91][69] * vector[91] +matrix[92][69] * vector[92] +matrix[93][69] * vector[93] +matrix[94][69] * vector[94] +matrix[95][69] * vector[95] +matrix[96][69] * vector[96] +matrix[97][69] * vector[97] +matrix[98][69] * vector[98] +matrix[99][69] * vector[99] +b[69];
assign result[70] = matrix[0][70] * vector[0] +matrix[1][70] * vector[1] +matrix[2][70] * vector[2] +matrix[3][70] * vector[3] +matrix[4][70] * vector[4] +matrix[5][70] * vector[5] +matrix[6][70] * vector[6] +matrix[7][70] * vector[7] +matrix[8][70] * vector[8] +matrix[9][70] * vector[9] +matrix[10][70] * vector[10] +matrix[11][70] * vector[11] +matrix[12][70] * vector[12] +matrix[13][70] * vector[13] +matrix[14][70] * vector[14] +matrix[15][70] * vector[15] +matrix[16][70] * vector[16] +matrix[17][70] * vector[17] +matrix[18][70] * vector[18] +matrix[19][70] * vector[19] +matrix[20][70] * vector[20] +matrix[21][70] * vector[21] +matrix[22][70] * vector[22] +matrix[23][70] * vector[23] +matrix[24][70] * vector[24] +matrix[25][70] * vector[25] +matrix[26][70] * vector[26] +matrix[27][70] * vector[27] +matrix[28][70] * vector[28] +matrix[29][70] * vector[29] +matrix[30][70] * vector[30] +matrix[31][70] * vector[31] +matrix[32][70] * vector[32] +matrix[33][70] * vector[33] +matrix[34][70] * vector[34] +matrix[35][70] * vector[35] +matrix[36][70] * vector[36] +matrix[37][70] * vector[37] +matrix[38][70] * vector[38] +matrix[39][70] * vector[39] +matrix[40][70] * vector[40] +matrix[41][70] * vector[41] +matrix[42][70] * vector[42] +matrix[43][70] * vector[43] +matrix[44][70] * vector[44] +matrix[45][70] * vector[45] +matrix[46][70] * vector[46] +matrix[47][70] * vector[47] +matrix[48][70] * vector[48] +matrix[49][70] * vector[49] +matrix[50][70] * vector[50] +matrix[51][70] * vector[51] +matrix[52][70] * vector[52] +matrix[53][70] * vector[53] +matrix[54][70] * vector[54] +matrix[55][70] * vector[55] +matrix[56][70] * vector[56] +matrix[57][70] * vector[57] +matrix[58][70] * vector[58] +matrix[59][70] * vector[59] +matrix[60][70] * vector[60] +matrix[61][70] * vector[61] +matrix[62][70] * vector[62] +matrix[63][70] * vector[63] +matrix[64][70] * vector[64] +matrix[65][70] * vector[65] +matrix[66][70] * vector[66] +matrix[67][70] * vector[67] +matrix[68][70] * vector[68] +matrix[69][70] * vector[69] +matrix[70][70] * vector[70] +matrix[71][70] * vector[71] +matrix[72][70] * vector[72] +matrix[73][70] * vector[73] +matrix[74][70] * vector[74] +matrix[75][70] * vector[75] +matrix[76][70] * vector[76] +matrix[77][70] * vector[77] +matrix[78][70] * vector[78] +matrix[79][70] * vector[79] +matrix[80][70] * vector[80] +matrix[81][70] * vector[81] +matrix[82][70] * vector[82] +matrix[83][70] * vector[83] +matrix[84][70] * vector[84] +matrix[85][70] * vector[85] +matrix[86][70] * vector[86] +matrix[87][70] * vector[87] +matrix[88][70] * vector[88] +matrix[89][70] * vector[89] +matrix[90][70] * vector[90] +matrix[91][70] * vector[91] +matrix[92][70] * vector[92] +matrix[93][70] * vector[93] +matrix[94][70] * vector[94] +matrix[95][70] * vector[95] +matrix[96][70] * vector[96] +matrix[97][70] * vector[97] +matrix[98][70] * vector[98] +matrix[99][70] * vector[99] +b[70];
assign result[71] = matrix[0][71] * vector[0] +matrix[1][71] * vector[1] +matrix[2][71] * vector[2] +matrix[3][71] * vector[3] +matrix[4][71] * vector[4] +matrix[5][71] * vector[5] +matrix[6][71] * vector[6] +matrix[7][71] * vector[7] +matrix[8][71] * vector[8] +matrix[9][71] * vector[9] +matrix[10][71] * vector[10] +matrix[11][71] * vector[11] +matrix[12][71] * vector[12] +matrix[13][71] * vector[13] +matrix[14][71] * vector[14] +matrix[15][71] * vector[15] +matrix[16][71] * vector[16] +matrix[17][71] * vector[17] +matrix[18][71] * vector[18] +matrix[19][71] * vector[19] +matrix[20][71] * vector[20] +matrix[21][71] * vector[21] +matrix[22][71] * vector[22] +matrix[23][71] * vector[23] +matrix[24][71] * vector[24] +matrix[25][71] * vector[25] +matrix[26][71] * vector[26] +matrix[27][71] * vector[27] +matrix[28][71] * vector[28] +matrix[29][71] * vector[29] +matrix[30][71] * vector[30] +matrix[31][71] * vector[31] +matrix[32][71] * vector[32] +matrix[33][71] * vector[33] +matrix[34][71] * vector[34] +matrix[35][71] * vector[35] +matrix[36][71] * vector[36] +matrix[37][71] * vector[37] +matrix[38][71] * vector[38] +matrix[39][71] * vector[39] +matrix[40][71] * vector[40] +matrix[41][71] * vector[41] +matrix[42][71] * vector[42] +matrix[43][71] * vector[43] +matrix[44][71] * vector[44] +matrix[45][71] * vector[45] +matrix[46][71] * vector[46] +matrix[47][71] * vector[47] +matrix[48][71] * vector[48] +matrix[49][71] * vector[49] +matrix[50][71] * vector[50] +matrix[51][71] * vector[51] +matrix[52][71] * vector[52] +matrix[53][71] * vector[53] +matrix[54][71] * vector[54] +matrix[55][71] * vector[55] +matrix[56][71] * vector[56] +matrix[57][71] * vector[57] +matrix[58][71] * vector[58] +matrix[59][71] * vector[59] +matrix[60][71] * vector[60] +matrix[61][71] * vector[61] +matrix[62][71] * vector[62] +matrix[63][71] * vector[63] +matrix[64][71] * vector[64] +matrix[65][71] * vector[65] +matrix[66][71] * vector[66] +matrix[67][71] * vector[67] +matrix[68][71] * vector[68] +matrix[69][71] * vector[69] +matrix[70][71] * vector[70] +matrix[71][71] * vector[71] +matrix[72][71] * vector[72] +matrix[73][71] * vector[73] +matrix[74][71] * vector[74] +matrix[75][71] * vector[75] +matrix[76][71] * vector[76] +matrix[77][71] * vector[77] +matrix[78][71] * vector[78] +matrix[79][71] * vector[79] +matrix[80][71] * vector[80] +matrix[81][71] * vector[81] +matrix[82][71] * vector[82] +matrix[83][71] * vector[83] +matrix[84][71] * vector[84] +matrix[85][71] * vector[85] +matrix[86][71] * vector[86] +matrix[87][71] * vector[87] +matrix[88][71] * vector[88] +matrix[89][71] * vector[89] +matrix[90][71] * vector[90] +matrix[91][71] * vector[91] +matrix[92][71] * vector[92] +matrix[93][71] * vector[93] +matrix[94][71] * vector[94] +matrix[95][71] * vector[95] +matrix[96][71] * vector[96] +matrix[97][71] * vector[97] +matrix[98][71] * vector[98] +matrix[99][71] * vector[99] +b[71];
assign result[72] = matrix[0][72] * vector[0] +matrix[1][72] * vector[1] +matrix[2][72] * vector[2] +matrix[3][72] * vector[3] +matrix[4][72] * vector[4] +matrix[5][72] * vector[5] +matrix[6][72] * vector[6] +matrix[7][72] * vector[7] +matrix[8][72] * vector[8] +matrix[9][72] * vector[9] +matrix[10][72] * vector[10] +matrix[11][72] * vector[11] +matrix[12][72] * vector[12] +matrix[13][72] * vector[13] +matrix[14][72] * vector[14] +matrix[15][72] * vector[15] +matrix[16][72] * vector[16] +matrix[17][72] * vector[17] +matrix[18][72] * vector[18] +matrix[19][72] * vector[19] +matrix[20][72] * vector[20] +matrix[21][72] * vector[21] +matrix[22][72] * vector[22] +matrix[23][72] * vector[23] +matrix[24][72] * vector[24] +matrix[25][72] * vector[25] +matrix[26][72] * vector[26] +matrix[27][72] * vector[27] +matrix[28][72] * vector[28] +matrix[29][72] * vector[29] +matrix[30][72] * vector[30] +matrix[31][72] * vector[31] +matrix[32][72] * vector[32] +matrix[33][72] * vector[33] +matrix[34][72] * vector[34] +matrix[35][72] * vector[35] +matrix[36][72] * vector[36] +matrix[37][72] * vector[37] +matrix[38][72] * vector[38] +matrix[39][72] * vector[39] +matrix[40][72] * vector[40] +matrix[41][72] * vector[41] +matrix[42][72] * vector[42] +matrix[43][72] * vector[43] +matrix[44][72] * vector[44] +matrix[45][72] * vector[45] +matrix[46][72] * vector[46] +matrix[47][72] * vector[47] +matrix[48][72] * vector[48] +matrix[49][72] * vector[49] +matrix[50][72] * vector[50] +matrix[51][72] * vector[51] +matrix[52][72] * vector[52] +matrix[53][72] * vector[53] +matrix[54][72] * vector[54] +matrix[55][72] * vector[55] +matrix[56][72] * vector[56] +matrix[57][72] * vector[57] +matrix[58][72] * vector[58] +matrix[59][72] * vector[59] +matrix[60][72] * vector[60] +matrix[61][72] * vector[61] +matrix[62][72] * vector[62] +matrix[63][72] * vector[63] +matrix[64][72] * vector[64] +matrix[65][72] * vector[65] +matrix[66][72] * vector[66] +matrix[67][72] * vector[67] +matrix[68][72] * vector[68] +matrix[69][72] * vector[69] +matrix[70][72] * vector[70] +matrix[71][72] * vector[71] +matrix[72][72] * vector[72] +matrix[73][72] * vector[73] +matrix[74][72] * vector[74] +matrix[75][72] * vector[75] +matrix[76][72] * vector[76] +matrix[77][72] * vector[77] +matrix[78][72] * vector[78] +matrix[79][72] * vector[79] +matrix[80][72] * vector[80] +matrix[81][72] * vector[81] +matrix[82][72] * vector[82] +matrix[83][72] * vector[83] +matrix[84][72] * vector[84] +matrix[85][72] * vector[85] +matrix[86][72] * vector[86] +matrix[87][72] * vector[87] +matrix[88][72] * vector[88] +matrix[89][72] * vector[89] +matrix[90][72] * vector[90] +matrix[91][72] * vector[91] +matrix[92][72] * vector[92] +matrix[93][72] * vector[93] +matrix[94][72] * vector[94] +matrix[95][72] * vector[95] +matrix[96][72] * vector[96] +matrix[97][72] * vector[97] +matrix[98][72] * vector[98] +matrix[99][72] * vector[99] +b[72];
assign result[73] = matrix[0][73] * vector[0] +matrix[1][73] * vector[1] +matrix[2][73] * vector[2] +matrix[3][73] * vector[3] +matrix[4][73] * vector[4] +matrix[5][73] * vector[5] +matrix[6][73] * vector[6] +matrix[7][73] * vector[7] +matrix[8][73] * vector[8] +matrix[9][73] * vector[9] +matrix[10][73] * vector[10] +matrix[11][73] * vector[11] +matrix[12][73] * vector[12] +matrix[13][73] * vector[13] +matrix[14][73] * vector[14] +matrix[15][73] * vector[15] +matrix[16][73] * vector[16] +matrix[17][73] * vector[17] +matrix[18][73] * vector[18] +matrix[19][73] * vector[19] +matrix[20][73] * vector[20] +matrix[21][73] * vector[21] +matrix[22][73] * vector[22] +matrix[23][73] * vector[23] +matrix[24][73] * vector[24] +matrix[25][73] * vector[25] +matrix[26][73] * vector[26] +matrix[27][73] * vector[27] +matrix[28][73] * vector[28] +matrix[29][73] * vector[29] +matrix[30][73] * vector[30] +matrix[31][73] * vector[31] +matrix[32][73] * vector[32] +matrix[33][73] * vector[33] +matrix[34][73] * vector[34] +matrix[35][73] * vector[35] +matrix[36][73] * vector[36] +matrix[37][73] * vector[37] +matrix[38][73] * vector[38] +matrix[39][73] * vector[39] +matrix[40][73] * vector[40] +matrix[41][73] * vector[41] +matrix[42][73] * vector[42] +matrix[43][73] * vector[43] +matrix[44][73] * vector[44] +matrix[45][73] * vector[45] +matrix[46][73] * vector[46] +matrix[47][73] * vector[47] +matrix[48][73] * vector[48] +matrix[49][73] * vector[49] +matrix[50][73] * vector[50] +matrix[51][73] * vector[51] +matrix[52][73] * vector[52] +matrix[53][73] * vector[53] +matrix[54][73] * vector[54] +matrix[55][73] * vector[55] +matrix[56][73] * vector[56] +matrix[57][73] * vector[57] +matrix[58][73] * vector[58] +matrix[59][73] * vector[59] +matrix[60][73] * vector[60] +matrix[61][73] * vector[61] +matrix[62][73] * vector[62] +matrix[63][73] * vector[63] +matrix[64][73] * vector[64] +matrix[65][73] * vector[65] +matrix[66][73] * vector[66] +matrix[67][73] * vector[67] +matrix[68][73] * vector[68] +matrix[69][73] * vector[69] +matrix[70][73] * vector[70] +matrix[71][73] * vector[71] +matrix[72][73] * vector[72] +matrix[73][73] * vector[73] +matrix[74][73] * vector[74] +matrix[75][73] * vector[75] +matrix[76][73] * vector[76] +matrix[77][73] * vector[77] +matrix[78][73] * vector[78] +matrix[79][73] * vector[79] +matrix[80][73] * vector[80] +matrix[81][73] * vector[81] +matrix[82][73] * vector[82] +matrix[83][73] * vector[83] +matrix[84][73] * vector[84] +matrix[85][73] * vector[85] +matrix[86][73] * vector[86] +matrix[87][73] * vector[87] +matrix[88][73] * vector[88] +matrix[89][73] * vector[89] +matrix[90][73] * vector[90] +matrix[91][73] * vector[91] +matrix[92][73] * vector[92] +matrix[93][73] * vector[93] +matrix[94][73] * vector[94] +matrix[95][73] * vector[95] +matrix[96][73] * vector[96] +matrix[97][73] * vector[97] +matrix[98][73] * vector[98] +matrix[99][73] * vector[99] +b[73];
assign result[74] = matrix[0][74] * vector[0] +matrix[1][74] * vector[1] +matrix[2][74] * vector[2] +matrix[3][74] * vector[3] +matrix[4][74] * vector[4] +matrix[5][74] * vector[5] +matrix[6][74] * vector[6] +matrix[7][74] * vector[7] +matrix[8][74] * vector[8] +matrix[9][74] * vector[9] +matrix[10][74] * vector[10] +matrix[11][74] * vector[11] +matrix[12][74] * vector[12] +matrix[13][74] * vector[13] +matrix[14][74] * vector[14] +matrix[15][74] * vector[15] +matrix[16][74] * vector[16] +matrix[17][74] * vector[17] +matrix[18][74] * vector[18] +matrix[19][74] * vector[19] +matrix[20][74] * vector[20] +matrix[21][74] * vector[21] +matrix[22][74] * vector[22] +matrix[23][74] * vector[23] +matrix[24][74] * vector[24] +matrix[25][74] * vector[25] +matrix[26][74] * vector[26] +matrix[27][74] * vector[27] +matrix[28][74] * vector[28] +matrix[29][74] * vector[29] +matrix[30][74] * vector[30] +matrix[31][74] * vector[31] +matrix[32][74] * vector[32] +matrix[33][74] * vector[33] +matrix[34][74] * vector[34] +matrix[35][74] * vector[35] +matrix[36][74] * vector[36] +matrix[37][74] * vector[37] +matrix[38][74] * vector[38] +matrix[39][74] * vector[39] +matrix[40][74] * vector[40] +matrix[41][74] * vector[41] +matrix[42][74] * vector[42] +matrix[43][74] * vector[43] +matrix[44][74] * vector[44] +matrix[45][74] * vector[45] +matrix[46][74] * vector[46] +matrix[47][74] * vector[47] +matrix[48][74] * vector[48] +matrix[49][74] * vector[49] +matrix[50][74] * vector[50] +matrix[51][74] * vector[51] +matrix[52][74] * vector[52] +matrix[53][74] * vector[53] +matrix[54][74] * vector[54] +matrix[55][74] * vector[55] +matrix[56][74] * vector[56] +matrix[57][74] * vector[57] +matrix[58][74] * vector[58] +matrix[59][74] * vector[59] +matrix[60][74] * vector[60] +matrix[61][74] * vector[61] +matrix[62][74] * vector[62] +matrix[63][74] * vector[63] +matrix[64][74] * vector[64] +matrix[65][74] * vector[65] +matrix[66][74] * vector[66] +matrix[67][74] * vector[67] +matrix[68][74] * vector[68] +matrix[69][74] * vector[69] +matrix[70][74] * vector[70] +matrix[71][74] * vector[71] +matrix[72][74] * vector[72] +matrix[73][74] * vector[73] +matrix[74][74] * vector[74] +matrix[75][74] * vector[75] +matrix[76][74] * vector[76] +matrix[77][74] * vector[77] +matrix[78][74] * vector[78] +matrix[79][74] * vector[79] +matrix[80][74] * vector[80] +matrix[81][74] * vector[81] +matrix[82][74] * vector[82] +matrix[83][74] * vector[83] +matrix[84][74] * vector[84] +matrix[85][74] * vector[85] +matrix[86][74] * vector[86] +matrix[87][74] * vector[87] +matrix[88][74] * vector[88] +matrix[89][74] * vector[89] +matrix[90][74] * vector[90] +matrix[91][74] * vector[91] +matrix[92][74] * vector[92] +matrix[93][74] * vector[93] +matrix[94][74] * vector[94] +matrix[95][74] * vector[95] +matrix[96][74] * vector[96] +matrix[97][74] * vector[97] +matrix[98][74] * vector[98] +matrix[99][74] * vector[99] +b[74];
assign result[75] = matrix[0][75] * vector[0] +matrix[1][75] * vector[1] +matrix[2][75] * vector[2] +matrix[3][75] * vector[3] +matrix[4][75] * vector[4] +matrix[5][75] * vector[5] +matrix[6][75] * vector[6] +matrix[7][75] * vector[7] +matrix[8][75] * vector[8] +matrix[9][75] * vector[9] +matrix[10][75] * vector[10] +matrix[11][75] * vector[11] +matrix[12][75] * vector[12] +matrix[13][75] * vector[13] +matrix[14][75] * vector[14] +matrix[15][75] * vector[15] +matrix[16][75] * vector[16] +matrix[17][75] * vector[17] +matrix[18][75] * vector[18] +matrix[19][75] * vector[19] +matrix[20][75] * vector[20] +matrix[21][75] * vector[21] +matrix[22][75] * vector[22] +matrix[23][75] * vector[23] +matrix[24][75] * vector[24] +matrix[25][75] * vector[25] +matrix[26][75] * vector[26] +matrix[27][75] * vector[27] +matrix[28][75] * vector[28] +matrix[29][75] * vector[29] +matrix[30][75] * vector[30] +matrix[31][75] * vector[31] +matrix[32][75] * vector[32] +matrix[33][75] * vector[33] +matrix[34][75] * vector[34] +matrix[35][75] * vector[35] +matrix[36][75] * vector[36] +matrix[37][75] * vector[37] +matrix[38][75] * vector[38] +matrix[39][75] * vector[39] +matrix[40][75] * vector[40] +matrix[41][75] * vector[41] +matrix[42][75] * vector[42] +matrix[43][75] * vector[43] +matrix[44][75] * vector[44] +matrix[45][75] * vector[45] +matrix[46][75] * vector[46] +matrix[47][75] * vector[47] +matrix[48][75] * vector[48] +matrix[49][75] * vector[49] +matrix[50][75] * vector[50] +matrix[51][75] * vector[51] +matrix[52][75] * vector[52] +matrix[53][75] * vector[53] +matrix[54][75] * vector[54] +matrix[55][75] * vector[55] +matrix[56][75] * vector[56] +matrix[57][75] * vector[57] +matrix[58][75] * vector[58] +matrix[59][75] * vector[59] +matrix[60][75] * vector[60] +matrix[61][75] * vector[61] +matrix[62][75] * vector[62] +matrix[63][75] * vector[63] +matrix[64][75] * vector[64] +matrix[65][75] * vector[65] +matrix[66][75] * vector[66] +matrix[67][75] * vector[67] +matrix[68][75] * vector[68] +matrix[69][75] * vector[69] +matrix[70][75] * vector[70] +matrix[71][75] * vector[71] +matrix[72][75] * vector[72] +matrix[73][75] * vector[73] +matrix[74][75] * vector[74] +matrix[75][75] * vector[75] +matrix[76][75] * vector[76] +matrix[77][75] * vector[77] +matrix[78][75] * vector[78] +matrix[79][75] * vector[79] +matrix[80][75] * vector[80] +matrix[81][75] * vector[81] +matrix[82][75] * vector[82] +matrix[83][75] * vector[83] +matrix[84][75] * vector[84] +matrix[85][75] * vector[85] +matrix[86][75] * vector[86] +matrix[87][75] * vector[87] +matrix[88][75] * vector[88] +matrix[89][75] * vector[89] +matrix[90][75] * vector[90] +matrix[91][75] * vector[91] +matrix[92][75] * vector[92] +matrix[93][75] * vector[93] +matrix[94][75] * vector[94] +matrix[95][75] * vector[95] +matrix[96][75] * vector[96] +matrix[97][75] * vector[97] +matrix[98][75] * vector[98] +matrix[99][75] * vector[99] +b[75];
assign result[76] = matrix[0][76] * vector[0] +matrix[1][76] * vector[1] +matrix[2][76] * vector[2] +matrix[3][76] * vector[3] +matrix[4][76] * vector[4] +matrix[5][76] * vector[5] +matrix[6][76] * vector[6] +matrix[7][76] * vector[7] +matrix[8][76] * vector[8] +matrix[9][76] * vector[9] +matrix[10][76] * vector[10] +matrix[11][76] * vector[11] +matrix[12][76] * vector[12] +matrix[13][76] * vector[13] +matrix[14][76] * vector[14] +matrix[15][76] * vector[15] +matrix[16][76] * vector[16] +matrix[17][76] * vector[17] +matrix[18][76] * vector[18] +matrix[19][76] * vector[19] +matrix[20][76] * vector[20] +matrix[21][76] * vector[21] +matrix[22][76] * vector[22] +matrix[23][76] * vector[23] +matrix[24][76] * vector[24] +matrix[25][76] * vector[25] +matrix[26][76] * vector[26] +matrix[27][76] * vector[27] +matrix[28][76] * vector[28] +matrix[29][76] * vector[29] +matrix[30][76] * vector[30] +matrix[31][76] * vector[31] +matrix[32][76] * vector[32] +matrix[33][76] * vector[33] +matrix[34][76] * vector[34] +matrix[35][76] * vector[35] +matrix[36][76] * vector[36] +matrix[37][76] * vector[37] +matrix[38][76] * vector[38] +matrix[39][76] * vector[39] +matrix[40][76] * vector[40] +matrix[41][76] * vector[41] +matrix[42][76] * vector[42] +matrix[43][76] * vector[43] +matrix[44][76] * vector[44] +matrix[45][76] * vector[45] +matrix[46][76] * vector[46] +matrix[47][76] * vector[47] +matrix[48][76] * vector[48] +matrix[49][76] * vector[49] +matrix[50][76] * vector[50] +matrix[51][76] * vector[51] +matrix[52][76] * vector[52] +matrix[53][76] * vector[53] +matrix[54][76] * vector[54] +matrix[55][76] * vector[55] +matrix[56][76] * vector[56] +matrix[57][76] * vector[57] +matrix[58][76] * vector[58] +matrix[59][76] * vector[59] +matrix[60][76] * vector[60] +matrix[61][76] * vector[61] +matrix[62][76] * vector[62] +matrix[63][76] * vector[63] +matrix[64][76] * vector[64] +matrix[65][76] * vector[65] +matrix[66][76] * vector[66] +matrix[67][76] * vector[67] +matrix[68][76] * vector[68] +matrix[69][76] * vector[69] +matrix[70][76] * vector[70] +matrix[71][76] * vector[71] +matrix[72][76] * vector[72] +matrix[73][76] * vector[73] +matrix[74][76] * vector[74] +matrix[75][76] * vector[75] +matrix[76][76] * vector[76] +matrix[77][76] * vector[77] +matrix[78][76] * vector[78] +matrix[79][76] * vector[79] +matrix[80][76] * vector[80] +matrix[81][76] * vector[81] +matrix[82][76] * vector[82] +matrix[83][76] * vector[83] +matrix[84][76] * vector[84] +matrix[85][76] * vector[85] +matrix[86][76] * vector[86] +matrix[87][76] * vector[87] +matrix[88][76] * vector[88] +matrix[89][76] * vector[89] +matrix[90][76] * vector[90] +matrix[91][76] * vector[91] +matrix[92][76] * vector[92] +matrix[93][76] * vector[93] +matrix[94][76] * vector[94] +matrix[95][76] * vector[95] +matrix[96][76] * vector[96] +matrix[97][76] * vector[97] +matrix[98][76] * vector[98] +matrix[99][76] * vector[99] +b[76];
assign result[77] = matrix[0][77] * vector[0] +matrix[1][77] * vector[1] +matrix[2][77] * vector[2] +matrix[3][77] * vector[3] +matrix[4][77] * vector[4] +matrix[5][77] * vector[5] +matrix[6][77] * vector[6] +matrix[7][77] * vector[7] +matrix[8][77] * vector[8] +matrix[9][77] * vector[9] +matrix[10][77] * vector[10] +matrix[11][77] * vector[11] +matrix[12][77] * vector[12] +matrix[13][77] * vector[13] +matrix[14][77] * vector[14] +matrix[15][77] * vector[15] +matrix[16][77] * vector[16] +matrix[17][77] * vector[17] +matrix[18][77] * vector[18] +matrix[19][77] * vector[19] +matrix[20][77] * vector[20] +matrix[21][77] * vector[21] +matrix[22][77] * vector[22] +matrix[23][77] * vector[23] +matrix[24][77] * vector[24] +matrix[25][77] * vector[25] +matrix[26][77] * vector[26] +matrix[27][77] * vector[27] +matrix[28][77] * vector[28] +matrix[29][77] * vector[29] +matrix[30][77] * vector[30] +matrix[31][77] * vector[31] +matrix[32][77] * vector[32] +matrix[33][77] * vector[33] +matrix[34][77] * vector[34] +matrix[35][77] * vector[35] +matrix[36][77] * vector[36] +matrix[37][77] * vector[37] +matrix[38][77] * vector[38] +matrix[39][77] * vector[39] +matrix[40][77] * vector[40] +matrix[41][77] * vector[41] +matrix[42][77] * vector[42] +matrix[43][77] * vector[43] +matrix[44][77] * vector[44] +matrix[45][77] * vector[45] +matrix[46][77] * vector[46] +matrix[47][77] * vector[47] +matrix[48][77] * vector[48] +matrix[49][77] * vector[49] +matrix[50][77] * vector[50] +matrix[51][77] * vector[51] +matrix[52][77] * vector[52] +matrix[53][77] * vector[53] +matrix[54][77] * vector[54] +matrix[55][77] * vector[55] +matrix[56][77] * vector[56] +matrix[57][77] * vector[57] +matrix[58][77] * vector[58] +matrix[59][77] * vector[59] +matrix[60][77] * vector[60] +matrix[61][77] * vector[61] +matrix[62][77] * vector[62] +matrix[63][77] * vector[63] +matrix[64][77] * vector[64] +matrix[65][77] * vector[65] +matrix[66][77] * vector[66] +matrix[67][77] * vector[67] +matrix[68][77] * vector[68] +matrix[69][77] * vector[69] +matrix[70][77] * vector[70] +matrix[71][77] * vector[71] +matrix[72][77] * vector[72] +matrix[73][77] * vector[73] +matrix[74][77] * vector[74] +matrix[75][77] * vector[75] +matrix[76][77] * vector[76] +matrix[77][77] * vector[77] +matrix[78][77] * vector[78] +matrix[79][77] * vector[79] +matrix[80][77] * vector[80] +matrix[81][77] * vector[81] +matrix[82][77] * vector[82] +matrix[83][77] * vector[83] +matrix[84][77] * vector[84] +matrix[85][77] * vector[85] +matrix[86][77] * vector[86] +matrix[87][77] * vector[87] +matrix[88][77] * vector[88] +matrix[89][77] * vector[89] +matrix[90][77] * vector[90] +matrix[91][77] * vector[91] +matrix[92][77] * vector[92] +matrix[93][77] * vector[93] +matrix[94][77] * vector[94] +matrix[95][77] * vector[95] +matrix[96][77] * vector[96] +matrix[97][77] * vector[97] +matrix[98][77] * vector[98] +matrix[99][77] * vector[99] +b[77];
assign result[78] = matrix[0][78] * vector[0] +matrix[1][78] * vector[1] +matrix[2][78] * vector[2] +matrix[3][78] * vector[3] +matrix[4][78] * vector[4] +matrix[5][78] * vector[5] +matrix[6][78] * vector[6] +matrix[7][78] * vector[7] +matrix[8][78] * vector[8] +matrix[9][78] * vector[9] +matrix[10][78] * vector[10] +matrix[11][78] * vector[11] +matrix[12][78] * vector[12] +matrix[13][78] * vector[13] +matrix[14][78] * vector[14] +matrix[15][78] * vector[15] +matrix[16][78] * vector[16] +matrix[17][78] * vector[17] +matrix[18][78] * vector[18] +matrix[19][78] * vector[19] +matrix[20][78] * vector[20] +matrix[21][78] * vector[21] +matrix[22][78] * vector[22] +matrix[23][78] * vector[23] +matrix[24][78] * vector[24] +matrix[25][78] * vector[25] +matrix[26][78] * vector[26] +matrix[27][78] * vector[27] +matrix[28][78] * vector[28] +matrix[29][78] * vector[29] +matrix[30][78] * vector[30] +matrix[31][78] * vector[31] +matrix[32][78] * vector[32] +matrix[33][78] * vector[33] +matrix[34][78] * vector[34] +matrix[35][78] * vector[35] +matrix[36][78] * vector[36] +matrix[37][78] * vector[37] +matrix[38][78] * vector[38] +matrix[39][78] * vector[39] +matrix[40][78] * vector[40] +matrix[41][78] * vector[41] +matrix[42][78] * vector[42] +matrix[43][78] * vector[43] +matrix[44][78] * vector[44] +matrix[45][78] * vector[45] +matrix[46][78] * vector[46] +matrix[47][78] * vector[47] +matrix[48][78] * vector[48] +matrix[49][78] * vector[49] +matrix[50][78] * vector[50] +matrix[51][78] * vector[51] +matrix[52][78] * vector[52] +matrix[53][78] * vector[53] +matrix[54][78] * vector[54] +matrix[55][78] * vector[55] +matrix[56][78] * vector[56] +matrix[57][78] * vector[57] +matrix[58][78] * vector[58] +matrix[59][78] * vector[59] +matrix[60][78] * vector[60] +matrix[61][78] * vector[61] +matrix[62][78] * vector[62] +matrix[63][78] * vector[63] +matrix[64][78] * vector[64] +matrix[65][78] * vector[65] +matrix[66][78] * vector[66] +matrix[67][78] * vector[67] +matrix[68][78] * vector[68] +matrix[69][78] * vector[69] +matrix[70][78] * vector[70] +matrix[71][78] * vector[71] +matrix[72][78] * vector[72] +matrix[73][78] * vector[73] +matrix[74][78] * vector[74] +matrix[75][78] * vector[75] +matrix[76][78] * vector[76] +matrix[77][78] * vector[77] +matrix[78][78] * vector[78] +matrix[79][78] * vector[79] +matrix[80][78] * vector[80] +matrix[81][78] * vector[81] +matrix[82][78] * vector[82] +matrix[83][78] * vector[83] +matrix[84][78] * vector[84] +matrix[85][78] * vector[85] +matrix[86][78] * vector[86] +matrix[87][78] * vector[87] +matrix[88][78] * vector[88] +matrix[89][78] * vector[89] +matrix[90][78] * vector[90] +matrix[91][78] * vector[91] +matrix[92][78] * vector[92] +matrix[93][78] * vector[93] +matrix[94][78] * vector[94] +matrix[95][78] * vector[95] +matrix[96][78] * vector[96] +matrix[97][78] * vector[97] +matrix[98][78] * vector[98] +matrix[99][78] * vector[99] +b[78];
assign result[79] = matrix[0][79] * vector[0] +matrix[1][79] * vector[1] +matrix[2][79] * vector[2] +matrix[3][79] * vector[3] +matrix[4][79] * vector[4] +matrix[5][79] * vector[5] +matrix[6][79] * vector[6] +matrix[7][79] * vector[7] +matrix[8][79] * vector[8] +matrix[9][79] * vector[9] +matrix[10][79] * vector[10] +matrix[11][79] * vector[11] +matrix[12][79] * vector[12] +matrix[13][79] * vector[13] +matrix[14][79] * vector[14] +matrix[15][79] * vector[15] +matrix[16][79] * vector[16] +matrix[17][79] * vector[17] +matrix[18][79] * vector[18] +matrix[19][79] * vector[19] +matrix[20][79] * vector[20] +matrix[21][79] * vector[21] +matrix[22][79] * vector[22] +matrix[23][79] * vector[23] +matrix[24][79] * vector[24] +matrix[25][79] * vector[25] +matrix[26][79] * vector[26] +matrix[27][79] * vector[27] +matrix[28][79] * vector[28] +matrix[29][79] * vector[29] +matrix[30][79] * vector[30] +matrix[31][79] * vector[31] +matrix[32][79] * vector[32] +matrix[33][79] * vector[33] +matrix[34][79] * vector[34] +matrix[35][79] * vector[35] +matrix[36][79] * vector[36] +matrix[37][79] * vector[37] +matrix[38][79] * vector[38] +matrix[39][79] * vector[39] +matrix[40][79] * vector[40] +matrix[41][79] * vector[41] +matrix[42][79] * vector[42] +matrix[43][79] * vector[43] +matrix[44][79] * vector[44] +matrix[45][79] * vector[45] +matrix[46][79] * vector[46] +matrix[47][79] * vector[47] +matrix[48][79] * vector[48] +matrix[49][79] * vector[49] +matrix[50][79] * vector[50] +matrix[51][79] * vector[51] +matrix[52][79] * vector[52] +matrix[53][79] * vector[53] +matrix[54][79] * vector[54] +matrix[55][79] * vector[55] +matrix[56][79] * vector[56] +matrix[57][79] * vector[57] +matrix[58][79] * vector[58] +matrix[59][79] * vector[59] +matrix[60][79] * vector[60] +matrix[61][79] * vector[61] +matrix[62][79] * vector[62] +matrix[63][79] * vector[63] +matrix[64][79] * vector[64] +matrix[65][79] * vector[65] +matrix[66][79] * vector[66] +matrix[67][79] * vector[67] +matrix[68][79] * vector[68] +matrix[69][79] * vector[69] +matrix[70][79] * vector[70] +matrix[71][79] * vector[71] +matrix[72][79] * vector[72] +matrix[73][79] * vector[73] +matrix[74][79] * vector[74] +matrix[75][79] * vector[75] +matrix[76][79] * vector[76] +matrix[77][79] * vector[77] +matrix[78][79] * vector[78] +matrix[79][79] * vector[79] +matrix[80][79] * vector[80] +matrix[81][79] * vector[81] +matrix[82][79] * vector[82] +matrix[83][79] * vector[83] +matrix[84][79] * vector[84] +matrix[85][79] * vector[85] +matrix[86][79] * vector[86] +matrix[87][79] * vector[87] +matrix[88][79] * vector[88] +matrix[89][79] * vector[89] +matrix[90][79] * vector[90] +matrix[91][79] * vector[91] +matrix[92][79] * vector[92] +matrix[93][79] * vector[93] +matrix[94][79] * vector[94] +matrix[95][79] * vector[95] +matrix[96][79] * vector[96] +matrix[97][79] * vector[97] +matrix[98][79] * vector[98] +matrix[99][79] * vector[99] +b[79];
assign result[80] = matrix[0][80] * vector[0] +matrix[1][80] * vector[1] +matrix[2][80] * vector[2] +matrix[3][80] * vector[3] +matrix[4][80] * vector[4] +matrix[5][80] * vector[5] +matrix[6][80] * vector[6] +matrix[7][80] * vector[7] +matrix[8][80] * vector[8] +matrix[9][80] * vector[9] +matrix[10][80] * vector[10] +matrix[11][80] * vector[11] +matrix[12][80] * vector[12] +matrix[13][80] * vector[13] +matrix[14][80] * vector[14] +matrix[15][80] * vector[15] +matrix[16][80] * vector[16] +matrix[17][80] * vector[17] +matrix[18][80] * vector[18] +matrix[19][80] * vector[19] +matrix[20][80] * vector[20] +matrix[21][80] * vector[21] +matrix[22][80] * vector[22] +matrix[23][80] * vector[23] +matrix[24][80] * vector[24] +matrix[25][80] * vector[25] +matrix[26][80] * vector[26] +matrix[27][80] * vector[27] +matrix[28][80] * vector[28] +matrix[29][80] * vector[29] +matrix[30][80] * vector[30] +matrix[31][80] * vector[31] +matrix[32][80] * vector[32] +matrix[33][80] * vector[33] +matrix[34][80] * vector[34] +matrix[35][80] * vector[35] +matrix[36][80] * vector[36] +matrix[37][80] * vector[37] +matrix[38][80] * vector[38] +matrix[39][80] * vector[39] +matrix[40][80] * vector[40] +matrix[41][80] * vector[41] +matrix[42][80] * vector[42] +matrix[43][80] * vector[43] +matrix[44][80] * vector[44] +matrix[45][80] * vector[45] +matrix[46][80] * vector[46] +matrix[47][80] * vector[47] +matrix[48][80] * vector[48] +matrix[49][80] * vector[49] +matrix[50][80] * vector[50] +matrix[51][80] * vector[51] +matrix[52][80] * vector[52] +matrix[53][80] * vector[53] +matrix[54][80] * vector[54] +matrix[55][80] * vector[55] +matrix[56][80] * vector[56] +matrix[57][80] * vector[57] +matrix[58][80] * vector[58] +matrix[59][80] * vector[59] +matrix[60][80] * vector[60] +matrix[61][80] * vector[61] +matrix[62][80] * vector[62] +matrix[63][80] * vector[63] +matrix[64][80] * vector[64] +matrix[65][80] * vector[65] +matrix[66][80] * vector[66] +matrix[67][80] * vector[67] +matrix[68][80] * vector[68] +matrix[69][80] * vector[69] +matrix[70][80] * vector[70] +matrix[71][80] * vector[71] +matrix[72][80] * vector[72] +matrix[73][80] * vector[73] +matrix[74][80] * vector[74] +matrix[75][80] * vector[75] +matrix[76][80] * vector[76] +matrix[77][80] * vector[77] +matrix[78][80] * vector[78] +matrix[79][80] * vector[79] +matrix[80][80] * vector[80] +matrix[81][80] * vector[81] +matrix[82][80] * vector[82] +matrix[83][80] * vector[83] +matrix[84][80] * vector[84] +matrix[85][80] * vector[85] +matrix[86][80] * vector[86] +matrix[87][80] * vector[87] +matrix[88][80] * vector[88] +matrix[89][80] * vector[89] +matrix[90][80] * vector[90] +matrix[91][80] * vector[91] +matrix[92][80] * vector[92] +matrix[93][80] * vector[93] +matrix[94][80] * vector[94] +matrix[95][80] * vector[95] +matrix[96][80] * vector[96] +matrix[97][80] * vector[97] +matrix[98][80] * vector[98] +matrix[99][80] * vector[99] +b[80];
assign result[81] = matrix[0][81] * vector[0] +matrix[1][81] * vector[1] +matrix[2][81] * vector[2] +matrix[3][81] * vector[3] +matrix[4][81] * vector[4] +matrix[5][81] * vector[5] +matrix[6][81] * vector[6] +matrix[7][81] * vector[7] +matrix[8][81] * vector[8] +matrix[9][81] * vector[9] +matrix[10][81] * vector[10] +matrix[11][81] * vector[11] +matrix[12][81] * vector[12] +matrix[13][81] * vector[13] +matrix[14][81] * vector[14] +matrix[15][81] * vector[15] +matrix[16][81] * vector[16] +matrix[17][81] * vector[17] +matrix[18][81] * vector[18] +matrix[19][81] * vector[19] +matrix[20][81] * vector[20] +matrix[21][81] * vector[21] +matrix[22][81] * vector[22] +matrix[23][81] * vector[23] +matrix[24][81] * vector[24] +matrix[25][81] * vector[25] +matrix[26][81] * vector[26] +matrix[27][81] * vector[27] +matrix[28][81] * vector[28] +matrix[29][81] * vector[29] +matrix[30][81] * vector[30] +matrix[31][81] * vector[31] +matrix[32][81] * vector[32] +matrix[33][81] * vector[33] +matrix[34][81] * vector[34] +matrix[35][81] * vector[35] +matrix[36][81] * vector[36] +matrix[37][81] * vector[37] +matrix[38][81] * vector[38] +matrix[39][81] * vector[39] +matrix[40][81] * vector[40] +matrix[41][81] * vector[41] +matrix[42][81] * vector[42] +matrix[43][81] * vector[43] +matrix[44][81] * vector[44] +matrix[45][81] * vector[45] +matrix[46][81] * vector[46] +matrix[47][81] * vector[47] +matrix[48][81] * vector[48] +matrix[49][81] * vector[49] +matrix[50][81] * vector[50] +matrix[51][81] * vector[51] +matrix[52][81] * vector[52] +matrix[53][81] * vector[53] +matrix[54][81] * vector[54] +matrix[55][81] * vector[55] +matrix[56][81] * vector[56] +matrix[57][81] * vector[57] +matrix[58][81] * vector[58] +matrix[59][81] * vector[59] +matrix[60][81] * vector[60] +matrix[61][81] * vector[61] +matrix[62][81] * vector[62] +matrix[63][81] * vector[63] +matrix[64][81] * vector[64] +matrix[65][81] * vector[65] +matrix[66][81] * vector[66] +matrix[67][81] * vector[67] +matrix[68][81] * vector[68] +matrix[69][81] * vector[69] +matrix[70][81] * vector[70] +matrix[71][81] * vector[71] +matrix[72][81] * vector[72] +matrix[73][81] * vector[73] +matrix[74][81] * vector[74] +matrix[75][81] * vector[75] +matrix[76][81] * vector[76] +matrix[77][81] * vector[77] +matrix[78][81] * vector[78] +matrix[79][81] * vector[79] +matrix[80][81] * vector[80] +matrix[81][81] * vector[81] +matrix[82][81] * vector[82] +matrix[83][81] * vector[83] +matrix[84][81] * vector[84] +matrix[85][81] * vector[85] +matrix[86][81] * vector[86] +matrix[87][81] * vector[87] +matrix[88][81] * vector[88] +matrix[89][81] * vector[89] +matrix[90][81] * vector[90] +matrix[91][81] * vector[91] +matrix[92][81] * vector[92] +matrix[93][81] * vector[93] +matrix[94][81] * vector[94] +matrix[95][81] * vector[95] +matrix[96][81] * vector[96] +matrix[97][81] * vector[97] +matrix[98][81] * vector[98] +matrix[99][81] * vector[99] +b[81];
assign result[82] = matrix[0][82] * vector[0] +matrix[1][82] * vector[1] +matrix[2][82] * vector[2] +matrix[3][82] * vector[3] +matrix[4][82] * vector[4] +matrix[5][82] * vector[5] +matrix[6][82] * vector[6] +matrix[7][82] * vector[7] +matrix[8][82] * vector[8] +matrix[9][82] * vector[9] +matrix[10][82] * vector[10] +matrix[11][82] * vector[11] +matrix[12][82] * vector[12] +matrix[13][82] * vector[13] +matrix[14][82] * vector[14] +matrix[15][82] * vector[15] +matrix[16][82] * vector[16] +matrix[17][82] * vector[17] +matrix[18][82] * vector[18] +matrix[19][82] * vector[19] +matrix[20][82] * vector[20] +matrix[21][82] * vector[21] +matrix[22][82] * vector[22] +matrix[23][82] * vector[23] +matrix[24][82] * vector[24] +matrix[25][82] * vector[25] +matrix[26][82] * vector[26] +matrix[27][82] * vector[27] +matrix[28][82] * vector[28] +matrix[29][82] * vector[29] +matrix[30][82] * vector[30] +matrix[31][82] * vector[31] +matrix[32][82] * vector[32] +matrix[33][82] * vector[33] +matrix[34][82] * vector[34] +matrix[35][82] * vector[35] +matrix[36][82] * vector[36] +matrix[37][82] * vector[37] +matrix[38][82] * vector[38] +matrix[39][82] * vector[39] +matrix[40][82] * vector[40] +matrix[41][82] * vector[41] +matrix[42][82] * vector[42] +matrix[43][82] * vector[43] +matrix[44][82] * vector[44] +matrix[45][82] * vector[45] +matrix[46][82] * vector[46] +matrix[47][82] * vector[47] +matrix[48][82] * vector[48] +matrix[49][82] * vector[49] +matrix[50][82] * vector[50] +matrix[51][82] * vector[51] +matrix[52][82] * vector[52] +matrix[53][82] * vector[53] +matrix[54][82] * vector[54] +matrix[55][82] * vector[55] +matrix[56][82] * vector[56] +matrix[57][82] * vector[57] +matrix[58][82] * vector[58] +matrix[59][82] * vector[59] +matrix[60][82] * vector[60] +matrix[61][82] * vector[61] +matrix[62][82] * vector[62] +matrix[63][82] * vector[63] +matrix[64][82] * vector[64] +matrix[65][82] * vector[65] +matrix[66][82] * vector[66] +matrix[67][82] * vector[67] +matrix[68][82] * vector[68] +matrix[69][82] * vector[69] +matrix[70][82] * vector[70] +matrix[71][82] * vector[71] +matrix[72][82] * vector[72] +matrix[73][82] * vector[73] +matrix[74][82] * vector[74] +matrix[75][82] * vector[75] +matrix[76][82] * vector[76] +matrix[77][82] * vector[77] +matrix[78][82] * vector[78] +matrix[79][82] * vector[79] +matrix[80][82] * vector[80] +matrix[81][82] * vector[81] +matrix[82][82] * vector[82] +matrix[83][82] * vector[83] +matrix[84][82] * vector[84] +matrix[85][82] * vector[85] +matrix[86][82] * vector[86] +matrix[87][82] * vector[87] +matrix[88][82] * vector[88] +matrix[89][82] * vector[89] +matrix[90][82] * vector[90] +matrix[91][82] * vector[91] +matrix[92][82] * vector[92] +matrix[93][82] * vector[93] +matrix[94][82] * vector[94] +matrix[95][82] * vector[95] +matrix[96][82] * vector[96] +matrix[97][82] * vector[97] +matrix[98][82] * vector[98] +matrix[99][82] * vector[99] +b[82];
assign result[83] = matrix[0][83] * vector[0] +matrix[1][83] * vector[1] +matrix[2][83] * vector[2] +matrix[3][83] * vector[3] +matrix[4][83] * vector[4] +matrix[5][83] * vector[5] +matrix[6][83] * vector[6] +matrix[7][83] * vector[7] +matrix[8][83] * vector[8] +matrix[9][83] * vector[9] +matrix[10][83] * vector[10] +matrix[11][83] * vector[11] +matrix[12][83] * vector[12] +matrix[13][83] * vector[13] +matrix[14][83] * vector[14] +matrix[15][83] * vector[15] +matrix[16][83] * vector[16] +matrix[17][83] * vector[17] +matrix[18][83] * vector[18] +matrix[19][83] * vector[19] +matrix[20][83] * vector[20] +matrix[21][83] * vector[21] +matrix[22][83] * vector[22] +matrix[23][83] * vector[23] +matrix[24][83] * vector[24] +matrix[25][83] * vector[25] +matrix[26][83] * vector[26] +matrix[27][83] * vector[27] +matrix[28][83] * vector[28] +matrix[29][83] * vector[29] +matrix[30][83] * vector[30] +matrix[31][83] * vector[31] +matrix[32][83] * vector[32] +matrix[33][83] * vector[33] +matrix[34][83] * vector[34] +matrix[35][83] * vector[35] +matrix[36][83] * vector[36] +matrix[37][83] * vector[37] +matrix[38][83] * vector[38] +matrix[39][83] * vector[39] +matrix[40][83] * vector[40] +matrix[41][83] * vector[41] +matrix[42][83] * vector[42] +matrix[43][83] * vector[43] +matrix[44][83] * vector[44] +matrix[45][83] * vector[45] +matrix[46][83] * vector[46] +matrix[47][83] * vector[47] +matrix[48][83] * vector[48] +matrix[49][83] * vector[49] +matrix[50][83] * vector[50] +matrix[51][83] * vector[51] +matrix[52][83] * vector[52] +matrix[53][83] * vector[53] +matrix[54][83] * vector[54] +matrix[55][83] * vector[55] +matrix[56][83] * vector[56] +matrix[57][83] * vector[57] +matrix[58][83] * vector[58] +matrix[59][83] * vector[59] +matrix[60][83] * vector[60] +matrix[61][83] * vector[61] +matrix[62][83] * vector[62] +matrix[63][83] * vector[63] +matrix[64][83] * vector[64] +matrix[65][83] * vector[65] +matrix[66][83] * vector[66] +matrix[67][83] * vector[67] +matrix[68][83] * vector[68] +matrix[69][83] * vector[69] +matrix[70][83] * vector[70] +matrix[71][83] * vector[71] +matrix[72][83] * vector[72] +matrix[73][83] * vector[73] +matrix[74][83] * vector[74] +matrix[75][83] * vector[75] +matrix[76][83] * vector[76] +matrix[77][83] * vector[77] +matrix[78][83] * vector[78] +matrix[79][83] * vector[79] +matrix[80][83] * vector[80] +matrix[81][83] * vector[81] +matrix[82][83] * vector[82] +matrix[83][83] * vector[83] +matrix[84][83] * vector[84] +matrix[85][83] * vector[85] +matrix[86][83] * vector[86] +matrix[87][83] * vector[87] +matrix[88][83] * vector[88] +matrix[89][83] * vector[89] +matrix[90][83] * vector[90] +matrix[91][83] * vector[91] +matrix[92][83] * vector[92] +matrix[93][83] * vector[93] +matrix[94][83] * vector[94] +matrix[95][83] * vector[95] +matrix[96][83] * vector[96] +matrix[97][83] * vector[97] +matrix[98][83] * vector[98] +matrix[99][83] * vector[99] +b[83];
assign result[84] = matrix[0][84] * vector[0] +matrix[1][84] * vector[1] +matrix[2][84] * vector[2] +matrix[3][84] * vector[3] +matrix[4][84] * vector[4] +matrix[5][84] * vector[5] +matrix[6][84] * vector[6] +matrix[7][84] * vector[7] +matrix[8][84] * vector[8] +matrix[9][84] * vector[9] +matrix[10][84] * vector[10] +matrix[11][84] * vector[11] +matrix[12][84] * vector[12] +matrix[13][84] * vector[13] +matrix[14][84] * vector[14] +matrix[15][84] * vector[15] +matrix[16][84] * vector[16] +matrix[17][84] * vector[17] +matrix[18][84] * vector[18] +matrix[19][84] * vector[19] +matrix[20][84] * vector[20] +matrix[21][84] * vector[21] +matrix[22][84] * vector[22] +matrix[23][84] * vector[23] +matrix[24][84] * vector[24] +matrix[25][84] * vector[25] +matrix[26][84] * vector[26] +matrix[27][84] * vector[27] +matrix[28][84] * vector[28] +matrix[29][84] * vector[29] +matrix[30][84] * vector[30] +matrix[31][84] * vector[31] +matrix[32][84] * vector[32] +matrix[33][84] * vector[33] +matrix[34][84] * vector[34] +matrix[35][84] * vector[35] +matrix[36][84] * vector[36] +matrix[37][84] * vector[37] +matrix[38][84] * vector[38] +matrix[39][84] * vector[39] +matrix[40][84] * vector[40] +matrix[41][84] * vector[41] +matrix[42][84] * vector[42] +matrix[43][84] * vector[43] +matrix[44][84] * vector[44] +matrix[45][84] * vector[45] +matrix[46][84] * vector[46] +matrix[47][84] * vector[47] +matrix[48][84] * vector[48] +matrix[49][84] * vector[49] +matrix[50][84] * vector[50] +matrix[51][84] * vector[51] +matrix[52][84] * vector[52] +matrix[53][84] * vector[53] +matrix[54][84] * vector[54] +matrix[55][84] * vector[55] +matrix[56][84] * vector[56] +matrix[57][84] * vector[57] +matrix[58][84] * vector[58] +matrix[59][84] * vector[59] +matrix[60][84] * vector[60] +matrix[61][84] * vector[61] +matrix[62][84] * vector[62] +matrix[63][84] * vector[63] +matrix[64][84] * vector[64] +matrix[65][84] * vector[65] +matrix[66][84] * vector[66] +matrix[67][84] * vector[67] +matrix[68][84] * vector[68] +matrix[69][84] * vector[69] +matrix[70][84] * vector[70] +matrix[71][84] * vector[71] +matrix[72][84] * vector[72] +matrix[73][84] * vector[73] +matrix[74][84] * vector[74] +matrix[75][84] * vector[75] +matrix[76][84] * vector[76] +matrix[77][84] * vector[77] +matrix[78][84] * vector[78] +matrix[79][84] * vector[79] +matrix[80][84] * vector[80] +matrix[81][84] * vector[81] +matrix[82][84] * vector[82] +matrix[83][84] * vector[83] +matrix[84][84] * vector[84] +matrix[85][84] * vector[85] +matrix[86][84] * vector[86] +matrix[87][84] * vector[87] +matrix[88][84] * vector[88] +matrix[89][84] * vector[89] +matrix[90][84] * vector[90] +matrix[91][84] * vector[91] +matrix[92][84] * vector[92] +matrix[93][84] * vector[93] +matrix[94][84] * vector[94] +matrix[95][84] * vector[95] +matrix[96][84] * vector[96] +matrix[97][84] * vector[97] +matrix[98][84] * vector[98] +matrix[99][84] * vector[99] +b[84];
assign result[85] = matrix[0][85] * vector[0] +matrix[1][85] * vector[1] +matrix[2][85] * vector[2] +matrix[3][85] * vector[3] +matrix[4][85] * vector[4] +matrix[5][85] * vector[5] +matrix[6][85] * vector[6] +matrix[7][85] * vector[7] +matrix[8][85] * vector[8] +matrix[9][85] * vector[9] +matrix[10][85] * vector[10] +matrix[11][85] * vector[11] +matrix[12][85] * vector[12] +matrix[13][85] * vector[13] +matrix[14][85] * vector[14] +matrix[15][85] * vector[15] +matrix[16][85] * vector[16] +matrix[17][85] * vector[17] +matrix[18][85] * vector[18] +matrix[19][85] * vector[19] +matrix[20][85] * vector[20] +matrix[21][85] * vector[21] +matrix[22][85] * vector[22] +matrix[23][85] * vector[23] +matrix[24][85] * vector[24] +matrix[25][85] * vector[25] +matrix[26][85] * vector[26] +matrix[27][85] * vector[27] +matrix[28][85] * vector[28] +matrix[29][85] * vector[29] +matrix[30][85] * vector[30] +matrix[31][85] * vector[31] +matrix[32][85] * vector[32] +matrix[33][85] * vector[33] +matrix[34][85] * vector[34] +matrix[35][85] * vector[35] +matrix[36][85] * vector[36] +matrix[37][85] * vector[37] +matrix[38][85] * vector[38] +matrix[39][85] * vector[39] +matrix[40][85] * vector[40] +matrix[41][85] * vector[41] +matrix[42][85] * vector[42] +matrix[43][85] * vector[43] +matrix[44][85] * vector[44] +matrix[45][85] * vector[45] +matrix[46][85] * vector[46] +matrix[47][85] * vector[47] +matrix[48][85] * vector[48] +matrix[49][85] * vector[49] +matrix[50][85] * vector[50] +matrix[51][85] * vector[51] +matrix[52][85] * vector[52] +matrix[53][85] * vector[53] +matrix[54][85] * vector[54] +matrix[55][85] * vector[55] +matrix[56][85] * vector[56] +matrix[57][85] * vector[57] +matrix[58][85] * vector[58] +matrix[59][85] * vector[59] +matrix[60][85] * vector[60] +matrix[61][85] * vector[61] +matrix[62][85] * vector[62] +matrix[63][85] * vector[63] +matrix[64][85] * vector[64] +matrix[65][85] * vector[65] +matrix[66][85] * vector[66] +matrix[67][85] * vector[67] +matrix[68][85] * vector[68] +matrix[69][85] * vector[69] +matrix[70][85] * vector[70] +matrix[71][85] * vector[71] +matrix[72][85] * vector[72] +matrix[73][85] * vector[73] +matrix[74][85] * vector[74] +matrix[75][85] * vector[75] +matrix[76][85] * vector[76] +matrix[77][85] * vector[77] +matrix[78][85] * vector[78] +matrix[79][85] * vector[79] +matrix[80][85] * vector[80] +matrix[81][85] * vector[81] +matrix[82][85] * vector[82] +matrix[83][85] * vector[83] +matrix[84][85] * vector[84] +matrix[85][85] * vector[85] +matrix[86][85] * vector[86] +matrix[87][85] * vector[87] +matrix[88][85] * vector[88] +matrix[89][85] * vector[89] +matrix[90][85] * vector[90] +matrix[91][85] * vector[91] +matrix[92][85] * vector[92] +matrix[93][85] * vector[93] +matrix[94][85] * vector[94] +matrix[95][85] * vector[95] +matrix[96][85] * vector[96] +matrix[97][85] * vector[97] +matrix[98][85] * vector[98] +matrix[99][85] * vector[99] +b[85];
assign result[86] = matrix[0][86] * vector[0] +matrix[1][86] * vector[1] +matrix[2][86] * vector[2] +matrix[3][86] * vector[3] +matrix[4][86] * vector[4] +matrix[5][86] * vector[5] +matrix[6][86] * vector[6] +matrix[7][86] * vector[7] +matrix[8][86] * vector[8] +matrix[9][86] * vector[9] +matrix[10][86] * vector[10] +matrix[11][86] * vector[11] +matrix[12][86] * vector[12] +matrix[13][86] * vector[13] +matrix[14][86] * vector[14] +matrix[15][86] * vector[15] +matrix[16][86] * vector[16] +matrix[17][86] * vector[17] +matrix[18][86] * vector[18] +matrix[19][86] * vector[19] +matrix[20][86] * vector[20] +matrix[21][86] * vector[21] +matrix[22][86] * vector[22] +matrix[23][86] * vector[23] +matrix[24][86] * vector[24] +matrix[25][86] * vector[25] +matrix[26][86] * vector[26] +matrix[27][86] * vector[27] +matrix[28][86] * vector[28] +matrix[29][86] * vector[29] +matrix[30][86] * vector[30] +matrix[31][86] * vector[31] +matrix[32][86] * vector[32] +matrix[33][86] * vector[33] +matrix[34][86] * vector[34] +matrix[35][86] * vector[35] +matrix[36][86] * vector[36] +matrix[37][86] * vector[37] +matrix[38][86] * vector[38] +matrix[39][86] * vector[39] +matrix[40][86] * vector[40] +matrix[41][86] * vector[41] +matrix[42][86] * vector[42] +matrix[43][86] * vector[43] +matrix[44][86] * vector[44] +matrix[45][86] * vector[45] +matrix[46][86] * vector[46] +matrix[47][86] * vector[47] +matrix[48][86] * vector[48] +matrix[49][86] * vector[49] +matrix[50][86] * vector[50] +matrix[51][86] * vector[51] +matrix[52][86] * vector[52] +matrix[53][86] * vector[53] +matrix[54][86] * vector[54] +matrix[55][86] * vector[55] +matrix[56][86] * vector[56] +matrix[57][86] * vector[57] +matrix[58][86] * vector[58] +matrix[59][86] * vector[59] +matrix[60][86] * vector[60] +matrix[61][86] * vector[61] +matrix[62][86] * vector[62] +matrix[63][86] * vector[63] +matrix[64][86] * vector[64] +matrix[65][86] * vector[65] +matrix[66][86] * vector[66] +matrix[67][86] * vector[67] +matrix[68][86] * vector[68] +matrix[69][86] * vector[69] +matrix[70][86] * vector[70] +matrix[71][86] * vector[71] +matrix[72][86] * vector[72] +matrix[73][86] * vector[73] +matrix[74][86] * vector[74] +matrix[75][86] * vector[75] +matrix[76][86] * vector[76] +matrix[77][86] * vector[77] +matrix[78][86] * vector[78] +matrix[79][86] * vector[79] +matrix[80][86] * vector[80] +matrix[81][86] * vector[81] +matrix[82][86] * vector[82] +matrix[83][86] * vector[83] +matrix[84][86] * vector[84] +matrix[85][86] * vector[85] +matrix[86][86] * vector[86] +matrix[87][86] * vector[87] +matrix[88][86] * vector[88] +matrix[89][86] * vector[89] +matrix[90][86] * vector[90] +matrix[91][86] * vector[91] +matrix[92][86] * vector[92] +matrix[93][86] * vector[93] +matrix[94][86] * vector[94] +matrix[95][86] * vector[95] +matrix[96][86] * vector[96] +matrix[97][86] * vector[97] +matrix[98][86] * vector[98] +matrix[99][86] * vector[99] +b[86];
assign result[87] = matrix[0][87] * vector[0] +matrix[1][87] * vector[1] +matrix[2][87] * vector[2] +matrix[3][87] * vector[3] +matrix[4][87] * vector[4] +matrix[5][87] * vector[5] +matrix[6][87] * vector[6] +matrix[7][87] * vector[7] +matrix[8][87] * vector[8] +matrix[9][87] * vector[9] +matrix[10][87] * vector[10] +matrix[11][87] * vector[11] +matrix[12][87] * vector[12] +matrix[13][87] * vector[13] +matrix[14][87] * vector[14] +matrix[15][87] * vector[15] +matrix[16][87] * vector[16] +matrix[17][87] * vector[17] +matrix[18][87] * vector[18] +matrix[19][87] * vector[19] +matrix[20][87] * vector[20] +matrix[21][87] * vector[21] +matrix[22][87] * vector[22] +matrix[23][87] * vector[23] +matrix[24][87] * vector[24] +matrix[25][87] * vector[25] +matrix[26][87] * vector[26] +matrix[27][87] * vector[27] +matrix[28][87] * vector[28] +matrix[29][87] * vector[29] +matrix[30][87] * vector[30] +matrix[31][87] * vector[31] +matrix[32][87] * vector[32] +matrix[33][87] * vector[33] +matrix[34][87] * vector[34] +matrix[35][87] * vector[35] +matrix[36][87] * vector[36] +matrix[37][87] * vector[37] +matrix[38][87] * vector[38] +matrix[39][87] * vector[39] +matrix[40][87] * vector[40] +matrix[41][87] * vector[41] +matrix[42][87] * vector[42] +matrix[43][87] * vector[43] +matrix[44][87] * vector[44] +matrix[45][87] * vector[45] +matrix[46][87] * vector[46] +matrix[47][87] * vector[47] +matrix[48][87] * vector[48] +matrix[49][87] * vector[49] +matrix[50][87] * vector[50] +matrix[51][87] * vector[51] +matrix[52][87] * vector[52] +matrix[53][87] * vector[53] +matrix[54][87] * vector[54] +matrix[55][87] * vector[55] +matrix[56][87] * vector[56] +matrix[57][87] * vector[57] +matrix[58][87] * vector[58] +matrix[59][87] * vector[59] +matrix[60][87] * vector[60] +matrix[61][87] * vector[61] +matrix[62][87] * vector[62] +matrix[63][87] * vector[63] +matrix[64][87] * vector[64] +matrix[65][87] * vector[65] +matrix[66][87] * vector[66] +matrix[67][87] * vector[67] +matrix[68][87] * vector[68] +matrix[69][87] * vector[69] +matrix[70][87] * vector[70] +matrix[71][87] * vector[71] +matrix[72][87] * vector[72] +matrix[73][87] * vector[73] +matrix[74][87] * vector[74] +matrix[75][87] * vector[75] +matrix[76][87] * vector[76] +matrix[77][87] * vector[77] +matrix[78][87] * vector[78] +matrix[79][87] * vector[79] +matrix[80][87] * vector[80] +matrix[81][87] * vector[81] +matrix[82][87] * vector[82] +matrix[83][87] * vector[83] +matrix[84][87] * vector[84] +matrix[85][87] * vector[85] +matrix[86][87] * vector[86] +matrix[87][87] * vector[87] +matrix[88][87] * vector[88] +matrix[89][87] * vector[89] +matrix[90][87] * vector[90] +matrix[91][87] * vector[91] +matrix[92][87] * vector[92] +matrix[93][87] * vector[93] +matrix[94][87] * vector[94] +matrix[95][87] * vector[95] +matrix[96][87] * vector[96] +matrix[97][87] * vector[97] +matrix[98][87] * vector[98] +matrix[99][87] * vector[99] +b[87];
assign result[88] = matrix[0][88] * vector[0] +matrix[1][88] * vector[1] +matrix[2][88] * vector[2] +matrix[3][88] * vector[3] +matrix[4][88] * vector[4] +matrix[5][88] * vector[5] +matrix[6][88] * vector[6] +matrix[7][88] * vector[7] +matrix[8][88] * vector[8] +matrix[9][88] * vector[9] +matrix[10][88] * vector[10] +matrix[11][88] * vector[11] +matrix[12][88] * vector[12] +matrix[13][88] * vector[13] +matrix[14][88] * vector[14] +matrix[15][88] * vector[15] +matrix[16][88] * vector[16] +matrix[17][88] * vector[17] +matrix[18][88] * vector[18] +matrix[19][88] * vector[19] +matrix[20][88] * vector[20] +matrix[21][88] * vector[21] +matrix[22][88] * vector[22] +matrix[23][88] * vector[23] +matrix[24][88] * vector[24] +matrix[25][88] * vector[25] +matrix[26][88] * vector[26] +matrix[27][88] * vector[27] +matrix[28][88] * vector[28] +matrix[29][88] * vector[29] +matrix[30][88] * vector[30] +matrix[31][88] * vector[31] +matrix[32][88] * vector[32] +matrix[33][88] * vector[33] +matrix[34][88] * vector[34] +matrix[35][88] * vector[35] +matrix[36][88] * vector[36] +matrix[37][88] * vector[37] +matrix[38][88] * vector[38] +matrix[39][88] * vector[39] +matrix[40][88] * vector[40] +matrix[41][88] * vector[41] +matrix[42][88] * vector[42] +matrix[43][88] * vector[43] +matrix[44][88] * vector[44] +matrix[45][88] * vector[45] +matrix[46][88] * vector[46] +matrix[47][88] * vector[47] +matrix[48][88] * vector[48] +matrix[49][88] * vector[49] +matrix[50][88] * vector[50] +matrix[51][88] * vector[51] +matrix[52][88] * vector[52] +matrix[53][88] * vector[53] +matrix[54][88] * vector[54] +matrix[55][88] * vector[55] +matrix[56][88] * vector[56] +matrix[57][88] * vector[57] +matrix[58][88] * vector[58] +matrix[59][88] * vector[59] +matrix[60][88] * vector[60] +matrix[61][88] * vector[61] +matrix[62][88] * vector[62] +matrix[63][88] * vector[63] +matrix[64][88] * vector[64] +matrix[65][88] * vector[65] +matrix[66][88] * vector[66] +matrix[67][88] * vector[67] +matrix[68][88] * vector[68] +matrix[69][88] * vector[69] +matrix[70][88] * vector[70] +matrix[71][88] * vector[71] +matrix[72][88] * vector[72] +matrix[73][88] * vector[73] +matrix[74][88] * vector[74] +matrix[75][88] * vector[75] +matrix[76][88] * vector[76] +matrix[77][88] * vector[77] +matrix[78][88] * vector[78] +matrix[79][88] * vector[79] +matrix[80][88] * vector[80] +matrix[81][88] * vector[81] +matrix[82][88] * vector[82] +matrix[83][88] * vector[83] +matrix[84][88] * vector[84] +matrix[85][88] * vector[85] +matrix[86][88] * vector[86] +matrix[87][88] * vector[87] +matrix[88][88] * vector[88] +matrix[89][88] * vector[89] +matrix[90][88] * vector[90] +matrix[91][88] * vector[91] +matrix[92][88] * vector[92] +matrix[93][88] * vector[93] +matrix[94][88] * vector[94] +matrix[95][88] * vector[95] +matrix[96][88] * vector[96] +matrix[97][88] * vector[97] +matrix[98][88] * vector[98] +matrix[99][88] * vector[99] +b[88];
assign result[89] = matrix[0][89] * vector[0] +matrix[1][89] * vector[1] +matrix[2][89] * vector[2] +matrix[3][89] * vector[3] +matrix[4][89] * vector[4] +matrix[5][89] * vector[5] +matrix[6][89] * vector[6] +matrix[7][89] * vector[7] +matrix[8][89] * vector[8] +matrix[9][89] * vector[9] +matrix[10][89] * vector[10] +matrix[11][89] * vector[11] +matrix[12][89] * vector[12] +matrix[13][89] * vector[13] +matrix[14][89] * vector[14] +matrix[15][89] * vector[15] +matrix[16][89] * vector[16] +matrix[17][89] * vector[17] +matrix[18][89] * vector[18] +matrix[19][89] * vector[19] +matrix[20][89] * vector[20] +matrix[21][89] * vector[21] +matrix[22][89] * vector[22] +matrix[23][89] * vector[23] +matrix[24][89] * vector[24] +matrix[25][89] * vector[25] +matrix[26][89] * vector[26] +matrix[27][89] * vector[27] +matrix[28][89] * vector[28] +matrix[29][89] * vector[29] +matrix[30][89] * vector[30] +matrix[31][89] * vector[31] +matrix[32][89] * vector[32] +matrix[33][89] * vector[33] +matrix[34][89] * vector[34] +matrix[35][89] * vector[35] +matrix[36][89] * vector[36] +matrix[37][89] * vector[37] +matrix[38][89] * vector[38] +matrix[39][89] * vector[39] +matrix[40][89] * vector[40] +matrix[41][89] * vector[41] +matrix[42][89] * vector[42] +matrix[43][89] * vector[43] +matrix[44][89] * vector[44] +matrix[45][89] * vector[45] +matrix[46][89] * vector[46] +matrix[47][89] * vector[47] +matrix[48][89] * vector[48] +matrix[49][89] * vector[49] +matrix[50][89] * vector[50] +matrix[51][89] * vector[51] +matrix[52][89] * vector[52] +matrix[53][89] * vector[53] +matrix[54][89] * vector[54] +matrix[55][89] * vector[55] +matrix[56][89] * vector[56] +matrix[57][89] * vector[57] +matrix[58][89] * vector[58] +matrix[59][89] * vector[59] +matrix[60][89] * vector[60] +matrix[61][89] * vector[61] +matrix[62][89] * vector[62] +matrix[63][89] * vector[63] +matrix[64][89] * vector[64] +matrix[65][89] * vector[65] +matrix[66][89] * vector[66] +matrix[67][89] * vector[67] +matrix[68][89] * vector[68] +matrix[69][89] * vector[69] +matrix[70][89] * vector[70] +matrix[71][89] * vector[71] +matrix[72][89] * vector[72] +matrix[73][89] * vector[73] +matrix[74][89] * vector[74] +matrix[75][89] * vector[75] +matrix[76][89] * vector[76] +matrix[77][89] * vector[77] +matrix[78][89] * vector[78] +matrix[79][89] * vector[79] +matrix[80][89] * vector[80] +matrix[81][89] * vector[81] +matrix[82][89] * vector[82] +matrix[83][89] * vector[83] +matrix[84][89] * vector[84] +matrix[85][89] * vector[85] +matrix[86][89] * vector[86] +matrix[87][89] * vector[87] +matrix[88][89] * vector[88] +matrix[89][89] * vector[89] +matrix[90][89] * vector[90] +matrix[91][89] * vector[91] +matrix[92][89] * vector[92] +matrix[93][89] * vector[93] +matrix[94][89] * vector[94] +matrix[95][89] * vector[95] +matrix[96][89] * vector[96] +matrix[97][89] * vector[97] +matrix[98][89] * vector[98] +matrix[99][89] * vector[99] +b[89];
assign result[90] = matrix[0][90] * vector[0] +matrix[1][90] * vector[1] +matrix[2][90] * vector[2] +matrix[3][90] * vector[3] +matrix[4][90] * vector[4] +matrix[5][90] * vector[5] +matrix[6][90] * vector[6] +matrix[7][90] * vector[7] +matrix[8][90] * vector[8] +matrix[9][90] * vector[9] +matrix[10][90] * vector[10] +matrix[11][90] * vector[11] +matrix[12][90] * vector[12] +matrix[13][90] * vector[13] +matrix[14][90] * vector[14] +matrix[15][90] * vector[15] +matrix[16][90] * vector[16] +matrix[17][90] * vector[17] +matrix[18][90] * vector[18] +matrix[19][90] * vector[19] +matrix[20][90] * vector[20] +matrix[21][90] * vector[21] +matrix[22][90] * vector[22] +matrix[23][90] * vector[23] +matrix[24][90] * vector[24] +matrix[25][90] * vector[25] +matrix[26][90] * vector[26] +matrix[27][90] * vector[27] +matrix[28][90] * vector[28] +matrix[29][90] * vector[29] +matrix[30][90] * vector[30] +matrix[31][90] * vector[31] +matrix[32][90] * vector[32] +matrix[33][90] * vector[33] +matrix[34][90] * vector[34] +matrix[35][90] * vector[35] +matrix[36][90] * vector[36] +matrix[37][90] * vector[37] +matrix[38][90] * vector[38] +matrix[39][90] * vector[39] +matrix[40][90] * vector[40] +matrix[41][90] * vector[41] +matrix[42][90] * vector[42] +matrix[43][90] * vector[43] +matrix[44][90] * vector[44] +matrix[45][90] * vector[45] +matrix[46][90] * vector[46] +matrix[47][90] * vector[47] +matrix[48][90] * vector[48] +matrix[49][90] * vector[49] +matrix[50][90] * vector[50] +matrix[51][90] * vector[51] +matrix[52][90] * vector[52] +matrix[53][90] * vector[53] +matrix[54][90] * vector[54] +matrix[55][90] * vector[55] +matrix[56][90] * vector[56] +matrix[57][90] * vector[57] +matrix[58][90] * vector[58] +matrix[59][90] * vector[59] +matrix[60][90] * vector[60] +matrix[61][90] * vector[61] +matrix[62][90] * vector[62] +matrix[63][90] * vector[63] +matrix[64][90] * vector[64] +matrix[65][90] * vector[65] +matrix[66][90] * vector[66] +matrix[67][90] * vector[67] +matrix[68][90] * vector[68] +matrix[69][90] * vector[69] +matrix[70][90] * vector[70] +matrix[71][90] * vector[71] +matrix[72][90] * vector[72] +matrix[73][90] * vector[73] +matrix[74][90] * vector[74] +matrix[75][90] * vector[75] +matrix[76][90] * vector[76] +matrix[77][90] * vector[77] +matrix[78][90] * vector[78] +matrix[79][90] * vector[79] +matrix[80][90] * vector[80] +matrix[81][90] * vector[81] +matrix[82][90] * vector[82] +matrix[83][90] * vector[83] +matrix[84][90] * vector[84] +matrix[85][90] * vector[85] +matrix[86][90] * vector[86] +matrix[87][90] * vector[87] +matrix[88][90] * vector[88] +matrix[89][90] * vector[89] +matrix[90][90] * vector[90] +matrix[91][90] * vector[91] +matrix[92][90] * vector[92] +matrix[93][90] * vector[93] +matrix[94][90] * vector[94] +matrix[95][90] * vector[95] +matrix[96][90] * vector[96] +matrix[97][90] * vector[97] +matrix[98][90] * vector[98] +matrix[99][90] * vector[99] +b[90];
assign result[91] = matrix[0][91] * vector[0] +matrix[1][91] * vector[1] +matrix[2][91] * vector[2] +matrix[3][91] * vector[3] +matrix[4][91] * vector[4] +matrix[5][91] * vector[5] +matrix[6][91] * vector[6] +matrix[7][91] * vector[7] +matrix[8][91] * vector[8] +matrix[9][91] * vector[9] +matrix[10][91] * vector[10] +matrix[11][91] * vector[11] +matrix[12][91] * vector[12] +matrix[13][91] * vector[13] +matrix[14][91] * vector[14] +matrix[15][91] * vector[15] +matrix[16][91] * vector[16] +matrix[17][91] * vector[17] +matrix[18][91] * vector[18] +matrix[19][91] * vector[19] +matrix[20][91] * vector[20] +matrix[21][91] * vector[21] +matrix[22][91] * vector[22] +matrix[23][91] * vector[23] +matrix[24][91] * vector[24] +matrix[25][91] * vector[25] +matrix[26][91] * vector[26] +matrix[27][91] * vector[27] +matrix[28][91] * vector[28] +matrix[29][91] * vector[29] +matrix[30][91] * vector[30] +matrix[31][91] * vector[31] +matrix[32][91] * vector[32] +matrix[33][91] * vector[33] +matrix[34][91] * vector[34] +matrix[35][91] * vector[35] +matrix[36][91] * vector[36] +matrix[37][91] * vector[37] +matrix[38][91] * vector[38] +matrix[39][91] * vector[39] +matrix[40][91] * vector[40] +matrix[41][91] * vector[41] +matrix[42][91] * vector[42] +matrix[43][91] * vector[43] +matrix[44][91] * vector[44] +matrix[45][91] * vector[45] +matrix[46][91] * vector[46] +matrix[47][91] * vector[47] +matrix[48][91] * vector[48] +matrix[49][91] * vector[49] +matrix[50][91] * vector[50] +matrix[51][91] * vector[51] +matrix[52][91] * vector[52] +matrix[53][91] * vector[53] +matrix[54][91] * vector[54] +matrix[55][91] * vector[55] +matrix[56][91] * vector[56] +matrix[57][91] * vector[57] +matrix[58][91] * vector[58] +matrix[59][91] * vector[59] +matrix[60][91] * vector[60] +matrix[61][91] * vector[61] +matrix[62][91] * vector[62] +matrix[63][91] * vector[63] +matrix[64][91] * vector[64] +matrix[65][91] * vector[65] +matrix[66][91] * vector[66] +matrix[67][91] * vector[67] +matrix[68][91] * vector[68] +matrix[69][91] * vector[69] +matrix[70][91] * vector[70] +matrix[71][91] * vector[71] +matrix[72][91] * vector[72] +matrix[73][91] * vector[73] +matrix[74][91] * vector[74] +matrix[75][91] * vector[75] +matrix[76][91] * vector[76] +matrix[77][91] * vector[77] +matrix[78][91] * vector[78] +matrix[79][91] * vector[79] +matrix[80][91] * vector[80] +matrix[81][91] * vector[81] +matrix[82][91] * vector[82] +matrix[83][91] * vector[83] +matrix[84][91] * vector[84] +matrix[85][91] * vector[85] +matrix[86][91] * vector[86] +matrix[87][91] * vector[87] +matrix[88][91] * vector[88] +matrix[89][91] * vector[89] +matrix[90][91] * vector[90] +matrix[91][91] * vector[91] +matrix[92][91] * vector[92] +matrix[93][91] * vector[93] +matrix[94][91] * vector[94] +matrix[95][91] * vector[95] +matrix[96][91] * vector[96] +matrix[97][91] * vector[97] +matrix[98][91] * vector[98] +matrix[99][91] * vector[99] +b[91];
assign result[92] = matrix[0][92] * vector[0] +matrix[1][92] * vector[1] +matrix[2][92] * vector[2] +matrix[3][92] * vector[3] +matrix[4][92] * vector[4] +matrix[5][92] * vector[5] +matrix[6][92] * vector[6] +matrix[7][92] * vector[7] +matrix[8][92] * vector[8] +matrix[9][92] * vector[9] +matrix[10][92] * vector[10] +matrix[11][92] * vector[11] +matrix[12][92] * vector[12] +matrix[13][92] * vector[13] +matrix[14][92] * vector[14] +matrix[15][92] * vector[15] +matrix[16][92] * vector[16] +matrix[17][92] * vector[17] +matrix[18][92] * vector[18] +matrix[19][92] * vector[19] +matrix[20][92] * vector[20] +matrix[21][92] * vector[21] +matrix[22][92] * vector[22] +matrix[23][92] * vector[23] +matrix[24][92] * vector[24] +matrix[25][92] * vector[25] +matrix[26][92] * vector[26] +matrix[27][92] * vector[27] +matrix[28][92] * vector[28] +matrix[29][92] * vector[29] +matrix[30][92] * vector[30] +matrix[31][92] * vector[31] +matrix[32][92] * vector[32] +matrix[33][92] * vector[33] +matrix[34][92] * vector[34] +matrix[35][92] * vector[35] +matrix[36][92] * vector[36] +matrix[37][92] * vector[37] +matrix[38][92] * vector[38] +matrix[39][92] * vector[39] +matrix[40][92] * vector[40] +matrix[41][92] * vector[41] +matrix[42][92] * vector[42] +matrix[43][92] * vector[43] +matrix[44][92] * vector[44] +matrix[45][92] * vector[45] +matrix[46][92] * vector[46] +matrix[47][92] * vector[47] +matrix[48][92] * vector[48] +matrix[49][92] * vector[49] +matrix[50][92] * vector[50] +matrix[51][92] * vector[51] +matrix[52][92] * vector[52] +matrix[53][92] * vector[53] +matrix[54][92] * vector[54] +matrix[55][92] * vector[55] +matrix[56][92] * vector[56] +matrix[57][92] * vector[57] +matrix[58][92] * vector[58] +matrix[59][92] * vector[59] +matrix[60][92] * vector[60] +matrix[61][92] * vector[61] +matrix[62][92] * vector[62] +matrix[63][92] * vector[63] +matrix[64][92] * vector[64] +matrix[65][92] * vector[65] +matrix[66][92] * vector[66] +matrix[67][92] * vector[67] +matrix[68][92] * vector[68] +matrix[69][92] * vector[69] +matrix[70][92] * vector[70] +matrix[71][92] * vector[71] +matrix[72][92] * vector[72] +matrix[73][92] * vector[73] +matrix[74][92] * vector[74] +matrix[75][92] * vector[75] +matrix[76][92] * vector[76] +matrix[77][92] * vector[77] +matrix[78][92] * vector[78] +matrix[79][92] * vector[79] +matrix[80][92] * vector[80] +matrix[81][92] * vector[81] +matrix[82][92] * vector[82] +matrix[83][92] * vector[83] +matrix[84][92] * vector[84] +matrix[85][92] * vector[85] +matrix[86][92] * vector[86] +matrix[87][92] * vector[87] +matrix[88][92] * vector[88] +matrix[89][92] * vector[89] +matrix[90][92] * vector[90] +matrix[91][92] * vector[91] +matrix[92][92] * vector[92] +matrix[93][92] * vector[93] +matrix[94][92] * vector[94] +matrix[95][92] * vector[95] +matrix[96][92] * vector[96] +matrix[97][92] * vector[97] +matrix[98][92] * vector[98] +matrix[99][92] * vector[99] +b[92];
assign result[93] = matrix[0][93] * vector[0] +matrix[1][93] * vector[1] +matrix[2][93] * vector[2] +matrix[3][93] * vector[3] +matrix[4][93] * vector[4] +matrix[5][93] * vector[5] +matrix[6][93] * vector[6] +matrix[7][93] * vector[7] +matrix[8][93] * vector[8] +matrix[9][93] * vector[9] +matrix[10][93] * vector[10] +matrix[11][93] * vector[11] +matrix[12][93] * vector[12] +matrix[13][93] * vector[13] +matrix[14][93] * vector[14] +matrix[15][93] * vector[15] +matrix[16][93] * vector[16] +matrix[17][93] * vector[17] +matrix[18][93] * vector[18] +matrix[19][93] * vector[19] +matrix[20][93] * vector[20] +matrix[21][93] * vector[21] +matrix[22][93] * vector[22] +matrix[23][93] * vector[23] +matrix[24][93] * vector[24] +matrix[25][93] * vector[25] +matrix[26][93] * vector[26] +matrix[27][93] * vector[27] +matrix[28][93] * vector[28] +matrix[29][93] * vector[29] +matrix[30][93] * vector[30] +matrix[31][93] * vector[31] +matrix[32][93] * vector[32] +matrix[33][93] * vector[33] +matrix[34][93] * vector[34] +matrix[35][93] * vector[35] +matrix[36][93] * vector[36] +matrix[37][93] * vector[37] +matrix[38][93] * vector[38] +matrix[39][93] * vector[39] +matrix[40][93] * vector[40] +matrix[41][93] * vector[41] +matrix[42][93] * vector[42] +matrix[43][93] * vector[43] +matrix[44][93] * vector[44] +matrix[45][93] * vector[45] +matrix[46][93] * vector[46] +matrix[47][93] * vector[47] +matrix[48][93] * vector[48] +matrix[49][93] * vector[49] +matrix[50][93] * vector[50] +matrix[51][93] * vector[51] +matrix[52][93] * vector[52] +matrix[53][93] * vector[53] +matrix[54][93] * vector[54] +matrix[55][93] * vector[55] +matrix[56][93] * vector[56] +matrix[57][93] * vector[57] +matrix[58][93] * vector[58] +matrix[59][93] * vector[59] +matrix[60][93] * vector[60] +matrix[61][93] * vector[61] +matrix[62][93] * vector[62] +matrix[63][93] * vector[63] +matrix[64][93] * vector[64] +matrix[65][93] * vector[65] +matrix[66][93] * vector[66] +matrix[67][93] * vector[67] +matrix[68][93] * vector[68] +matrix[69][93] * vector[69] +matrix[70][93] * vector[70] +matrix[71][93] * vector[71] +matrix[72][93] * vector[72] +matrix[73][93] * vector[73] +matrix[74][93] * vector[74] +matrix[75][93] * vector[75] +matrix[76][93] * vector[76] +matrix[77][93] * vector[77] +matrix[78][93] * vector[78] +matrix[79][93] * vector[79] +matrix[80][93] * vector[80] +matrix[81][93] * vector[81] +matrix[82][93] * vector[82] +matrix[83][93] * vector[83] +matrix[84][93] * vector[84] +matrix[85][93] * vector[85] +matrix[86][93] * vector[86] +matrix[87][93] * vector[87] +matrix[88][93] * vector[88] +matrix[89][93] * vector[89] +matrix[90][93] * vector[90] +matrix[91][93] * vector[91] +matrix[92][93] * vector[92] +matrix[93][93] * vector[93] +matrix[94][93] * vector[94] +matrix[95][93] * vector[95] +matrix[96][93] * vector[96] +matrix[97][93] * vector[97] +matrix[98][93] * vector[98] +matrix[99][93] * vector[99] +b[93];
assign result[94] = matrix[0][94] * vector[0] +matrix[1][94] * vector[1] +matrix[2][94] * vector[2] +matrix[3][94] * vector[3] +matrix[4][94] * vector[4] +matrix[5][94] * vector[5] +matrix[6][94] * vector[6] +matrix[7][94] * vector[7] +matrix[8][94] * vector[8] +matrix[9][94] * vector[9] +matrix[10][94] * vector[10] +matrix[11][94] * vector[11] +matrix[12][94] * vector[12] +matrix[13][94] * vector[13] +matrix[14][94] * vector[14] +matrix[15][94] * vector[15] +matrix[16][94] * vector[16] +matrix[17][94] * vector[17] +matrix[18][94] * vector[18] +matrix[19][94] * vector[19] +matrix[20][94] * vector[20] +matrix[21][94] * vector[21] +matrix[22][94] * vector[22] +matrix[23][94] * vector[23] +matrix[24][94] * vector[24] +matrix[25][94] * vector[25] +matrix[26][94] * vector[26] +matrix[27][94] * vector[27] +matrix[28][94] * vector[28] +matrix[29][94] * vector[29] +matrix[30][94] * vector[30] +matrix[31][94] * vector[31] +matrix[32][94] * vector[32] +matrix[33][94] * vector[33] +matrix[34][94] * vector[34] +matrix[35][94] * vector[35] +matrix[36][94] * vector[36] +matrix[37][94] * vector[37] +matrix[38][94] * vector[38] +matrix[39][94] * vector[39] +matrix[40][94] * vector[40] +matrix[41][94] * vector[41] +matrix[42][94] * vector[42] +matrix[43][94] * vector[43] +matrix[44][94] * vector[44] +matrix[45][94] * vector[45] +matrix[46][94] * vector[46] +matrix[47][94] * vector[47] +matrix[48][94] * vector[48] +matrix[49][94] * vector[49] +matrix[50][94] * vector[50] +matrix[51][94] * vector[51] +matrix[52][94] * vector[52] +matrix[53][94] * vector[53] +matrix[54][94] * vector[54] +matrix[55][94] * vector[55] +matrix[56][94] * vector[56] +matrix[57][94] * vector[57] +matrix[58][94] * vector[58] +matrix[59][94] * vector[59] +matrix[60][94] * vector[60] +matrix[61][94] * vector[61] +matrix[62][94] * vector[62] +matrix[63][94] * vector[63] +matrix[64][94] * vector[64] +matrix[65][94] * vector[65] +matrix[66][94] * vector[66] +matrix[67][94] * vector[67] +matrix[68][94] * vector[68] +matrix[69][94] * vector[69] +matrix[70][94] * vector[70] +matrix[71][94] * vector[71] +matrix[72][94] * vector[72] +matrix[73][94] * vector[73] +matrix[74][94] * vector[74] +matrix[75][94] * vector[75] +matrix[76][94] * vector[76] +matrix[77][94] * vector[77] +matrix[78][94] * vector[78] +matrix[79][94] * vector[79] +matrix[80][94] * vector[80] +matrix[81][94] * vector[81] +matrix[82][94] * vector[82] +matrix[83][94] * vector[83] +matrix[84][94] * vector[84] +matrix[85][94] * vector[85] +matrix[86][94] * vector[86] +matrix[87][94] * vector[87] +matrix[88][94] * vector[88] +matrix[89][94] * vector[89] +matrix[90][94] * vector[90] +matrix[91][94] * vector[91] +matrix[92][94] * vector[92] +matrix[93][94] * vector[93] +matrix[94][94] * vector[94] +matrix[95][94] * vector[95] +matrix[96][94] * vector[96] +matrix[97][94] * vector[97] +matrix[98][94] * vector[98] +matrix[99][94] * vector[99] +b[94];
assign result[95] = matrix[0][95] * vector[0] +matrix[1][95] * vector[1] +matrix[2][95] * vector[2] +matrix[3][95] * vector[3] +matrix[4][95] * vector[4] +matrix[5][95] * vector[5] +matrix[6][95] * vector[6] +matrix[7][95] * vector[7] +matrix[8][95] * vector[8] +matrix[9][95] * vector[9] +matrix[10][95] * vector[10] +matrix[11][95] * vector[11] +matrix[12][95] * vector[12] +matrix[13][95] * vector[13] +matrix[14][95] * vector[14] +matrix[15][95] * vector[15] +matrix[16][95] * vector[16] +matrix[17][95] * vector[17] +matrix[18][95] * vector[18] +matrix[19][95] * vector[19] +matrix[20][95] * vector[20] +matrix[21][95] * vector[21] +matrix[22][95] * vector[22] +matrix[23][95] * vector[23] +matrix[24][95] * vector[24] +matrix[25][95] * vector[25] +matrix[26][95] * vector[26] +matrix[27][95] * vector[27] +matrix[28][95] * vector[28] +matrix[29][95] * vector[29] +matrix[30][95] * vector[30] +matrix[31][95] * vector[31] +matrix[32][95] * vector[32] +matrix[33][95] * vector[33] +matrix[34][95] * vector[34] +matrix[35][95] * vector[35] +matrix[36][95] * vector[36] +matrix[37][95] * vector[37] +matrix[38][95] * vector[38] +matrix[39][95] * vector[39] +matrix[40][95] * vector[40] +matrix[41][95] * vector[41] +matrix[42][95] * vector[42] +matrix[43][95] * vector[43] +matrix[44][95] * vector[44] +matrix[45][95] * vector[45] +matrix[46][95] * vector[46] +matrix[47][95] * vector[47] +matrix[48][95] * vector[48] +matrix[49][95] * vector[49] +matrix[50][95] * vector[50] +matrix[51][95] * vector[51] +matrix[52][95] * vector[52] +matrix[53][95] * vector[53] +matrix[54][95] * vector[54] +matrix[55][95] * vector[55] +matrix[56][95] * vector[56] +matrix[57][95] * vector[57] +matrix[58][95] * vector[58] +matrix[59][95] * vector[59] +matrix[60][95] * vector[60] +matrix[61][95] * vector[61] +matrix[62][95] * vector[62] +matrix[63][95] * vector[63] +matrix[64][95] * vector[64] +matrix[65][95] * vector[65] +matrix[66][95] * vector[66] +matrix[67][95] * vector[67] +matrix[68][95] * vector[68] +matrix[69][95] * vector[69] +matrix[70][95] * vector[70] +matrix[71][95] * vector[71] +matrix[72][95] * vector[72] +matrix[73][95] * vector[73] +matrix[74][95] * vector[74] +matrix[75][95] * vector[75] +matrix[76][95] * vector[76] +matrix[77][95] * vector[77] +matrix[78][95] * vector[78] +matrix[79][95] * vector[79] +matrix[80][95] * vector[80] +matrix[81][95] * vector[81] +matrix[82][95] * vector[82] +matrix[83][95] * vector[83] +matrix[84][95] * vector[84] +matrix[85][95] * vector[85] +matrix[86][95] * vector[86] +matrix[87][95] * vector[87] +matrix[88][95] * vector[88] +matrix[89][95] * vector[89] +matrix[90][95] * vector[90] +matrix[91][95] * vector[91] +matrix[92][95] * vector[92] +matrix[93][95] * vector[93] +matrix[94][95] * vector[94] +matrix[95][95] * vector[95] +matrix[96][95] * vector[96] +matrix[97][95] * vector[97] +matrix[98][95] * vector[98] +matrix[99][95] * vector[99] +b[95];
assign result[96] = matrix[0][96] * vector[0] +matrix[1][96] * vector[1] +matrix[2][96] * vector[2] +matrix[3][96] * vector[3] +matrix[4][96] * vector[4] +matrix[5][96] * vector[5] +matrix[6][96] * vector[6] +matrix[7][96] * vector[7] +matrix[8][96] * vector[8] +matrix[9][96] * vector[9] +matrix[10][96] * vector[10] +matrix[11][96] * vector[11] +matrix[12][96] * vector[12] +matrix[13][96] * vector[13] +matrix[14][96] * vector[14] +matrix[15][96] * vector[15] +matrix[16][96] * vector[16] +matrix[17][96] * vector[17] +matrix[18][96] * vector[18] +matrix[19][96] * vector[19] +matrix[20][96] * vector[20] +matrix[21][96] * vector[21] +matrix[22][96] * vector[22] +matrix[23][96] * vector[23] +matrix[24][96] * vector[24] +matrix[25][96] * vector[25] +matrix[26][96] * vector[26] +matrix[27][96] * vector[27] +matrix[28][96] * vector[28] +matrix[29][96] * vector[29] +matrix[30][96] * vector[30] +matrix[31][96] * vector[31] +matrix[32][96] * vector[32] +matrix[33][96] * vector[33] +matrix[34][96] * vector[34] +matrix[35][96] * vector[35] +matrix[36][96] * vector[36] +matrix[37][96] * vector[37] +matrix[38][96] * vector[38] +matrix[39][96] * vector[39] +matrix[40][96] * vector[40] +matrix[41][96] * vector[41] +matrix[42][96] * vector[42] +matrix[43][96] * vector[43] +matrix[44][96] * vector[44] +matrix[45][96] * vector[45] +matrix[46][96] * vector[46] +matrix[47][96] * vector[47] +matrix[48][96] * vector[48] +matrix[49][96] * vector[49] +matrix[50][96] * vector[50] +matrix[51][96] * vector[51] +matrix[52][96] * vector[52] +matrix[53][96] * vector[53] +matrix[54][96] * vector[54] +matrix[55][96] * vector[55] +matrix[56][96] * vector[56] +matrix[57][96] * vector[57] +matrix[58][96] * vector[58] +matrix[59][96] * vector[59] +matrix[60][96] * vector[60] +matrix[61][96] * vector[61] +matrix[62][96] * vector[62] +matrix[63][96] * vector[63] +matrix[64][96] * vector[64] +matrix[65][96] * vector[65] +matrix[66][96] * vector[66] +matrix[67][96] * vector[67] +matrix[68][96] * vector[68] +matrix[69][96] * vector[69] +matrix[70][96] * vector[70] +matrix[71][96] * vector[71] +matrix[72][96] * vector[72] +matrix[73][96] * vector[73] +matrix[74][96] * vector[74] +matrix[75][96] * vector[75] +matrix[76][96] * vector[76] +matrix[77][96] * vector[77] +matrix[78][96] * vector[78] +matrix[79][96] * vector[79] +matrix[80][96] * vector[80] +matrix[81][96] * vector[81] +matrix[82][96] * vector[82] +matrix[83][96] * vector[83] +matrix[84][96] * vector[84] +matrix[85][96] * vector[85] +matrix[86][96] * vector[86] +matrix[87][96] * vector[87] +matrix[88][96] * vector[88] +matrix[89][96] * vector[89] +matrix[90][96] * vector[90] +matrix[91][96] * vector[91] +matrix[92][96] * vector[92] +matrix[93][96] * vector[93] +matrix[94][96] * vector[94] +matrix[95][96] * vector[95] +matrix[96][96] * vector[96] +matrix[97][96] * vector[97] +matrix[98][96] * vector[98] +matrix[99][96] * vector[99] +b[96];
assign result[97] = matrix[0][97] * vector[0] +matrix[1][97] * vector[1] +matrix[2][97] * vector[2] +matrix[3][97] * vector[3] +matrix[4][97] * vector[4] +matrix[5][97] * vector[5] +matrix[6][97] * vector[6] +matrix[7][97] * vector[7] +matrix[8][97] * vector[8] +matrix[9][97] * vector[9] +matrix[10][97] * vector[10] +matrix[11][97] * vector[11] +matrix[12][97] * vector[12] +matrix[13][97] * vector[13] +matrix[14][97] * vector[14] +matrix[15][97] * vector[15] +matrix[16][97] * vector[16] +matrix[17][97] * vector[17] +matrix[18][97] * vector[18] +matrix[19][97] * vector[19] +matrix[20][97] * vector[20] +matrix[21][97] * vector[21] +matrix[22][97] * vector[22] +matrix[23][97] * vector[23] +matrix[24][97] * vector[24] +matrix[25][97] * vector[25] +matrix[26][97] * vector[26] +matrix[27][97] * vector[27] +matrix[28][97] * vector[28] +matrix[29][97] * vector[29] +matrix[30][97] * vector[30] +matrix[31][97] * vector[31] +matrix[32][97] * vector[32] +matrix[33][97] * vector[33] +matrix[34][97] * vector[34] +matrix[35][97] * vector[35] +matrix[36][97] * vector[36] +matrix[37][97] * vector[37] +matrix[38][97] * vector[38] +matrix[39][97] * vector[39] +matrix[40][97] * vector[40] +matrix[41][97] * vector[41] +matrix[42][97] * vector[42] +matrix[43][97] * vector[43] +matrix[44][97] * vector[44] +matrix[45][97] * vector[45] +matrix[46][97] * vector[46] +matrix[47][97] * vector[47] +matrix[48][97] * vector[48] +matrix[49][97] * vector[49] +matrix[50][97] * vector[50] +matrix[51][97] * vector[51] +matrix[52][97] * vector[52] +matrix[53][97] * vector[53] +matrix[54][97] * vector[54] +matrix[55][97] * vector[55] +matrix[56][97] * vector[56] +matrix[57][97] * vector[57] +matrix[58][97] * vector[58] +matrix[59][97] * vector[59] +matrix[60][97] * vector[60] +matrix[61][97] * vector[61] +matrix[62][97] * vector[62] +matrix[63][97] * vector[63] +matrix[64][97] * vector[64] +matrix[65][97] * vector[65] +matrix[66][97] * vector[66] +matrix[67][97] * vector[67] +matrix[68][97] * vector[68] +matrix[69][97] * vector[69] +matrix[70][97] * vector[70] +matrix[71][97] * vector[71] +matrix[72][97] * vector[72] +matrix[73][97] * vector[73] +matrix[74][97] * vector[74] +matrix[75][97] * vector[75] +matrix[76][97] * vector[76] +matrix[77][97] * vector[77] +matrix[78][97] * vector[78] +matrix[79][97] * vector[79] +matrix[80][97] * vector[80] +matrix[81][97] * vector[81] +matrix[82][97] * vector[82] +matrix[83][97] * vector[83] +matrix[84][97] * vector[84] +matrix[85][97] * vector[85] +matrix[86][97] * vector[86] +matrix[87][97] * vector[87] +matrix[88][97] * vector[88] +matrix[89][97] * vector[89] +matrix[90][97] * vector[90] +matrix[91][97] * vector[91] +matrix[92][97] * vector[92] +matrix[93][97] * vector[93] +matrix[94][97] * vector[94] +matrix[95][97] * vector[95] +matrix[96][97] * vector[96] +matrix[97][97] * vector[97] +matrix[98][97] * vector[98] +matrix[99][97] * vector[99] +b[97];
assign result[98] = matrix[0][98] * vector[0] +matrix[1][98] * vector[1] +matrix[2][98] * vector[2] +matrix[3][98] * vector[3] +matrix[4][98] * vector[4] +matrix[5][98] * vector[5] +matrix[6][98] * vector[6] +matrix[7][98] * vector[7] +matrix[8][98] * vector[8] +matrix[9][98] * vector[9] +matrix[10][98] * vector[10] +matrix[11][98] * vector[11] +matrix[12][98] * vector[12] +matrix[13][98] * vector[13] +matrix[14][98] * vector[14] +matrix[15][98] * vector[15] +matrix[16][98] * vector[16] +matrix[17][98] * vector[17] +matrix[18][98] * vector[18] +matrix[19][98] * vector[19] +matrix[20][98] * vector[20] +matrix[21][98] * vector[21] +matrix[22][98] * vector[22] +matrix[23][98] * vector[23] +matrix[24][98] * vector[24] +matrix[25][98] * vector[25] +matrix[26][98] * vector[26] +matrix[27][98] * vector[27] +matrix[28][98] * vector[28] +matrix[29][98] * vector[29] +matrix[30][98] * vector[30] +matrix[31][98] * vector[31] +matrix[32][98] * vector[32] +matrix[33][98] * vector[33] +matrix[34][98] * vector[34] +matrix[35][98] * vector[35] +matrix[36][98] * vector[36] +matrix[37][98] * vector[37] +matrix[38][98] * vector[38] +matrix[39][98] * vector[39] +matrix[40][98] * vector[40] +matrix[41][98] * vector[41] +matrix[42][98] * vector[42] +matrix[43][98] * vector[43] +matrix[44][98] * vector[44] +matrix[45][98] * vector[45] +matrix[46][98] * vector[46] +matrix[47][98] * vector[47] +matrix[48][98] * vector[48] +matrix[49][98] * vector[49] +matrix[50][98] * vector[50] +matrix[51][98] * vector[51] +matrix[52][98] * vector[52] +matrix[53][98] * vector[53] +matrix[54][98] * vector[54] +matrix[55][98] * vector[55] +matrix[56][98] * vector[56] +matrix[57][98] * vector[57] +matrix[58][98] * vector[58] +matrix[59][98] * vector[59] +matrix[60][98] * vector[60] +matrix[61][98] * vector[61] +matrix[62][98] * vector[62] +matrix[63][98] * vector[63] +matrix[64][98] * vector[64] +matrix[65][98] * vector[65] +matrix[66][98] * vector[66] +matrix[67][98] * vector[67] +matrix[68][98] * vector[68] +matrix[69][98] * vector[69] +matrix[70][98] * vector[70] +matrix[71][98] * vector[71] +matrix[72][98] * vector[72] +matrix[73][98] * vector[73] +matrix[74][98] * vector[74] +matrix[75][98] * vector[75] +matrix[76][98] * vector[76] +matrix[77][98] * vector[77] +matrix[78][98] * vector[78] +matrix[79][98] * vector[79] +matrix[80][98] * vector[80] +matrix[81][98] * vector[81] +matrix[82][98] * vector[82] +matrix[83][98] * vector[83] +matrix[84][98] * vector[84] +matrix[85][98] * vector[85] +matrix[86][98] * vector[86] +matrix[87][98] * vector[87] +matrix[88][98] * vector[88] +matrix[89][98] * vector[89] +matrix[90][98] * vector[90] +matrix[91][98] * vector[91] +matrix[92][98] * vector[92] +matrix[93][98] * vector[93] +matrix[94][98] * vector[94] +matrix[95][98] * vector[95] +matrix[96][98] * vector[96] +matrix[97][98] * vector[97] +matrix[98][98] * vector[98] +matrix[99][98] * vector[99] +b[98];
assign result[99] = matrix[0][99] * vector[0] +matrix[1][99] * vector[1] +matrix[2][99] * vector[2] +matrix[3][99] * vector[3] +matrix[4][99] * vector[4] +matrix[5][99] * vector[5] +matrix[6][99] * vector[6] +matrix[7][99] * vector[7] +matrix[8][99] * vector[8] +matrix[9][99] * vector[9] +matrix[10][99] * vector[10] +matrix[11][99] * vector[11] +matrix[12][99] * vector[12] +matrix[13][99] * vector[13] +matrix[14][99] * vector[14] +matrix[15][99] * vector[15] +matrix[16][99] * vector[16] +matrix[17][99] * vector[17] +matrix[18][99] * vector[18] +matrix[19][99] * vector[19] +matrix[20][99] * vector[20] +matrix[21][99] * vector[21] +matrix[22][99] * vector[22] +matrix[23][99] * vector[23] +matrix[24][99] * vector[24] +matrix[25][99] * vector[25] +matrix[26][99] * vector[26] +matrix[27][99] * vector[27] +matrix[28][99] * vector[28] +matrix[29][99] * vector[29] +matrix[30][99] * vector[30] +matrix[31][99] * vector[31] +matrix[32][99] * vector[32] +matrix[33][99] * vector[33] +matrix[34][99] * vector[34] +matrix[35][99] * vector[35] +matrix[36][99] * vector[36] +matrix[37][99] * vector[37] +matrix[38][99] * vector[38] +matrix[39][99] * vector[39] +matrix[40][99] * vector[40] +matrix[41][99] * vector[41] +matrix[42][99] * vector[42] +matrix[43][99] * vector[43] +matrix[44][99] * vector[44] +matrix[45][99] * vector[45] +matrix[46][99] * vector[46] +matrix[47][99] * vector[47] +matrix[48][99] * vector[48] +matrix[49][99] * vector[49] +matrix[50][99] * vector[50] +matrix[51][99] * vector[51] +matrix[52][99] * vector[52] +matrix[53][99] * vector[53] +matrix[54][99] * vector[54] +matrix[55][99] * vector[55] +matrix[56][99] * vector[56] +matrix[57][99] * vector[57] +matrix[58][99] * vector[58] +matrix[59][99] * vector[59] +matrix[60][99] * vector[60] +matrix[61][99] * vector[61] +matrix[62][99] * vector[62] +matrix[63][99] * vector[63] +matrix[64][99] * vector[64] +matrix[65][99] * vector[65] +matrix[66][99] * vector[66] +matrix[67][99] * vector[67] +matrix[68][99] * vector[68] +matrix[69][99] * vector[69] +matrix[70][99] * vector[70] +matrix[71][99] * vector[71] +matrix[72][99] * vector[72] +matrix[73][99] * vector[73] +matrix[74][99] * vector[74] +matrix[75][99] * vector[75] +matrix[76][99] * vector[76] +matrix[77][99] * vector[77] +matrix[78][99] * vector[78] +matrix[79][99] * vector[79] +matrix[80][99] * vector[80] +matrix[81][99] * vector[81] +matrix[82][99] * vector[82] +matrix[83][99] * vector[83] +matrix[84][99] * vector[84] +matrix[85][99] * vector[85] +matrix[86][99] * vector[86] +matrix[87][99] * vector[87] +matrix[88][99] * vector[88] +matrix[89][99] * vector[89] +matrix[90][99] * vector[90] +matrix[91][99] * vector[91] +matrix[92][99] * vector[92] +matrix[93][99] * vector[93] +matrix[94][99] * vector[94] +matrix[95][99] * vector[95] +matrix[96][99] * vector[96] +matrix[97][99] * vector[97] +matrix[98][99] * vector[98] +matrix[99][99] * vector[99] +b[99];
assign result[100] = matrix[0][100] * vector[0] +matrix[1][100] * vector[1] +matrix[2][100] * vector[2] +matrix[3][100] * vector[3] +matrix[4][100] * vector[4] +matrix[5][100] * vector[5] +matrix[6][100] * vector[6] +matrix[7][100] * vector[7] +matrix[8][100] * vector[8] +matrix[9][100] * vector[9] +matrix[10][100] * vector[10] +matrix[11][100] * vector[11] +matrix[12][100] * vector[12] +matrix[13][100] * vector[13] +matrix[14][100] * vector[14] +matrix[15][100] * vector[15] +matrix[16][100] * vector[16] +matrix[17][100] * vector[17] +matrix[18][100] * vector[18] +matrix[19][100] * vector[19] +matrix[20][100] * vector[20] +matrix[21][100] * vector[21] +matrix[22][100] * vector[22] +matrix[23][100] * vector[23] +matrix[24][100] * vector[24] +matrix[25][100] * vector[25] +matrix[26][100] * vector[26] +matrix[27][100] * vector[27] +matrix[28][100] * vector[28] +matrix[29][100] * vector[29] +matrix[30][100] * vector[30] +matrix[31][100] * vector[31] +matrix[32][100] * vector[32] +matrix[33][100] * vector[33] +matrix[34][100] * vector[34] +matrix[35][100] * vector[35] +matrix[36][100] * vector[36] +matrix[37][100] * vector[37] +matrix[38][100] * vector[38] +matrix[39][100] * vector[39] +matrix[40][100] * vector[40] +matrix[41][100] * vector[41] +matrix[42][100] * vector[42] +matrix[43][100] * vector[43] +matrix[44][100] * vector[44] +matrix[45][100] * vector[45] +matrix[46][100] * vector[46] +matrix[47][100] * vector[47] +matrix[48][100] * vector[48] +matrix[49][100] * vector[49] +matrix[50][100] * vector[50] +matrix[51][100] * vector[51] +matrix[52][100] * vector[52] +matrix[53][100] * vector[53] +matrix[54][100] * vector[54] +matrix[55][100] * vector[55] +matrix[56][100] * vector[56] +matrix[57][100] * vector[57] +matrix[58][100] * vector[58] +matrix[59][100] * vector[59] +matrix[60][100] * vector[60] +matrix[61][100] * vector[61] +matrix[62][100] * vector[62] +matrix[63][100] * vector[63] +matrix[64][100] * vector[64] +matrix[65][100] * vector[65] +matrix[66][100] * vector[66] +matrix[67][100] * vector[67] +matrix[68][100] * vector[68] +matrix[69][100] * vector[69] +matrix[70][100] * vector[70] +matrix[71][100] * vector[71] +matrix[72][100] * vector[72] +matrix[73][100] * vector[73] +matrix[74][100] * vector[74] +matrix[75][100] * vector[75] +matrix[76][100] * vector[76] +matrix[77][100] * vector[77] +matrix[78][100] * vector[78] +matrix[79][100] * vector[79] +matrix[80][100] * vector[80] +matrix[81][100] * vector[81] +matrix[82][100] * vector[82] +matrix[83][100] * vector[83] +matrix[84][100] * vector[84] +matrix[85][100] * vector[85] +matrix[86][100] * vector[86] +matrix[87][100] * vector[87] +matrix[88][100] * vector[88] +matrix[89][100] * vector[89] +matrix[90][100] * vector[90] +matrix[91][100] * vector[91] +matrix[92][100] * vector[92] +matrix[93][100] * vector[93] +matrix[94][100] * vector[94] +matrix[95][100] * vector[95] +matrix[96][100] * vector[96] +matrix[97][100] * vector[97] +matrix[98][100] * vector[98] +matrix[99][100] * vector[99] +b[100];
assign result[101] = matrix[0][101] * vector[0] +matrix[1][101] * vector[1] +matrix[2][101] * vector[2] +matrix[3][101] * vector[3] +matrix[4][101] * vector[4] +matrix[5][101] * vector[5] +matrix[6][101] * vector[6] +matrix[7][101] * vector[7] +matrix[8][101] * vector[8] +matrix[9][101] * vector[9] +matrix[10][101] * vector[10] +matrix[11][101] * vector[11] +matrix[12][101] * vector[12] +matrix[13][101] * vector[13] +matrix[14][101] * vector[14] +matrix[15][101] * vector[15] +matrix[16][101] * vector[16] +matrix[17][101] * vector[17] +matrix[18][101] * vector[18] +matrix[19][101] * vector[19] +matrix[20][101] * vector[20] +matrix[21][101] * vector[21] +matrix[22][101] * vector[22] +matrix[23][101] * vector[23] +matrix[24][101] * vector[24] +matrix[25][101] * vector[25] +matrix[26][101] * vector[26] +matrix[27][101] * vector[27] +matrix[28][101] * vector[28] +matrix[29][101] * vector[29] +matrix[30][101] * vector[30] +matrix[31][101] * vector[31] +matrix[32][101] * vector[32] +matrix[33][101] * vector[33] +matrix[34][101] * vector[34] +matrix[35][101] * vector[35] +matrix[36][101] * vector[36] +matrix[37][101] * vector[37] +matrix[38][101] * vector[38] +matrix[39][101] * vector[39] +matrix[40][101] * vector[40] +matrix[41][101] * vector[41] +matrix[42][101] * vector[42] +matrix[43][101] * vector[43] +matrix[44][101] * vector[44] +matrix[45][101] * vector[45] +matrix[46][101] * vector[46] +matrix[47][101] * vector[47] +matrix[48][101] * vector[48] +matrix[49][101] * vector[49] +matrix[50][101] * vector[50] +matrix[51][101] * vector[51] +matrix[52][101] * vector[52] +matrix[53][101] * vector[53] +matrix[54][101] * vector[54] +matrix[55][101] * vector[55] +matrix[56][101] * vector[56] +matrix[57][101] * vector[57] +matrix[58][101] * vector[58] +matrix[59][101] * vector[59] +matrix[60][101] * vector[60] +matrix[61][101] * vector[61] +matrix[62][101] * vector[62] +matrix[63][101] * vector[63] +matrix[64][101] * vector[64] +matrix[65][101] * vector[65] +matrix[66][101] * vector[66] +matrix[67][101] * vector[67] +matrix[68][101] * vector[68] +matrix[69][101] * vector[69] +matrix[70][101] * vector[70] +matrix[71][101] * vector[71] +matrix[72][101] * vector[72] +matrix[73][101] * vector[73] +matrix[74][101] * vector[74] +matrix[75][101] * vector[75] +matrix[76][101] * vector[76] +matrix[77][101] * vector[77] +matrix[78][101] * vector[78] +matrix[79][101] * vector[79] +matrix[80][101] * vector[80] +matrix[81][101] * vector[81] +matrix[82][101] * vector[82] +matrix[83][101] * vector[83] +matrix[84][101] * vector[84] +matrix[85][101] * vector[85] +matrix[86][101] * vector[86] +matrix[87][101] * vector[87] +matrix[88][101] * vector[88] +matrix[89][101] * vector[89] +matrix[90][101] * vector[90] +matrix[91][101] * vector[91] +matrix[92][101] * vector[92] +matrix[93][101] * vector[93] +matrix[94][101] * vector[94] +matrix[95][101] * vector[95] +matrix[96][101] * vector[96] +matrix[97][101] * vector[97] +matrix[98][101] * vector[98] +matrix[99][101] * vector[99] +b[101];
assign result[102] = matrix[0][102] * vector[0] +matrix[1][102] * vector[1] +matrix[2][102] * vector[2] +matrix[3][102] * vector[3] +matrix[4][102] * vector[4] +matrix[5][102] * vector[5] +matrix[6][102] * vector[6] +matrix[7][102] * vector[7] +matrix[8][102] * vector[8] +matrix[9][102] * vector[9] +matrix[10][102] * vector[10] +matrix[11][102] * vector[11] +matrix[12][102] * vector[12] +matrix[13][102] * vector[13] +matrix[14][102] * vector[14] +matrix[15][102] * vector[15] +matrix[16][102] * vector[16] +matrix[17][102] * vector[17] +matrix[18][102] * vector[18] +matrix[19][102] * vector[19] +matrix[20][102] * vector[20] +matrix[21][102] * vector[21] +matrix[22][102] * vector[22] +matrix[23][102] * vector[23] +matrix[24][102] * vector[24] +matrix[25][102] * vector[25] +matrix[26][102] * vector[26] +matrix[27][102] * vector[27] +matrix[28][102] * vector[28] +matrix[29][102] * vector[29] +matrix[30][102] * vector[30] +matrix[31][102] * vector[31] +matrix[32][102] * vector[32] +matrix[33][102] * vector[33] +matrix[34][102] * vector[34] +matrix[35][102] * vector[35] +matrix[36][102] * vector[36] +matrix[37][102] * vector[37] +matrix[38][102] * vector[38] +matrix[39][102] * vector[39] +matrix[40][102] * vector[40] +matrix[41][102] * vector[41] +matrix[42][102] * vector[42] +matrix[43][102] * vector[43] +matrix[44][102] * vector[44] +matrix[45][102] * vector[45] +matrix[46][102] * vector[46] +matrix[47][102] * vector[47] +matrix[48][102] * vector[48] +matrix[49][102] * vector[49] +matrix[50][102] * vector[50] +matrix[51][102] * vector[51] +matrix[52][102] * vector[52] +matrix[53][102] * vector[53] +matrix[54][102] * vector[54] +matrix[55][102] * vector[55] +matrix[56][102] * vector[56] +matrix[57][102] * vector[57] +matrix[58][102] * vector[58] +matrix[59][102] * vector[59] +matrix[60][102] * vector[60] +matrix[61][102] * vector[61] +matrix[62][102] * vector[62] +matrix[63][102] * vector[63] +matrix[64][102] * vector[64] +matrix[65][102] * vector[65] +matrix[66][102] * vector[66] +matrix[67][102] * vector[67] +matrix[68][102] * vector[68] +matrix[69][102] * vector[69] +matrix[70][102] * vector[70] +matrix[71][102] * vector[71] +matrix[72][102] * vector[72] +matrix[73][102] * vector[73] +matrix[74][102] * vector[74] +matrix[75][102] * vector[75] +matrix[76][102] * vector[76] +matrix[77][102] * vector[77] +matrix[78][102] * vector[78] +matrix[79][102] * vector[79] +matrix[80][102] * vector[80] +matrix[81][102] * vector[81] +matrix[82][102] * vector[82] +matrix[83][102] * vector[83] +matrix[84][102] * vector[84] +matrix[85][102] * vector[85] +matrix[86][102] * vector[86] +matrix[87][102] * vector[87] +matrix[88][102] * vector[88] +matrix[89][102] * vector[89] +matrix[90][102] * vector[90] +matrix[91][102] * vector[91] +matrix[92][102] * vector[92] +matrix[93][102] * vector[93] +matrix[94][102] * vector[94] +matrix[95][102] * vector[95] +matrix[96][102] * vector[96] +matrix[97][102] * vector[97] +matrix[98][102] * vector[98] +matrix[99][102] * vector[99] +b[102];
assign result[103] = matrix[0][103] * vector[0] +matrix[1][103] * vector[1] +matrix[2][103] * vector[2] +matrix[3][103] * vector[3] +matrix[4][103] * vector[4] +matrix[5][103] * vector[5] +matrix[6][103] * vector[6] +matrix[7][103] * vector[7] +matrix[8][103] * vector[8] +matrix[9][103] * vector[9] +matrix[10][103] * vector[10] +matrix[11][103] * vector[11] +matrix[12][103] * vector[12] +matrix[13][103] * vector[13] +matrix[14][103] * vector[14] +matrix[15][103] * vector[15] +matrix[16][103] * vector[16] +matrix[17][103] * vector[17] +matrix[18][103] * vector[18] +matrix[19][103] * vector[19] +matrix[20][103] * vector[20] +matrix[21][103] * vector[21] +matrix[22][103] * vector[22] +matrix[23][103] * vector[23] +matrix[24][103] * vector[24] +matrix[25][103] * vector[25] +matrix[26][103] * vector[26] +matrix[27][103] * vector[27] +matrix[28][103] * vector[28] +matrix[29][103] * vector[29] +matrix[30][103] * vector[30] +matrix[31][103] * vector[31] +matrix[32][103] * vector[32] +matrix[33][103] * vector[33] +matrix[34][103] * vector[34] +matrix[35][103] * vector[35] +matrix[36][103] * vector[36] +matrix[37][103] * vector[37] +matrix[38][103] * vector[38] +matrix[39][103] * vector[39] +matrix[40][103] * vector[40] +matrix[41][103] * vector[41] +matrix[42][103] * vector[42] +matrix[43][103] * vector[43] +matrix[44][103] * vector[44] +matrix[45][103] * vector[45] +matrix[46][103] * vector[46] +matrix[47][103] * vector[47] +matrix[48][103] * vector[48] +matrix[49][103] * vector[49] +matrix[50][103] * vector[50] +matrix[51][103] * vector[51] +matrix[52][103] * vector[52] +matrix[53][103] * vector[53] +matrix[54][103] * vector[54] +matrix[55][103] * vector[55] +matrix[56][103] * vector[56] +matrix[57][103] * vector[57] +matrix[58][103] * vector[58] +matrix[59][103] * vector[59] +matrix[60][103] * vector[60] +matrix[61][103] * vector[61] +matrix[62][103] * vector[62] +matrix[63][103] * vector[63] +matrix[64][103] * vector[64] +matrix[65][103] * vector[65] +matrix[66][103] * vector[66] +matrix[67][103] * vector[67] +matrix[68][103] * vector[68] +matrix[69][103] * vector[69] +matrix[70][103] * vector[70] +matrix[71][103] * vector[71] +matrix[72][103] * vector[72] +matrix[73][103] * vector[73] +matrix[74][103] * vector[74] +matrix[75][103] * vector[75] +matrix[76][103] * vector[76] +matrix[77][103] * vector[77] +matrix[78][103] * vector[78] +matrix[79][103] * vector[79] +matrix[80][103] * vector[80] +matrix[81][103] * vector[81] +matrix[82][103] * vector[82] +matrix[83][103] * vector[83] +matrix[84][103] * vector[84] +matrix[85][103] * vector[85] +matrix[86][103] * vector[86] +matrix[87][103] * vector[87] +matrix[88][103] * vector[88] +matrix[89][103] * vector[89] +matrix[90][103] * vector[90] +matrix[91][103] * vector[91] +matrix[92][103] * vector[92] +matrix[93][103] * vector[93] +matrix[94][103] * vector[94] +matrix[95][103] * vector[95] +matrix[96][103] * vector[96] +matrix[97][103] * vector[97] +matrix[98][103] * vector[98] +matrix[99][103] * vector[99] +b[103];
assign result[104] = matrix[0][104] * vector[0] +matrix[1][104] * vector[1] +matrix[2][104] * vector[2] +matrix[3][104] * vector[3] +matrix[4][104] * vector[4] +matrix[5][104] * vector[5] +matrix[6][104] * vector[6] +matrix[7][104] * vector[7] +matrix[8][104] * vector[8] +matrix[9][104] * vector[9] +matrix[10][104] * vector[10] +matrix[11][104] * vector[11] +matrix[12][104] * vector[12] +matrix[13][104] * vector[13] +matrix[14][104] * vector[14] +matrix[15][104] * vector[15] +matrix[16][104] * vector[16] +matrix[17][104] * vector[17] +matrix[18][104] * vector[18] +matrix[19][104] * vector[19] +matrix[20][104] * vector[20] +matrix[21][104] * vector[21] +matrix[22][104] * vector[22] +matrix[23][104] * vector[23] +matrix[24][104] * vector[24] +matrix[25][104] * vector[25] +matrix[26][104] * vector[26] +matrix[27][104] * vector[27] +matrix[28][104] * vector[28] +matrix[29][104] * vector[29] +matrix[30][104] * vector[30] +matrix[31][104] * vector[31] +matrix[32][104] * vector[32] +matrix[33][104] * vector[33] +matrix[34][104] * vector[34] +matrix[35][104] * vector[35] +matrix[36][104] * vector[36] +matrix[37][104] * vector[37] +matrix[38][104] * vector[38] +matrix[39][104] * vector[39] +matrix[40][104] * vector[40] +matrix[41][104] * vector[41] +matrix[42][104] * vector[42] +matrix[43][104] * vector[43] +matrix[44][104] * vector[44] +matrix[45][104] * vector[45] +matrix[46][104] * vector[46] +matrix[47][104] * vector[47] +matrix[48][104] * vector[48] +matrix[49][104] * vector[49] +matrix[50][104] * vector[50] +matrix[51][104] * vector[51] +matrix[52][104] * vector[52] +matrix[53][104] * vector[53] +matrix[54][104] * vector[54] +matrix[55][104] * vector[55] +matrix[56][104] * vector[56] +matrix[57][104] * vector[57] +matrix[58][104] * vector[58] +matrix[59][104] * vector[59] +matrix[60][104] * vector[60] +matrix[61][104] * vector[61] +matrix[62][104] * vector[62] +matrix[63][104] * vector[63] +matrix[64][104] * vector[64] +matrix[65][104] * vector[65] +matrix[66][104] * vector[66] +matrix[67][104] * vector[67] +matrix[68][104] * vector[68] +matrix[69][104] * vector[69] +matrix[70][104] * vector[70] +matrix[71][104] * vector[71] +matrix[72][104] * vector[72] +matrix[73][104] * vector[73] +matrix[74][104] * vector[74] +matrix[75][104] * vector[75] +matrix[76][104] * vector[76] +matrix[77][104] * vector[77] +matrix[78][104] * vector[78] +matrix[79][104] * vector[79] +matrix[80][104] * vector[80] +matrix[81][104] * vector[81] +matrix[82][104] * vector[82] +matrix[83][104] * vector[83] +matrix[84][104] * vector[84] +matrix[85][104] * vector[85] +matrix[86][104] * vector[86] +matrix[87][104] * vector[87] +matrix[88][104] * vector[88] +matrix[89][104] * vector[89] +matrix[90][104] * vector[90] +matrix[91][104] * vector[91] +matrix[92][104] * vector[92] +matrix[93][104] * vector[93] +matrix[94][104] * vector[94] +matrix[95][104] * vector[95] +matrix[96][104] * vector[96] +matrix[97][104] * vector[97] +matrix[98][104] * vector[98] +matrix[99][104] * vector[99] +b[104];
assign result[105] = matrix[0][105] * vector[0] +matrix[1][105] * vector[1] +matrix[2][105] * vector[2] +matrix[3][105] * vector[3] +matrix[4][105] * vector[4] +matrix[5][105] * vector[5] +matrix[6][105] * vector[6] +matrix[7][105] * vector[7] +matrix[8][105] * vector[8] +matrix[9][105] * vector[9] +matrix[10][105] * vector[10] +matrix[11][105] * vector[11] +matrix[12][105] * vector[12] +matrix[13][105] * vector[13] +matrix[14][105] * vector[14] +matrix[15][105] * vector[15] +matrix[16][105] * vector[16] +matrix[17][105] * vector[17] +matrix[18][105] * vector[18] +matrix[19][105] * vector[19] +matrix[20][105] * vector[20] +matrix[21][105] * vector[21] +matrix[22][105] * vector[22] +matrix[23][105] * vector[23] +matrix[24][105] * vector[24] +matrix[25][105] * vector[25] +matrix[26][105] * vector[26] +matrix[27][105] * vector[27] +matrix[28][105] * vector[28] +matrix[29][105] * vector[29] +matrix[30][105] * vector[30] +matrix[31][105] * vector[31] +matrix[32][105] * vector[32] +matrix[33][105] * vector[33] +matrix[34][105] * vector[34] +matrix[35][105] * vector[35] +matrix[36][105] * vector[36] +matrix[37][105] * vector[37] +matrix[38][105] * vector[38] +matrix[39][105] * vector[39] +matrix[40][105] * vector[40] +matrix[41][105] * vector[41] +matrix[42][105] * vector[42] +matrix[43][105] * vector[43] +matrix[44][105] * vector[44] +matrix[45][105] * vector[45] +matrix[46][105] * vector[46] +matrix[47][105] * vector[47] +matrix[48][105] * vector[48] +matrix[49][105] * vector[49] +matrix[50][105] * vector[50] +matrix[51][105] * vector[51] +matrix[52][105] * vector[52] +matrix[53][105] * vector[53] +matrix[54][105] * vector[54] +matrix[55][105] * vector[55] +matrix[56][105] * vector[56] +matrix[57][105] * vector[57] +matrix[58][105] * vector[58] +matrix[59][105] * vector[59] +matrix[60][105] * vector[60] +matrix[61][105] * vector[61] +matrix[62][105] * vector[62] +matrix[63][105] * vector[63] +matrix[64][105] * vector[64] +matrix[65][105] * vector[65] +matrix[66][105] * vector[66] +matrix[67][105] * vector[67] +matrix[68][105] * vector[68] +matrix[69][105] * vector[69] +matrix[70][105] * vector[70] +matrix[71][105] * vector[71] +matrix[72][105] * vector[72] +matrix[73][105] * vector[73] +matrix[74][105] * vector[74] +matrix[75][105] * vector[75] +matrix[76][105] * vector[76] +matrix[77][105] * vector[77] +matrix[78][105] * vector[78] +matrix[79][105] * vector[79] +matrix[80][105] * vector[80] +matrix[81][105] * vector[81] +matrix[82][105] * vector[82] +matrix[83][105] * vector[83] +matrix[84][105] * vector[84] +matrix[85][105] * vector[85] +matrix[86][105] * vector[86] +matrix[87][105] * vector[87] +matrix[88][105] * vector[88] +matrix[89][105] * vector[89] +matrix[90][105] * vector[90] +matrix[91][105] * vector[91] +matrix[92][105] * vector[92] +matrix[93][105] * vector[93] +matrix[94][105] * vector[94] +matrix[95][105] * vector[95] +matrix[96][105] * vector[96] +matrix[97][105] * vector[97] +matrix[98][105] * vector[98] +matrix[99][105] * vector[99] +b[105];
assign result[106] = matrix[0][106] * vector[0] +matrix[1][106] * vector[1] +matrix[2][106] * vector[2] +matrix[3][106] * vector[3] +matrix[4][106] * vector[4] +matrix[5][106] * vector[5] +matrix[6][106] * vector[6] +matrix[7][106] * vector[7] +matrix[8][106] * vector[8] +matrix[9][106] * vector[9] +matrix[10][106] * vector[10] +matrix[11][106] * vector[11] +matrix[12][106] * vector[12] +matrix[13][106] * vector[13] +matrix[14][106] * vector[14] +matrix[15][106] * vector[15] +matrix[16][106] * vector[16] +matrix[17][106] * vector[17] +matrix[18][106] * vector[18] +matrix[19][106] * vector[19] +matrix[20][106] * vector[20] +matrix[21][106] * vector[21] +matrix[22][106] * vector[22] +matrix[23][106] * vector[23] +matrix[24][106] * vector[24] +matrix[25][106] * vector[25] +matrix[26][106] * vector[26] +matrix[27][106] * vector[27] +matrix[28][106] * vector[28] +matrix[29][106] * vector[29] +matrix[30][106] * vector[30] +matrix[31][106] * vector[31] +matrix[32][106] * vector[32] +matrix[33][106] * vector[33] +matrix[34][106] * vector[34] +matrix[35][106] * vector[35] +matrix[36][106] * vector[36] +matrix[37][106] * vector[37] +matrix[38][106] * vector[38] +matrix[39][106] * vector[39] +matrix[40][106] * vector[40] +matrix[41][106] * vector[41] +matrix[42][106] * vector[42] +matrix[43][106] * vector[43] +matrix[44][106] * vector[44] +matrix[45][106] * vector[45] +matrix[46][106] * vector[46] +matrix[47][106] * vector[47] +matrix[48][106] * vector[48] +matrix[49][106] * vector[49] +matrix[50][106] * vector[50] +matrix[51][106] * vector[51] +matrix[52][106] * vector[52] +matrix[53][106] * vector[53] +matrix[54][106] * vector[54] +matrix[55][106] * vector[55] +matrix[56][106] * vector[56] +matrix[57][106] * vector[57] +matrix[58][106] * vector[58] +matrix[59][106] * vector[59] +matrix[60][106] * vector[60] +matrix[61][106] * vector[61] +matrix[62][106] * vector[62] +matrix[63][106] * vector[63] +matrix[64][106] * vector[64] +matrix[65][106] * vector[65] +matrix[66][106] * vector[66] +matrix[67][106] * vector[67] +matrix[68][106] * vector[68] +matrix[69][106] * vector[69] +matrix[70][106] * vector[70] +matrix[71][106] * vector[71] +matrix[72][106] * vector[72] +matrix[73][106] * vector[73] +matrix[74][106] * vector[74] +matrix[75][106] * vector[75] +matrix[76][106] * vector[76] +matrix[77][106] * vector[77] +matrix[78][106] * vector[78] +matrix[79][106] * vector[79] +matrix[80][106] * vector[80] +matrix[81][106] * vector[81] +matrix[82][106] * vector[82] +matrix[83][106] * vector[83] +matrix[84][106] * vector[84] +matrix[85][106] * vector[85] +matrix[86][106] * vector[86] +matrix[87][106] * vector[87] +matrix[88][106] * vector[88] +matrix[89][106] * vector[89] +matrix[90][106] * vector[90] +matrix[91][106] * vector[91] +matrix[92][106] * vector[92] +matrix[93][106] * vector[93] +matrix[94][106] * vector[94] +matrix[95][106] * vector[95] +matrix[96][106] * vector[96] +matrix[97][106] * vector[97] +matrix[98][106] * vector[98] +matrix[99][106] * vector[99] +b[106];
assign result[107] = matrix[0][107] * vector[0] +matrix[1][107] * vector[1] +matrix[2][107] * vector[2] +matrix[3][107] * vector[3] +matrix[4][107] * vector[4] +matrix[5][107] * vector[5] +matrix[6][107] * vector[6] +matrix[7][107] * vector[7] +matrix[8][107] * vector[8] +matrix[9][107] * vector[9] +matrix[10][107] * vector[10] +matrix[11][107] * vector[11] +matrix[12][107] * vector[12] +matrix[13][107] * vector[13] +matrix[14][107] * vector[14] +matrix[15][107] * vector[15] +matrix[16][107] * vector[16] +matrix[17][107] * vector[17] +matrix[18][107] * vector[18] +matrix[19][107] * vector[19] +matrix[20][107] * vector[20] +matrix[21][107] * vector[21] +matrix[22][107] * vector[22] +matrix[23][107] * vector[23] +matrix[24][107] * vector[24] +matrix[25][107] * vector[25] +matrix[26][107] * vector[26] +matrix[27][107] * vector[27] +matrix[28][107] * vector[28] +matrix[29][107] * vector[29] +matrix[30][107] * vector[30] +matrix[31][107] * vector[31] +matrix[32][107] * vector[32] +matrix[33][107] * vector[33] +matrix[34][107] * vector[34] +matrix[35][107] * vector[35] +matrix[36][107] * vector[36] +matrix[37][107] * vector[37] +matrix[38][107] * vector[38] +matrix[39][107] * vector[39] +matrix[40][107] * vector[40] +matrix[41][107] * vector[41] +matrix[42][107] * vector[42] +matrix[43][107] * vector[43] +matrix[44][107] * vector[44] +matrix[45][107] * vector[45] +matrix[46][107] * vector[46] +matrix[47][107] * vector[47] +matrix[48][107] * vector[48] +matrix[49][107] * vector[49] +matrix[50][107] * vector[50] +matrix[51][107] * vector[51] +matrix[52][107] * vector[52] +matrix[53][107] * vector[53] +matrix[54][107] * vector[54] +matrix[55][107] * vector[55] +matrix[56][107] * vector[56] +matrix[57][107] * vector[57] +matrix[58][107] * vector[58] +matrix[59][107] * vector[59] +matrix[60][107] * vector[60] +matrix[61][107] * vector[61] +matrix[62][107] * vector[62] +matrix[63][107] * vector[63] +matrix[64][107] * vector[64] +matrix[65][107] * vector[65] +matrix[66][107] * vector[66] +matrix[67][107] * vector[67] +matrix[68][107] * vector[68] +matrix[69][107] * vector[69] +matrix[70][107] * vector[70] +matrix[71][107] * vector[71] +matrix[72][107] * vector[72] +matrix[73][107] * vector[73] +matrix[74][107] * vector[74] +matrix[75][107] * vector[75] +matrix[76][107] * vector[76] +matrix[77][107] * vector[77] +matrix[78][107] * vector[78] +matrix[79][107] * vector[79] +matrix[80][107] * vector[80] +matrix[81][107] * vector[81] +matrix[82][107] * vector[82] +matrix[83][107] * vector[83] +matrix[84][107] * vector[84] +matrix[85][107] * vector[85] +matrix[86][107] * vector[86] +matrix[87][107] * vector[87] +matrix[88][107] * vector[88] +matrix[89][107] * vector[89] +matrix[90][107] * vector[90] +matrix[91][107] * vector[91] +matrix[92][107] * vector[92] +matrix[93][107] * vector[93] +matrix[94][107] * vector[94] +matrix[95][107] * vector[95] +matrix[96][107] * vector[96] +matrix[97][107] * vector[97] +matrix[98][107] * vector[98] +matrix[99][107] * vector[99] +b[107];
assign result[108] = matrix[0][108] * vector[0] +matrix[1][108] * vector[1] +matrix[2][108] * vector[2] +matrix[3][108] * vector[3] +matrix[4][108] * vector[4] +matrix[5][108] * vector[5] +matrix[6][108] * vector[6] +matrix[7][108] * vector[7] +matrix[8][108] * vector[8] +matrix[9][108] * vector[9] +matrix[10][108] * vector[10] +matrix[11][108] * vector[11] +matrix[12][108] * vector[12] +matrix[13][108] * vector[13] +matrix[14][108] * vector[14] +matrix[15][108] * vector[15] +matrix[16][108] * vector[16] +matrix[17][108] * vector[17] +matrix[18][108] * vector[18] +matrix[19][108] * vector[19] +matrix[20][108] * vector[20] +matrix[21][108] * vector[21] +matrix[22][108] * vector[22] +matrix[23][108] * vector[23] +matrix[24][108] * vector[24] +matrix[25][108] * vector[25] +matrix[26][108] * vector[26] +matrix[27][108] * vector[27] +matrix[28][108] * vector[28] +matrix[29][108] * vector[29] +matrix[30][108] * vector[30] +matrix[31][108] * vector[31] +matrix[32][108] * vector[32] +matrix[33][108] * vector[33] +matrix[34][108] * vector[34] +matrix[35][108] * vector[35] +matrix[36][108] * vector[36] +matrix[37][108] * vector[37] +matrix[38][108] * vector[38] +matrix[39][108] * vector[39] +matrix[40][108] * vector[40] +matrix[41][108] * vector[41] +matrix[42][108] * vector[42] +matrix[43][108] * vector[43] +matrix[44][108] * vector[44] +matrix[45][108] * vector[45] +matrix[46][108] * vector[46] +matrix[47][108] * vector[47] +matrix[48][108] * vector[48] +matrix[49][108] * vector[49] +matrix[50][108] * vector[50] +matrix[51][108] * vector[51] +matrix[52][108] * vector[52] +matrix[53][108] * vector[53] +matrix[54][108] * vector[54] +matrix[55][108] * vector[55] +matrix[56][108] * vector[56] +matrix[57][108] * vector[57] +matrix[58][108] * vector[58] +matrix[59][108] * vector[59] +matrix[60][108] * vector[60] +matrix[61][108] * vector[61] +matrix[62][108] * vector[62] +matrix[63][108] * vector[63] +matrix[64][108] * vector[64] +matrix[65][108] * vector[65] +matrix[66][108] * vector[66] +matrix[67][108] * vector[67] +matrix[68][108] * vector[68] +matrix[69][108] * vector[69] +matrix[70][108] * vector[70] +matrix[71][108] * vector[71] +matrix[72][108] * vector[72] +matrix[73][108] * vector[73] +matrix[74][108] * vector[74] +matrix[75][108] * vector[75] +matrix[76][108] * vector[76] +matrix[77][108] * vector[77] +matrix[78][108] * vector[78] +matrix[79][108] * vector[79] +matrix[80][108] * vector[80] +matrix[81][108] * vector[81] +matrix[82][108] * vector[82] +matrix[83][108] * vector[83] +matrix[84][108] * vector[84] +matrix[85][108] * vector[85] +matrix[86][108] * vector[86] +matrix[87][108] * vector[87] +matrix[88][108] * vector[88] +matrix[89][108] * vector[89] +matrix[90][108] * vector[90] +matrix[91][108] * vector[91] +matrix[92][108] * vector[92] +matrix[93][108] * vector[93] +matrix[94][108] * vector[94] +matrix[95][108] * vector[95] +matrix[96][108] * vector[96] +matrix[97][108] * vector[97] +matrix[98][108] * vector[98] +matrix[99][108] * vector[99] +b[108];
assign result[109] = matrix[0][109] * vector[0] +matrix[1][109] * vector[1] +matrix[2][109] * vector[2] +matrix[3][109] * vector[3] +matrix[4][109] * vector[4] +matrix[5][109] * vector[5] +matrix[6][109] * vector[6] +matrix[7][109] * vector[7] +matrix[8][109] * vector[8] +matrix[9][109] * vector[9] +matrix[10][109] * vector[10] +matrix[11][109] * vector[11] +matrix[12][109] * vector[12] +matrix[13][109] * vector[13] +matrix[14][109] * vector[14] +matrix[15][109] * vector[15] +matrix[16][109] * vector[16] +matrix[17][109] * vector[17] +matrix[18][109] * vector[18] +matrix[19][109] * vector[19] +matrix[20][109] * vector[20] +matrix[21][109] * vector[21] +matrix[22][109] * vector[22] +matrix[23][109] * vector[23] +matrix[24][109] * vector[24] +matrix[25][109] * vector[25] +matrix[26][109] * vector[26] +matrix[27][109] * vector[27] +matrix[28][109] * vector[28] +matrix[29][109] * vector[29] +matrix[30][109] * vector[30] +matrix[31][109] * vector[31] +matrix[32][109] * vector[32] +matrix[33][109] * vector[33] +matrix[34][109] * vector[34] +matrix[35][109] * vector[35] +matrix[36][109] * vector[36] +matrix[37][109] * vector[37] +matrix[38][109] * vector[38] +matrix[39][109] * vector[39] +matrix[40][109] * vector[40] +matrix[41][109] * vector[41] +matrix[42][109] * vector[42] +matrix[43][109] * vector[43] +matrix[44][109] * vector[44] +matrix[45][109] * vector[45] +matrix[46][109] * vector[46] +matrix[47][109] * vector[47] +matrix[48][109] * vector[48] +matrix[49][109] * vector[49] +matrix[50][109] * vector[50] +matrix[51][109] * vector[51] +matrix[52][109] * vector[52] +matrix[53][109] * vector[53] +matrix[54][109] * vector[54] +matrix[55][109] * vector[55] +matrix[56][109] * vector[56] +matrix[57][109] * vector[57] +matrix[58][109] * vector[58] +matrix[59][109] * vector[59] +matrix[60][109] * vector[60] +matrix[61][109] * vector[61] +matrix[62][109] * vector[62] +matrix[63][109] * vector[63] +matrix[64][109] * vector[64] +matrix[65][109] * vector[65] +matrix[66][109] * vector[66] +matrix[67][109] * vector[67] +matrix[68][109] * vector[68] +matrix[69][109] * vector[69] +matrix[70][109] * vector[70] +matrix[71][109] * vector[71] +matrix[72][109] * vector[72] +matrix[73][109] * vector[73] +matrix[74][109] * vector[74] +matrix[75][109] * vector[75] +matrix[76][109] * vector[76] +matrix[77][109] * vector[77] +matrix[78][109] * vector[78] +matrix[79][109] * vector[79] +matrix[80][109] * vector[80] +matrix[81][109] * vector[81] +matrix[82][109] * vector[82] +matrix[83][109] * vector[83] +matrix[84][109] * vector[84] +matrix[85][109] * vector[85] +matrix[86][109] * vector[86] +matrix[87][109] * vector[87] +matrix[88][109] * vector[88] +matrix[89][109] * vector[89] +matrix[90][109] * vector[90] +matrix[91][109] * vector[91] +matrix[92][109] * vector[92] +matrix[93][109] * vector[93] +matrix[94][109] * vector[94] +matrix[95][109] * vector[95] +matrix[96][109] * vector[96] +matrix[97][109] * vector[97] +matrix[98][109] * vector[98] +matrix[99][109] * vector[99] +b[109];
assign result[110] = matrix[0][110] * vector[0] +matrix[1][110] * vector[1] +matrix[2][110] * vector[2] +matrix[3][110] * vector[3] +matrix[4][110] * vector[4] +matrix[5][110] * vector[5] +matrix[6][110] * vector[6] +matrix[7][110] * vector[7] +matrix[8][110] * vector[8] +matrix[9][110] * vector[9] +matrix[10][110] * vector[10] +matrix[11][110] * vector[11] +matrix[12][110] * vector[12] +matrix[13][110] * vector[13] +matrix[14][110] * vector[14] +matrix[15][110] * vector[15] +matrix[16][110] * vector[16] +matrix[17][110] * vector[17] +matrix[18][110] * vector[18] +matrix[19][110] * vector[19] +matrix[20][110] * vector[20] +matrix[21][110] * vector[21] +matrix[22][110] * vector[22] +matrix[23][110] * vector[23] +matrix[24][110] * vector[24] +matrix[25][110] * vector[25] +matrix[26][110] * vector[26] +matrix[27][110] * vector[27] +matrix[28][110] * vector[28] +matrix[29][110] * vector[29] +matrix[30][110] * vector[30] +matrix[31][110] * vector[31] +matrix[32][110] * vector[32] +matrix[33][110] * vector[33] +matrix[34][110] * vector[34] +matrix[35][110] * vector[35] +matrix[36][110] * vector[36] +matrix[37][110] * vector[37] +matrix[38][110] * vector[38] +matrix[39][110] * vector[39] +matrix[40][110] * vector[40] +matrix[41][110] * vector[41] +matrix[42][110] * vector[42] +matrix[43][110] * vector[43] +matrix[44][110] * vector[44] +matrix[45][110] * vector[45] +matrix[46][110] * vector[46] +matrix[47][110] * vector[47] +matrix[48][110] * vector[48] +matrix[49][110] * vector[49] +matrix[50][110] * vector[50] +matrix[51][110] * vector[51] +matrix[52][110] * vector[52] +matrix[53][110] * vector[53] +matrix[54][110] * vector[54] +matrix[55][110] * vector[55] +matrix[56][110] * vector[56] +matrix[57][110] * vector[57] +matrix[58][110] * vector[58] +matrix[59][110] * vector[59] +matrix[60][110] * vector[60] +matrix[61][110] * vector[61] +matrix[62][110] * vector[62] +matrix[63][110] * vector[63] +matrix[64][110] * vector[64] +matrix[65][110] * vector[65] +matrix[66][110] * vector[66] +matrix[67][110] * vector[67] +matrix[68][110] * vector[68] +matrix[69][110] * vector[69] +matrix[70][110] * vector[70] +matrix[71][110] * vector[71] +matrix[72][110] * vector[72] +matrix[73][110] * vector[73] +matrix[74][110] * vector[74] +matrix[75][110] * vector[75] +matrix[76][110] * vector[76] +matrix[77][110] * vector[77] +matrix[78][110] * vector[78] +matrix[79][110] * vector[79] +matrix[80][110] * vector[80] +matrix[81][110] * vector[81] +matrix[82][110] * vector[82] +matrix[83][110] * vector[83] +matrix[84][110] * vector[84] +matrix[85][110] * vector[85] +matrix[86][110] * vector[86] +matrix[87][110] * vector[87] +matrix[88][110] * vector[88] +matrix[89][110] * vector[89] +matrix[90][110] * vector[90] +matrix[91][110] * vector[91] +matrix[92][110] * vector[92] +matrix[93][110] * vector[93] +matrix[94][110] * vector[94] +matrix[95][110] * vector[95] +matrix[96][110] * vector[96] +matrix[97][110] * vector[97] +matrix[98][110] * vector[98] +matrix[99][110] * vector[99] +b[110];
assign result[111] = matrix[0][111] * vector[0] +matrix[1][111] * vector[1] +matrix[2][111] * vector[2] +matrix[3][111] * vector[3] +matrix[4][111] * vector[4] +matrix[5][111] * vector[5] +matrix[6][111] * vector[6] +matrix[7][111] * vector[7] +matrix[8][111] * vector[8] +matrix[9][111] * vector[9] +matrix[10][111] * vector[10] +matrix[11][111] * vector[11] +matrix[12][111] * vector[12] +matrix[13][111] * vector[13] +matrix[14][111] * vector[14] +matrix[15][111] * vector[15] +matrix[16][111] * vector[16] +matrix[17][111] * vector[17] +matrix[18][111] * vector[18] +matrix[19][111] * vector[19] +matrix[20][111] * vector[20] +matrix[21][111] * vector[21] +matrix[22][111] * vector[22] +matrix[23][111] * vector[23] +matrix[24][111] * vector[24] +matrix[25][111] * vector[25] +matrix[26][111] * vector[26] +matrix[27][111] * vector[27] +matrix[28][111] * vector[28] +matrix[29][111] * vector[29] +matrix[30][111] * vector[30] +matrix[31][111] * vector[31] +matrix[32][111] * vector[32] +matrix[33][111] * vector[33] +matrix[34][111] * vector[34] +matrix[35][111] * vector[35] +matrix[36][111] * vector[36] +matrix[37][111] * vector[37] +matrix[38][111] * vector[38] +matrix[39][111] * vector[39] +matrix[40][111] * vector[40] +matrix[41][111] * vector[41] +matrix[42][111] * vector[42] +matrix[43][111] * vector[43] +matrix[44][111] * vector[44] +matrix[45][111] * vector[45] +matrix[46][111] * vector[46] +matrix[47][111] * vector[47] +matrix[48][111] * vector[48] +matrix[49][111] * vector[49] +matrix[50][111] * vector[50] +matrix[51][111] * vector[51] +matrix[52][111] * vector[52] +matrix[53][111] * vector[53] +matrix[54][111] * vector[54] +matrix[55][111] * vector[55] +matrix[56][111] * vector[56] +matrix[57][111] * vector[57] +matrix[58][111] * vector[58] +matrix[59][111] * vector[59] +matrix[60][111] * vector[60] +matrix[61][111] * vector[61] +matrix[62][111] * vector[62] +matrix[63][111] * vector[63] +matrix[64][111] * vector[64] +matrix[65][111] * vector[65] +matrix[66][111] * vector[66] +matrix[67][111] * vector[67] +matrix[68][111] * vector[68] +matrix[69][111] * vector[69] +matrix[70][111] * vector[70] +matrix[71][111] * vector[71] +matrix[72][111] * vector[72] +matrix[73][111] * vector[73] +matrix[74][111] * vector[74] +matrix[75][111] * vector[75] +matrix[76][111] * vector[76] +matrix[77][111] * vector[77] +matrix[78][111] * vector[78] +matrix[79][111] * vector[79] +matrix[80][111] * vector[80] +matrix[81][111] * vector[81] +matrix[82][111] * vector[82] +matrix[83][111] * vector[83] +matrix[84][111] * vector[84] +matrix[85][111] * vector[85] +matrix[86][111] * vector[86] +matrix[87][111] * vector[87] +matrix[88][111] * vector[88] +matrix[89][111] * vector[89] +matrix[90][111] * vector[90] +matrix[91][111] * vector[91] +matrix[92][111] * vector[92] +matrix[93][111] * vector[93] +matrix[94][111] * vector[94] +matrix[95][111] * vector[95] +matrix[96][111] * vector[96] +matrix[97][111] * vector[97] +matrix[98][111] * vector[98] +matrix[99][111] * vector[99] +b[111];
assign result[112] = matrix[0][112] * vector[0] +matrix[1][112] * vector[1] +matrix[2][112] * vector[2] +matrix[3][112] * vector[3] +matrix[4][112] * vector[4] +matrix[5][112] * vector[5] +matrix[6][112] * vector[6] +matrix[7][112] * vector[7] +matrix[8][112] * vector[8] +matrix[9][112] * vector[9] +matrix[10][112] * vector[10] +matrix[11][112] * vector[11] +matrix[12][112] * vector[12] +matrix[13][112] * vector[13] +matrix[14][112] * vector[14] +matrix[15][112] * vector[15] +matrix[16][112] * vector[16] +matrix[17][112] * vector[17] +matrix[18][112] * vector[18] +matrix[19][112] * vector[19] +matrix[20][112] * vector[20] +matrix[21][112] * vector[21] +matrix[22][112] * vector[22] +matrix[23][112] * vector[23] +matrix[24][112] * vector[24] +matrix[25][112] * vector[25] +matrix[26][112] * vector[26] +matrix[27][112] * vector[27] +matrix[28][112] * vector[28] +matrix[29][112] * vector[29] +matrix[30][112] * vector[30] +matrix[31][112] * vector[31] +matrix[32][112] * vector[32] +matrix[33][112] * vector[33] +matrix[34][112] * vector[34] +matrix[35][112] * vector[35] +matrix[36][112] * vector[36] +matrix[37][112] * vector[37] +matrix[38][112] * vector[38] +matrix[39][112] * vector[39] +matrix[40][112] * vector[40] +matrix[41][112] * vector[41] +matrix[42][112] * vector[42] +matrix[43][112] * vector[43] +matrix[44][112] * vector[44] +matrix[45][112] * vector[45] +matrix[46][112] * vector[46] +matrix[47][112] * vector[47] +matrix[48][112] * vector[48] +matrix[49][112] * vector[49] +matrix[50][112] * vector[50] +matrix[51][112] * vector[51] +matrix[52][112] * vector[52] +matrix[53][112] * vector[53] +matrix[54][112] * vector[54] +matrix[55][112] * vector[55] +matrix[56][112] * vector[56] +matrix[57][112] * vector[57] +matrix[58][112] * vector[58] +matrix[59][112] * vector[59] +matrix[60][112] * vector[60] +matrix[61][112] * vector[61] +matrix[62][112] * vector[62] +matrix[63][112] * vector[63] +matrix[64][112] * vector[64] +matrix[65][112] * vector[65] +matrix[66][112] * vector[66] +matrix[67][112] * vector[67] +matrix[68][112] * vector[68] +matrix[69][112] * vector[69] +matrix[70][112] * vector[70] +matrix[71][112] * vector[71] +matrix[72][112] * vector[72] +matrix[73][112] * vector[73] +matrix[74][112] * vector[74] +matrix[75][112] * vector[75] +matrix[76][112] * vector[76] +matrix[77][112] * vector[77] +matrix[78][112] * vector[78] +matrix[79][112] * vector[79] +matrix[80][112] * vector[80] +matrix[81][112] * vector[81] +matrix[82][112] * vector[82] +matrix[83][112] * vector[83] +matrix[84][112] * vector[84] +matrix[85][112] * vector[85] +matrix[86][112] * vector[86] +matrix[87][112] * vector[87] +matrix[88][112] * vector[88] +matrix[89][112] * vector[89] +matrix[90][112] * vector[90] +matrix[91][112] * vector[91] +matrix[92][112] * vector[92] +matrix[93][112] * vector[93] +matrix[94][112] * vector[94] +matrix[95][112] * vector[95] +matrix[96][112] * vector[96] +matrix[97][112] * vector[97] +matrix[98][112] * vector[98] +matrix[99][112] * vector[99] +b[112];
assign result[113] = matrix[0][113] * vector[0] +matrix[1][113] * vector[1] +matrix[2][113] * vector[2] +matrix[3][113] * vector[3] +matrix[4][113] * vector[4] +matrix[5][113] * vector[5] +matrix[6][113] * vector[6] +matrix[7][113] * vector[7] +matrix[8][113] * vector[8] +matrix[9][113] * vector[9] +matrix[10][113] * vector[10] +matrix[11][113] * vector[11] +matrix[12][113] * vector[12] +matrix[13][113] * vector[13] +matrix[14][113] * vector[14] +matrix[15][113] * vector[15] +matrix[16][113] * vector[16] +matrix[17][113] * vector[17] +matrix[18][113] * vector[18] +matrix[19][113] * vector[19] +matrix[20][113] * vector[20] +matrix[21][113] * vector[21] +matrix[22][113] * vector[22] +matrix[23][113] * vector[23] +matrix[24][113] * vector[24] +matrix[25][113] * vector[25] +matrix[26][113] * vector[26] +matrix[27][113] * vector[27] +matrix[28][113] * vector[28] +matrix[29][113] * vector[29] +matrix[30][113] * vector[30] +matrix[31][113] * vector[31] +matrix[32][113] * vector[32] +matrix[33][113] * vector[33] +matrix[34][113] * vector[34] +matrix[35][113] * vector[35] +matrix[36][113] * vector[36] +matrix[37][113] * vector[37] +matrix[38][113] * vector[38] +matrix[39][113] * vector[39] +matrix[40][113] * vector[40] +matrix[41][113] * vector[41] +matrix[42][113] * vector[42] +matrix[43][113] * vector[43] +matrix[44][113] * vector[44] +matrix[45][113] * vector[45] +matrix[46][113] * vector[46] +matrix[47][113] * vector[47] +matrix[48][113] * vector[48] +matrix[49][113] * vector[49] +matrix[50][113] * vector[50] +matrix[51][113] * vector[51] +matrix[52][113] * vector[52] +matrix[53][113] * vector[53] +matrix[54][113] * vector[54] +matrix[55][113] * vector[55] +matrix[56][113] * vector[56] +matrix[57][113] * vector[57] +matrix[58][113] * vector[58] +matrix[59][113] * vector[59] +matrix[60][113] * vector[60] +matrix[61][113] * vector[61] +matrix[62][113] * vector[62] +matrix[63][113] * vector[63] +matrix[64][113] * vector[64] +matrix[65][113] * vector[65] +matrix[66][113] * vector[66] +matrix[67][113] * vector[67] +matrix[68][113] * vector[68] +matrix[69][113] * vector[69] +matrix[70][113] * vector[70] +matrix[71][113] * vector[71] +matrix[72][113] * vector[72] +matrix[73][113] * vector[73] +matrix[74][113] * vector[74] +matrix[75][113] * vector[75] +matrix[76][113] * vector[76] +matrix[77][113] * vector[77] +matrix[78][113] * vector[78] +matrix[79][113] * vector[79] +matrix[80][113] * vector[80] +matrix[81][113] * vector[81] +matrix[82][113] * vector[82] +matrix[83][113] * vector[83] +matrix[84][113] * vector[84] +matrix[85][113] * vector[85] +matrix[86][113] * vector[86] +matrix[87][113] * vector[87] +matrix[88][113] * vector[88] +matrix[89][113] * vector[89] +matrix[90][113] * vector[90] +matrix[91][113] * vector[91] +matrix[92][113] * vector[92] +matrix[93][113] * vector[93] +matrix[94][113] * vector[94] +matrix[95][113] * vector[95] +matrix[96][113] * vector[96] +matrix[97][113] * vector[97] +matrix[98][113] * vector[98] +matrix[99][113] * vector[99] +b[113];
assign result[114] = matrix[0][114] * vector[0] +matrix[1][114] * vector[1] +matrix[2][114] * vector[2] +matrix[3][114] * vector[3] +matrix[4][114] * vector[4] +matrix[5][114] * vector[5] +matrix[6][114] * vector[6] +matrix[7][114] * vector[7] +matrix[8][114] * vector[8] +matrix[9][114] * vector[9] +matrix[10][114] * vector[10] +matrix[11][114] * vector[11] +matrix[12][114] * vector[12] +matrix[13][114] * vector[13] +matrix[14][114] * vector[14] +matrix[15][114] * vector[15] +matrix[16][114] * vector[16] +matrix[17][114] * vector[17] +matrix[18][114] * vector[18] +matrix[19][114] * vector[19] +matrix[20][114] * vector[20] +matrix[21][114] * vector[21] +matrix[22][114] * vector[22] +matrix[23][114] * vector[23] +matrix[24][114] * vector[24] +matrix[25][114] * vector[25] +matrix[26][114] * vector[26] +matrix[27][114] * vector[27] +matrix[28][114] * vector[28] +matrix[29][114] * vector[29] +matrix[30][114] * vector[30] +matrix[31][114] * vector[31] +matrix[32][114] * vector[32] +matrix[33][114] * vector[33] +matrix[34][114] * vector[34] +matrix[35][114] * vector[35] +matrix[36][114] * vector[36] +matrix[37][114] * vector[37] +matrix[38][114] * vector[38] +matrix[39][114] * vector[39] +matrix[40][114] * vector[40] +matrix[41][114] * vector[41] +matrix[42][114] * vector[42] +matrix[43][114] * vector[43] +matrix[44][114] * vector[44] +matrix[45][114] * vector[45] +matrix[46][114] * vector[46] +matrix[47][114] * vector[47] +matrix[48][114] * vector[48] +matrix[49][114] * vector[49] +matrix[50][114] * vector[50] +matrix[51][114] * vector[51] +matrix[52][114] * vector[52] +matrix[53][114] * vector[53] +matrix[54][114] * vector[54] +matrix[55][114] * vector[55] +matrix[56][114] * vector[56] +matrix[57][114] * vector[57] +matrix[58][114] * vector[58] +matrix[59][114] * vector[59] +matrix[60][114] * vector[60] +matrix[61][114] * vector[61] +matrix[62][114] * vector[62] +matrix[63][114] * vector[63] +matrix[64][114] * vector[64] +matrix[65][114] * vector[65] +matrix[66][114] * vector[66] +matrix[67][114] * vector[67] +matrix[68][114] * vector[68] +matrix[69][114] * vector[69] +matrix[70][114] * vector[70] +matrix[71][114] * vector[71] +matrix[72][114] * vector[72] +matrix[73][114] * vector[73] +matrix[74][114] * vector[74] +matrix[75][114] * vector[75] +matrix[76][114] * vector[76] +matrix[77][114] * vector[77] +matrix[78][114] * vector[78] +matrix[79][114] * vector[79] +matrix[80][114] * vector[80] +matrix[81][114] * vector[81] +matrix[82][114] * vector[82] +matrix[83][114] * vector[83] +matrix[84][114] * vector[84] +matrix[85][114] * vector[85] +matrix[86][114] * vector[86] +matrix[87][114] * vector[87] +matrix[88][114] * vector[88] +matrix[89][114] * vector[89] +matrix[90][114] * vector[90] +matrix[91][114] * vector[91] +matrix[92][114] * vector[92] +matrix[93][114] * vector[93] +matrix[94][114] * vector[94] +matrix[95][114] * vector[95] +matrix[96][114] * vector[96] +matrix[97][114] * vector[97] +matrix[98][114] * vector[98] +matrix[99][114] * vector[99] +b[114];
assign result[115] = matrix[0][115] * vector[0] +matrix[1][115] * vector[1] +matrix[2][115] * vector[2] +matrix[3][115] * vector[3] +matrix[4][115] * vector[4] +matrix[5][115] * vector[5] +matrix[6][115] * vector[6] +matrix[7][115] * vector[7] +matrix[8][115] * vector[8] +matrix[9][115] * vector[9] +matrix[10][115] * vector[10] +matrix[11][115] * vector[11] +matrix[12][115] * vector[12] +matrix[13][115] * vector[13] +matrix[14][115] * vector[14] +matrix[15][115] * vector[15] +matrix[16][115] * vector[16] +matrix[17][115] * vector[17] +matrix[18][115] * vector[18] +matrix[19][115] * vector[19] +matrix[20][115] * vector[20] +matrix[21][115] * vector[21] +matrix[22][115] * vector[22] +matrix[23][115] * vector[23] +matrix[24][115] * vector[24] +matrix[25][115] * vector[25] +matrix[26][115] * vector[26] +matrix[27][115] * vector[27] +matrix[28][115] * vector[28] +matrix[29][115] * vector[29] +matrix[30][115] * vector[30] +matrix[31][115] * vector[31] +matrix[32][115] * vector[32] +matrix[33][115] * vector[33] +matrix[34][115] * vector[34] +matrix[35][115] * vector[35] +matrix[36][115] * vector[36] +matrix[37][115] * vector[37] +matrix[38][115] * vector[38] +matrix[39][115] * vector[39] +matrix[40][115] * vector[40] +matrix[41][115] * vector[41] +matrix[42][115] * vector[42] +matrix[43][115] * vector[43] +matrix[44][115] * vector[44] +matrix[45][115] * vector[45] +matrix[46][115] * vector[46] +matrix[47][115] * vector[47] +matrix[48][115] * vector[48] +matrix[49][115] * vector[49] +matrix[50][115] * vector[50] +matrix[51][115] * vector[51] +matrix[52][115] * vector[52] +matrix[53][115] * vector[53] +matrix[54][115] * vector[54] +matrix[55][115] * vector[55] +matrix[56][115] * vector[56] +matrix[57][115] * vector[57] +matrix[58][115] * vector[58] +matrix[59][115] * vector[59] +matrix[60][115] * vector[60] +matrix[61][115] * vector[61] +matrix[62][115] * vector[62] +matrix[63][115] * vector[63] +matrix[64][115] * vector[64] +matrix[65][115] * vector[65] +matrix[66][115] * vector[66] +matrix[67][115] * vector[67] +matrix[68][115] * vector[68] +matrix[69][115] * vector[69] +matrix[70][115] * vector[70] +matrix[71][115] * vector[71] +matrix[72][115] * vector[72] +matrix[73][115] * vector[73] +matrix[74][115] * vector[74] +matrix[75][115] * vector[75] +matrix[76][115] * vector[76] +matrix[77][115] * vector[77] +matrix[78][115] * vector[78] +matrix[79][115] * vector[79] +matrix[80][115] * vector[80] +matrix[81][115] * vector[81] +matrix[82][115] * vector[82] +matrix[83][115] * vector[83] +matrix[84][115] * vector[84] +matrix[85][115] * vector[85] +matrix[86][115] * vector[86] +matrix[87][115] * vector[87] +matrix[88][115] * vector[88] +matrix[89][115] * vector[89] +matrix[90][115] * vector[90] +matrix[91][115] * vector[91] +matrix[92][115] * vector[92] +matrix[93][115] * vector[93] +matrix[94][115] * vector[94] +matrix[95][115] * vector[95] +matrix[96][115] * vector[96] +matrix[97][115] * vector[97] +matrix[98][115] * vector[98] +matrix[99][115] * vector[99] +b[115];
assign result[116] = matrix[0][116] * vector[0] +matrix[1][116] * vector[1] +matrix[2][116] * vector[2] +matrix[3][116] * vector[3] +matrix[4][116] * vector[4] +matrix[5][116] * vector[5] +matrix[6][116] * vector[6] +matrix[7][116] * vector[7] +matrix[8][116] * vector[8] +matrix[9][116] * vector[9] +matrix[10][116] * vector[10] +matrix[11][116] * vector[11] +matrix[12][116] * vector[12] +matrix[13][116] * vector[13] +matrix[14][116] * vector[14] +matrix[15][116] * vector[15] +matrix[16][116] * vector[16] +matrix[17][116] * vector[17] +matrix[18][116] * vector[18] +matrix[19][116] * vector[19] +matrix[20][116] * vector[20] +matrix[21][116] * vector[21] +matrix[22][116] * vector[22] +matrix[23][116] * vector[23] +matrix[24][116] * vector[24] +matrix[25][116] * vector[25] +matrix[26][116] * vector[26] +matrix[27][116] * vector[27] +matrix[28][116] * vector[28] +matrix[29][116] * vector[29] +matrix[30][116] * vector[30] +matrix[31][116] * vector[31] +matrix[32][116] * vector[32] +matrix[33][116] * vector[33] +matrix[34][116] * vector[34] +matrix[35][116] * vector[35] +matrix[36][116] * vector[36] +matrix[37][116] * vector[37] +matrix[38][116] * vector[38] +matrix[39][116] * vector[39] +matrix[40][116] * vector[40] +matrix[41][116] * vector[41] +matrix[42][116] * vector[42] +matrix[43][116] * vector[43] +matrix[44][116] * vector[44] +matrix[45][116] * vector[45] +matrix[46][116] * vector[46] +matrix[47][116] * vector[47] +matrix[48][116] * vector[48] +matrix[49][116] * vector[49] +matrix[50][116] * vector[50] +matrix[51][116] * vector[51] +matrix[52][116] * vector[52] +matrix[53][116] * vector[53] +matrix[54][116] * vector[54] +matrix[55][116] * vector[55] +matrix[56][116] * vector[56] +matrix[57][116] * vector[57] +matrix[58][116] * vector[58] +matrix[59][116] * vector[59] +matrix[60][116] * vector[60] +matrix[61][116] * vector[61] +matrix[62][116] * vector[62] +matrix[63][116] * vector[63] +matrix[64][116] * vector[64] +matrix[65][116] * vector[65] +matrix[66][116] * vector[66] +matrix[67][116] * vector[67] +matrix[68][116] * vector[68] +matrix[69][116] * vector[69] +matrix[70][116] * vector[70] +matrix[71][116] * vector[71] +matrix[72][116] * vector[72] +matrix[73][116] * vector[73] +matrix[74][116] * vector[74] +matrix[75][116] * vector[75] +matrix[76][116] * vector[76] +matrix[77][116] * vector[77] +matrix[78][116] * vector[78] +matrix[79][116] * vector[79] +matrix[80][116] * vector[80] +matrix[81][116] * vector[81] +matrix[82][116] * vector[82] +matrix[83][116] * vector[83] +matrix[84][116] * vector[84] +matrix[85][116] * vector[85] +matrix[86][116] * vector[86] +matrix[87][116] * vector[87] +matrix[88][116] * vector[88] +matrix[89][116] * vector[89] +matrix[90][116] * vector[90] +matrix[91][116] * vector[91] +matrix[92][116] * vector[92] +matrix[93][116] * vector[93] +matrix[94][116] * vector[94] +matrix[95][116] * vector[95] +matrix[96][116] * vector[96] +matrix[97][116] * vector[97] +matrix[98][116] * vector[98] +matrix[99][116] * vector[99] +b[116];
assign result[117] = matrix[0][117] * vector[0] +matrix[1][117] * vector[1] +matrix[2][117] * vector[2] +matrix[3][117] * vector[3] +matrix[4][117] * vector[4] +matrix[5][117] * vector[5] +matrix[6][117] * vector[6] +matrix[7][117] * vector[7] +matrix[8][117] * vector[8] +matrix[9][117] * vector[9] +matrix[10][117] * vector[10] +matrix[11][117] * vector[11] +matrix[12][117] * vector[12] +matrix[13][117] * vector[13] +matrix[14][117] * vector[14] +matrix[15][117] * vector[15] +matrix[16][117] * vector[16] +matrix[17][117] * vector[17] +matrix[18][117] * vector[18] +matrix[19][117] * vector[19] +matrix[20][117] * vector[20] +matrix[21][117] * vector[21] +matrix[22][117] * vector[22] +matrix[23][117] * vector[23] +matrix[24][117] * vector[24] +matrix[25][117] * vector[25] +matrix[26][117] * vector[26] +matrix[27][117] * vector[27] +matrix[28][117] * vector[28] +matrix[29][117] * vector[29] +matrix[30][117] * vector[30] +matrix[31][117] * vector[31] +matrix[32][117] * vector[32] +matrix[33][117] * vector[33] +matrix[34][117] * vector[34] +matrix[35][117] * vector[35] +matrix[36][117] * vector[36] +matrix[37][117] * vector[37] +matrix[38][117] * vector[38] +matrix[39][117] * vector[39] +matrix[40][117] * vector[40] +matrix[41][117] * vector[41] +matrix[42][117] * vector[42] +matrix[43][117] * vector[43] +matrix[44][117] * vector[44] +matrix[45][117] * vector[45] +matrix[46][117] * vector[46] +matrix[47][117] * vector[47] +matrix[48][117] * vector[48] +matrix[49][117] * vector[49] +matrix[50][117] * vector[50] +matrix[51][117] * vector[51] +matrix[52][117] * vector[52] +matrix[53][117] * vector[53] +matrix[54][117] * vector[54] +matrix[55][117] * vector[55] +matrix[56][117] * vector[56] +matrix[57][117] * vector[57] +matrix[58][117] * vector[58] +matrix[59][117] * vector[59] +matrix[60][117] * vector[60] +matrix[61][117] * vector[61] +matrix[62][117] * vector[62] +matrix[63][117] * vector[63] +matrix[64][117] * vector[64] +matrix[65][117] * vector[65] +matrix[66][117] * vector[66] +matrix[67][117] * vector[67] +matrix[68][117] * vector[68] +matrix[69][117] * vector[69] +matrix[70][117] * vector[70] +matrix[71][117] * vector[71] +matrix[72][117] * vector[72] +matrix[73][117] * vector[73] +matrix[74][117] * vector[74] +matrix[75][117] * vector[75] +matrix[76][117] * vector[76] +matrix[77][117] * vector[77] +matrix[78][117] * vector[78] +matrix[79][117] * vector[79] +matrix[80][117] * vector[80] +matrix[81][117] * vector[81] +matrix[82][117] * vector[82] +matrix[83][117] * vector[83] +matrix[84][117] * vector[84] +matrix[85][117] * vector[85] +matrix[86][117] * vector[86] +matrix[87][117] * vector[87] +matrix[88][117] * vector[88] +matrix[89][117] * vector[89] +matrix[90][117] * vector[90] +matrix[91][117] * vector[91] +matrix[92][117] * vector[92] +matrix[93][117] * vector[93] +matrix[94][117] * vector[94] +matrix[95][117] * vector[95] +matrix[96][117] * vector[96] +matrix[97][117] * vector[97] +matrix[98][117] * vector[98] +matrix[99][117] * vector[99] +b[117];
assign result[118] = matrix[0][118] * vector[0] +matrix[1][118] * vector[1] +matrix[2][118] * vector[2] +matrix[3][118] * vector[3] +matrix[4][118] * vector[4] +matrix[5][118] * vector[5] +matrix[6][118] * vector[6] +matrix[7][118] * vector[7] +matrix[8][118] * vector[8] +matrix[9][118] * vector[9] +matrix[10][118] * vector[10] +matrix[11][118] * vector[11] +matrix[12][118] * vector[12] +matrix[13][118] * vector[13] +matrix[14][118] * vector[14] +matrix[15][118] * vector[15] +matrix[16][118] * vector[16] +matrix[17][118] * vector[17] +matrix[18][118] * vector[18] +matrix[19][118] * vector[19] +matrix[20][118] * vector[20] +matrix[21][118] * vector[21] +matrix[22][118] * vector[22] +matrix[23][118] * vector[23] +matrix[24][118] * vector[24] +matrix[25][118] * vector[25] +matrix[26][118] * vector[26] +matrix[27][118] * vector[27] +matrix[28][118] * vector[28] +matrix[29][118] * vector[29] +matrix[30][118] * vector[30] +matrix[31][118] * vector[31] +matrix[32][118] * vector[32] +matrix[33][118] * vector[33] +matrix[34][118] * vector[34] +matrix[35][118] * vector[35] +matrix[36][118] * vector[36] +matrix[37][118] * vector[37] +matrix[38][118] * vector[38] +matrix[39][118] * vector[39] +matrix[40][118] * vector[40] +matrix[41][118] * vector[41] +matrix[42][118] * vector[42] +matrix[43][118] * vector[43] +matrix[44][118] * vector[44] +matrix[45][118] * vector[45] +matrix[46][118] * vector[46] +matrix[47][118] * vector[47] +matrix[48][118] * vector[48] +matrix[49][118] * vector[49] +matrix[50][118] * vector[50] +matrix[51][118] * vector[51] +matrix[52][118] * vector[52] +matrix[53][118] * vector[53] +matrix[54][118] * vector[54] +matrix[55][118] * vector[55] +matrix[56][118] * vector[56] +matrix[57][118] * vector[57] +matrix[58][118] * vector[58] +matrix[59][118] * vector[59] +matrix[60][118] * vector[60] +matrix[61][118] * vector[61] +matrix[62][118] * vector[62] +matrix[63][118] * vector[63] +matrix[64][118] * vector[64] +matrix[65][118] * vector[65] +matrix[66][118] * vector[66] +matrix[67][118] * vector[67] +matrix[68][118] * vector[68] +matrix[69][118] * vector[69] +matrix[70][118] * vector[70] +matrix[71][118] * vector[71] +matrix[72][118] * vector[72] +matrix[73][118] * vector[73] +matrix[74][118] * vector[74] +matrix[75][118] * vector[75] +matrix[76][118] * vector[76] +matrix[77][118] * vector[77] +matrix[78][118] * vector[78] +matrix[79][118] * vector[79] +matrix[80][118] * vector[80] +matrix[81][118] * vector[81] +matrix[82][118] * vector[82] +matrix[83][118] * vector[83] +matrix[84][118] * vector[84] +matrix[85][118] * vector[85] +matrix[86][118] * vector[86] +matrix[87][118] * vector[87] +matrix[88][118] * vector[88] +matrix[89][118] * vector[89] +matrix[90][118] * vector[90] +matrix[91][118] * vector[91] +matrix[92][118] * vector[92] +matrix[93][118] * vector[93] +matrix[94][118] * vector[94] +matrix[95][118] * vector[95] +matrix[96][118] * vector[96] +matrix[97][118] * vector[97] +matrix[98][118] * vector[98] +matrix[99][118] * vector[99] +b[118];
assign result[119] = matrix[0][119] * vector[0] +matrix[1][119] * vector[1] +matrix[2][119] * vector[2] +matrix[3][119] * vector[3] +matrix[4][119] * vector[4] +matrix[5][119] * vector[5] +matrix[6][119] * vector[6] +matrix[7][119] * vector[7] +matrix[8][119] * vector[8] +matrix[9][119] * vector[9] +matrix[10][119] * vector[10] +matrix[11][119] * vector[11] +matrix[12][119] * vector[12] +matrix[13][119] * vector[13] +matrix[14][119] * vector[14] +matrix[15][119] * vector[15] +matrix[16][119] * vector[16] +matrix[17][119] * vector[17] +matrix[18][119] * vector[18] +matrix[19][119] * vector[19] +matrix[20][119] * vector[20] +matrix[21][119] * vector[21] +matrix[22][119] * vector[22] +matrix[23][119] * vector[23] +matrix[24][119] * vector[24] +matrix[25][119] * vector[25] +matrix[26][119] * vector[26] +matrix[27][119] * vector[27] +matrix[28][119] * vector[28] +matrix[29][119] * vector[29] +matrix[30][119] * vector[30] +matrix[31][119] * vector[31] +matrix[32][119] * vector[32] +matrix[33][119] * vector[33] +matrix[34][119] * vector[34] +matrix[35][119] * vector[35] +matrix[36][119] * vector[36] +matrix[37][119] * vector[37] +matrix[38][119] * vector[38] +matrix[39][119] * vector[39] +matrix[40][119] * vector[40] +matrix[41][119] * vector[41] +matrix[42][119] * vector[42] +matrix[43][119] * vector[43] +matrix[44][119] * vector[44] +matrix[45][119] * vector[45] +matrix[46][119] * vector[46] +matrix[47][119] * vector[47] +matrix[48][119] * vector[48] +matrix[49][119] * vector[49] +matrix[50][119] * vector[50] +matrix[51][119] * vector[51] +matrix[52][119] * vector[52] +matrix[53][119] * vector[53] +matrix[54][119] * vector[54] +matrix[55][119] * vector[55] +matrix[56][119] * vector[56] +matrix[57][119] * vector[57] +matrix[58][119] * vector[58] +matrix[59][119] * vector[59] +matrix[60][119] * vector[60] +matrix[61][119] * vector[61] +matrix[62][119] * vector[62] +matrix[63][119] * vector[63] +matrix[64][119] * vector[64] +matrix[65][119] * vector[65] +matrix[66][119] * vector[66] +matrix[67][119] * vector[67] +matrix[68][119] * vector[68] +matrix[69][119] * vector[69] +matrix[70][119] * vector[70] +matrix[71][119] * vector[71] +matrix[72][119] * vector[72] +matrix[73][119] * vector[73] +matrix[74][119] * vector[74] +matrix[75][119] * vector[75] +matrix[76][119] * vector[76] +matrix[77][119] * vector[77] +matrix[78][119] * vector[78] +matrix[79][119] * vector[79] +matrix[80][119] * vector[80] +matrix[81][119] * vector[81] +matrix[82][119] * vector[82] +matrix[83][119] * vector[83] +matrix[84][119] * vector[84] +matrix[85][119] * vector[85] +matrix[86][119] * vector[86] +matrix[87][119] * vector[87] +matrix[88][119] * vector[88] +matrix[89][119] * vector[89] +matrix[90][119] * vector[90] +matrix[91][119] * vector[91] +matrix[92][119] * vector[92] +matrix[93][119] * vector[93] +matrix[94][119] * vector[94] +matrix[95][119] * vector[95] +matrix[96][119] * vector[96] +matrix[97][119] * vector[97] +matrix[98][119] * vector[98] +matrix[99][119] * vector[99] +b[119];
assign result[120] = matrix[0][120] * vector[0] +matrix[1][120] * vector[1] +matrix[2][120] * vector[2] +matrix[3][120] * vector[3] +matrix[4][120] * vector[4] +matrix[5][120] * vector[5] +matrix[6][120] * vector[6] +matrix[7][120] * vector[7] +matrix[8][120] * vector[8] +matrix[9][120] * vector[9] +matrix[10][120] * vector[10] +matrix[11][120] * vector[11] +matrix[12][120] * vector[12] +matrix[13][120] * vector[13] +matrix[14][120] * vector[14] +matrix[15][120] * vector[15] +matrix[16][120] * vector[16] +matrix[17][120] * vector[17] +matrix[18][120] * vector[18] +matrix[19][120] * vector[19] +matrix[20][120] * vector[20] +matrix[21][120] * vector[21] +matrix[22][120] * vector[22] +matrix[23][120] * vector[23] +matrix[24][120] * vector[24] +matrix[25][120] * vector[25] +matrix[26][120] * vector[26] +matrix[27][120] * vector[27] +matrix[28][120] * vector[28] +matrix[29][120] * vector[29] +matrix[30][120] * vector[30] +matrix[31][120] * vector[31] +matrix[32][120] * vector[32] +matrix[33][120] * vector[33] +matrix[34][120] * vector[34] +matrix[35][120] * vector[35] +matrix[36][120] * vector[36] +matrix[37][120] * vector[37] +matrix[38][120] * vector[38] +matrix[39][120] * vector[39] +matrix[40][120] * vector[40] +matrix[41][120] * vector[41] +matrix[42][120] * vector[42] +matrix[43][120] * vector[43] +matrix[44][120] * vector[44] +matrix[45][120] * vector[45] +matrix[46][120] * vector[46] +matrix[47][120] * vector[47] +matrix[48][120] * vector[48] +matrix[49][120] * vector[49] +matrix[50][120] * vector[50] +matrix[51][120] * vector[51] +matrix[52][120] * vector[52] +matrix[53][120] * vector[53] +matrix[54][120] * vector[54] +matrix[55][120] * vector[55] +matrix[56][120] * vector[56] +matrix[57][120] * vector[57] +matrix[58][120] * vector[58] +matrix[59][120] * vector[59] +matrix[60][120] * vector[60] +matrix[61][120] * vector[61] +matrix[62][120] * vector[62] +matrix[63][120] * vector[63] +matrix[64][120] * vector[64] +matrix[65][120] * vector[65] +matrix[66][120] * vector[66] +matrix[67][120] * vector[67] +matrix[68][120] * vector[68] +matrix[69][120] * vector[69] +matrix[70][120] * vector[70] +matrix[71][120] * vector[71] +matrix[72][120] * vector[72] +matrix[73][120] * vector[73] +matrix[74][120] * vector[74] +matrix[75][120] * vector[75] +matrix[76][120] * vector[76] +matrix[77][120] * vector[77] +matrix[78][120] * vector[78] +matrix[79][120] * vector[79] +matrix[80][120] * vector[80] +matrix[81][120] * vector[81] +matrix[82][120] * vector[82] +matrix[83][120] * vector[83] +matrix[84][120] * vector[84] +matrix[85][120] * vector[85] +matrix[86][120] * vector[86] +matrix[87][120] * vector[87] +matrix[88][120] * vector[88] +matrix[89][120] * vector[89] +matrix[90][120] * vector[90] +matrix[91][120] * vector[91] +matrix[92][120] * vector[92] +matrix[93][120] * vector[93] +matrix[94][120] * vector[94] +matrix[95][120] * vector[95] +matrix[96][120] * vector[96] +matrix[97][120] * vector[97] +matrix[98][120] * vector[98] +matrix[99][120] * vector[99] +b[120];
assign result[121] = matrix[0][121] * vector[0] +matrix[1][121] * vector[1] +matrix[2][121] * vector[2] +matrix[3][121] * vector[3] +matrix[4][121] * vector[4] +matrix[5][121] * vector[5] +matrix[6][121] * vector[6] +matrix[7][121] * vector[7] +matrix[8][121] * vector[8] +matrix[9][121] * vector[9] +matrix[10][121] * vector[10] +matrix[11][121] * vector[11] +matrix[12][121] * vector[12] +matrix[13][121] * vector[13] +matrix[14][121] * vector[14] +matrix[15][121] * vector[15] +matrix[16][121] * vector[16] +matrix[17][121] * vector[17] +matrix[18][121] * vector[18] +matrix[19][121] * vector[19] +matrix[20][121] * vector[20] +matrix[21][121] * vector[21] +matrix[22][121] * vector[22] +matrix[23][121] * vector[23] +matrix[24][121] * vector[24] +matrix[25][121] * vector[25] +matrix[26][121] * vector[26] +matrix[27][121] * vector[27] +matrix[28][121] * vector[28] +matrix[29][121] * vector[29] +matrix[30][121] * vector[30] +matrix[31][121] * vector[31] +matrix[32][121] * vector[32] +matrix[33][121] * vector[33] +matrix[34][121] * vector[34] +matrix[35][121] * vector[35] +matrix[36][121] * vector[36] +matrix[37][121] * vector[37] +matrix[38][121] * vector[38] +matrix[39][121] * vector[39] +matrix[40][121] * vector[40] +matrix[41][121] * vector[41] +matrix[42][121] * vector[42] +matrix[43][121] * vector[43] +matrix[44][121] * vector[44] +matrix[45][121] * vector[45] +matrix[46][121] * vector[46] +matrix[47][121] * vector[47] +matrix[48][121] * vector[48] +matrix[49][121] * vector[49] +matrix[50][121] * vector[50] +matrix[51][121] * vector[51] +matrix[52][121] * vector[52] +matrix[53][121] * vector[53] +matrix[54][121] * vector[54] +matrix[55][121] * vector[55] +matrix[56][121] * vector[56] +matrix[57][121] * vector[57] +matrix[58][121] * vector[58] +matrix[59][121] * vector[59] +matrix[60][121] * vector[60] +matrix[61][121] * vector[61] +matrix[62][121] * vector[62] +matrix[63][121] * vector[63] +matrix[64][121] * vector[64] +matrix[65][121] * vector[65] +matrix[66][121] * vector[66] +matrix[67][121] * vector[67] +matrix[68][121] * vector[68] +matrix[69][121] * vector[69] +matrix[70][121] * vector[70] +matrix[71][121] * vector[71] +matrix[72][121] * vector[72] +matrix[73][121] * vector[73] +matrix[74][121] * vector[74] +matrix[75][121] * vector[75] +matrix[76][121] * vector[76] +matrix[77][121] * vector[77] +matrix[78][121] * vector[78] +matrix[79][121] * vector[79] +matrix[80][121] * vector[80] +matrix[81][121] * vector[81] +matrix[82][121] * vector[82] +matrix[83][121] * vector[83] +matrix[84][121] * vector[84] +matrix[85][121] * vector[85] +matrix[86][121] * vector[86] +matrix[87][121] * vector[87] +matrix[88][121] * vector[88] +matrix[89][121] * vector[89] +matrix[90][121] * vector[90] +matrix[91][121] * vector[91] +matrix[92][121] * vector[92] +matrix[93][121] * vector[93] +matrix[94][121] * vector[94] +matrix[95][121] * vector[95] +matrix[96][121] * vector[96] +matrix[97][121] * vector[97] +matrix[98][121] * vector[98] +matrix[99][121] * vector[99] +b[121];
assign result[122] = matrix[0][122] * vector[0] +matrix[1][122] * vector[1] +matrix[2][122] * vector[2] +matrix[3][122] * vector[3] +matrix[4][122] * vector[4] +matrix[5][122] * vector[5] +matrix[6][122] * vector[6] +matrix[7][122] * vector[7] +matrix[8][122] * vector[8] +matrix[9][122] * vector[9] +matrix[10][122] * vector[10] +matrix[11][122] * vector[11] +matrix[12][122] * vector[12] +matrix[13][122] * vector[13] +matrix[14][122] * vector[14] +matrix[15][122] * vector[15] +matrix[16][122] * vector[16] +matrix[17][122] * vector[17] +matrix[18][122] * vector[18] +matrix[19][122] * vector[19] +matrix[20][122] * vector[20] +matrix[21][122] * vector[21] +matrix[22][122] * vector[22] +matrix[23][122] * vector[23] +matrix[24][122] * vector[24] +matrix[25][122] * vector[25] +matrix[26][122] * vector[26] +matrix[27][122] * vector[27] +matrix[28][122] * vector[28] +matrix[29][122] * vector[29] +matrix[30][122] * vector[30] +matrix[31][122] * vector[31] +matrix[32][122] * vector[32] +matrix[33][122] * vector[33] +matrix[34][122] * vector[34] +matrix[35][122] * vector[35] +matrix[36][122] * vector[36] +matrix[37][122] * vector[37] +matrix[38][122] * vector[38] +matrix[39][122] * vector[39] +matrix[40][122] * vector[40] +matrix[41][122] * vector[41] +matrix[42][122] * vector[42] +matrix[43][122] * vector[43] +matrix[44][122] * vector[44] +matrix[45][122] * vector[45] +matrix[46][122] * vector[46] +matrix[47][122] * vector[47] +matrix[48][122] * vector[48] +matrix[49][122] * vector[49] +matrix[50][122] * vector[50] +matrix[51][122] * vector[51] +matrix[52][122] * vector[52] +matrix[53][122] * vector[53] +matrix[54][122] * vector[54] +matrix[55][122] * vector[55] +matrix[56][122] * vector[56] +matrix[57][122] * vector[57] +matrix[58][122] * vector[58] +matrix[59][122] * vector[59] +matrix[60][122] * vector[60] +matrix[61][122] * vector[61] +matrix[62][122] * vector[62] +matrix[63][122] * vector[63] +matrix[64][122] * vector[64] +matrix[65][122] * vector[65] +matrix[66][122] * vector[66] +matrix[67][122] * vector[67] +matrix[68][122] * vector[68] +matrix[69][122] * vector[69] +matrix[70][122] * vector[70] +matrix[71][122] * vector[71] +matrix[72][122] * vector[72] +matrix[73][122] * vector[73] +matrix[74][122] * vector[74] +matrix[75][122] * vector[75] +matrix[76][122] * vector[76] +matrix[77][122] * vector[77] +matrix[78][122] * vector[78] +matrix[79][122] * vector[79] +matrix[80][122] * vector[80] +matrix[81][122] * vector[81] +matrix[82][122] * vector[82] +matrix[83][122] * vector[83] +matrix[84][122] * vector[84] +matrix[85][122] * vector[85] +matrix[86][122] * vector[86] +matrix[87][122] * vector[87] +matrix[88][122] * vector[88] +matrix[89][122] * vector[89] +matrix[90][122] * vector[90] +matrix[91][122] * vector[91] +matrix[92][122] * vector[92] +matrix[93][122] * vector[93] +matrix[94][122] * vector[94] +matrix[95][122] * vector[95] +matrix[96][122] * vector[96] +matrix[97][122] * vector[97] +matrix[98][122] * vector[98] +matrix[99][122] * vector[99] +b[122];
assign result[123] = matrix[0][123] * vector[0] +matrix[1][123] * vector[1] +matrix[2][123] * vector[2] +matrix[3][123] * vector[3] +matrix[4][123] * vector[4] +matrix[5][123] * vector[5] +matrix[6][123] * vector[6] +matrix[7][123] * vector[7] +matrix[8][123] * vector[8] +matrix[9][123] * vector[9] +matrix[10][123] * vector[10] +matrix[11][123] * vector[11] +matrix[12][123] * vector[12] +matrix[13][123] * vector[13] +matrix[14][123] * vector[14] +matrix[15][123] * vector[15] +matrix[16][123] * vector[16] +matrix[17][123] * vector[17] +matrix[18][123] * vector[18] +matrix[19][123] * vector[19] +matrix[20][123] * vector[20] +matrix[21][123] * vector[21] +matrix[22][123] * vector[22] +matrix[23][123] * vector[23] +matrix[24][123] * vector[24] +matrix[25][123] * vector[25] +matrix[26][123] * vector[26] +matrix[27][123] * vector[27] +matrix[28][123] * vector[28] +matrix[29][123] * vector[29] +matrix[30][123] * vector[30] +matrix[31][123] * vector[31] +matrix[32][123] * vector[32] +matrix[33][123] * vector[33] +matrix[34][123] * vector[34] +matrix[35][123] * vector[35] +matrix[36][123] * vector[36] +matrix[37][123] * vector[37] +matrix[38][123] * vector[38] +matrix[39][123] * vector[39] +matrix[40][123] * vector[40] +matrix[41][123] * vector[41] +matrix[42][123] * vector[42] +matrix[43][123] * vector[43] +matrix[44][123] * vector[44] +matrix[45][123] * vector[45] +matrix[46][123] * vector[46] +matrix[47][123] * vector[47] +matrix[48][123] * vector[48] +matrix[49][123] * vector[49] +matrix[50][123] * vector[50] +matrix[51][123] * vector[51] +matrix[52][123] * vector[52] +matrix[53][123] * vector[53] +matrix[54][123] * vector[54] +matrix[55][123] * vector[55] +matrix[56][123] * vector[56] +matrix[57][123] * vector[57] +matrix[58][123] * vector[58] +matrix[59][123] * vector[59] +matrix[60][123] * vector[60] +matrix[61][123] * vector[61] +matrix[62][123] * vector[62] +matrix[63][123] * vector[63] +matrix[64][123] * vector[64] +matrix[65][123] * vector[65] +matrix[66][123] * vector[66] +matrix[67][123] * vector[67] +matrix[68][123] * vector[68] +matrix[69][123] * vector[69] +matrix[70][123] * vector[70] +matrix[71][123] * vector[71] +matrix[72][123] * vector[72] +matrix[73][123] * vector[73] +matrix[74][123] * vector[74] +matrix[75][123] * vector[75] +matrix[76][123] * vector[76] +matrix[77][123] * vector[77] +matrix[78][123] * vector[78] +matrix[79][123] * vector[79] +matrix[80][123] * vector[80] +matrix[81][123] * vector[81] +matrix[82][123] * vector[82] +matrix[83][123] * vector[83] +matrix[84][123] * vector[84] +matrix[85][123] * vector[85] +matrix[86][123] * vector[86] +matrix[87][123] * vector[87] +matrix[88][123] * vector[88] +matrix[89][123] * vector[89] +matrix[90][123] * vector[90] +matrix[91][123] * vector[91] +matrix[92][123] * vector[92] +matrix[93][123] * vector[93] +matrix[94][123] * vector[94] +matrix[95][123] * vector[95] +matrix[96][123] * vector[96] +matrix[97][123] * vector[97] +matrix[98][123] * vector[98] +matrix[99][123] * vector[99] +b[123];
assign result[124] = matrix[0][124] * vector[0] +matrix[1][124] * vector[1] +matrix[2][124] * vector[2] +matrix[3][124] * vector[3] +matrix[4][124] * vector[4] +matrix[5][124] * vector[5] +matrix[6][124] * vector[6] +matrix[7][124] * vector[7] +matrix[8][124] * vector[8] +matrix[9][124] * vector[9] +matrix[10][124] * vector[10] +matrix[11][124] * vector[11] +matrix[12][124] * vector[12] +matrix[13][124] * vector[13] +matrix[14][124] * vector[14] +matrix[15][124] * vector[15] +matrix[16][124] * vector[16] +matrix[17][124] * vector[17] +matrix[18][124] * vector[18] +matrix[19][124] * vector[19] +matrix[20][124] * vector[20] +matrix[21][124] * vector[21] +matrix[22][124] * vector[22] +matrix[23][124] * vector[23] +matrix[24][124] * vector[24] +matrix[25][124] * vector[25] +matrix[26][124] * vector[26] +matrix[27][124] * vector[27] +matrix[28][124] * vector[28] +matrix[29][124] * vector[29] +matrix[30][124] * vector[30] +matrix[31][124] * vector[31] +matrix[32][124] * vector[32] +matrix[33][124] * vector[33] +matrix[34][124] * vector[34] +matrix[35][124] * vector[35] +matrix[36][124] * vector[36] +matrix[37][124] * vector[37] +matrix[38][124] * vector[38] +matrix[39][124] * vector[39] +matrix[40][124] * vector[40] +matrix[41][124] * vector[41] +matrix[42][124] * vector[42] +matrix[43][124] * vector[43] +matrix[44][124] * vector[44] +matrix[45][124] * vector[45] +matrix[46][124] * vector[46] +matrix[47][124] * vector[47] +matrix[48][124] * vector[48] +matrix[49][124] * vector[49] +matrix[50][124] * vector[50] +matrix[51][124] * vector[51] +matrix[52][124] * vector[52] +matrix[53][124] * vector[53] +matrix[54][124] * vector[54] +matrix[55][124] * vector[55] +matrix[56][124] * vector[56] +matrix[57][124] * vector[57] +matrix[58][124] * vector[58] +matrix[59][124] * vector[59] +matrix[60][124] * vector[60] +matrix[61][124] * vector[61] +matrix[62][124] * vector[62] +matrix[63][124] * vector[63] +matrix[64][124] * vector[64] +matrix[65][124] * vector[65] +matrix[66][124] * vector[66] +matrix[67][124] * vector[67] +matrix[68][124] * vector[68] +matrix[69][124] * vector[69] +matrix[70][124] * vector[70] +matrix[71][124] * vector[71] +matrix[72][124] * vector[72] +matrix[73][124] * vector[73] +matrix[74][124] * vector[74] +matrix[75][124] * vector[75] +matrix[76][124] * vector[76] +matrix[77][124] * vector[77] +matrix[78][124] * vector[78] +matrix[79][124] * vector[79] +matrix[80][124] * vector[80] +matrix[81][124] * vector[81] +matrix[82][124] * vector[82] +matrix[83][124] * vector[83] +matrix[84][124] * vector[84] +matrix[85][124] * vector[85] +matrix[86][124] * vector[86] +matrix[87][124] * vector[87] +matrix[88][124] * vector[88] +matrix[89][124] * vector[89] +matrix[90][124] * vector[90] +matrix[91][124] * vector[91] +matrix[92][124] * vector[92] +matrix[93][124] * vector[93] +matrix[94][124] * vector[94] +matrix[95][124] * vector[95] +matrix[96][124] * vector[96] +matrix[97][124] * vector[97] +matrix[98][124] * vector[98] +matrix[99][124] * vector[99] +b[124];
assign result[125] = matrix[0][125] * vector[0] +matrix[1][125] * vector[1] +matrix[2][125] * vector[2] +matrix[3][125] * vector[3] +matrix[4][125] * vector[4] +matrix[5][125] * vector[5] +matrix[6][125] * vector[6] +matrix[7][125] * vector[7] +matrix[8][125] * vector[8] +matrix[9][125] * vector[9] +matrix[10][125] * vector[10] +matrix[11][125] * vector[11] +matrix[12][125] * vector[12] +matrix[13][125] * vector[13] +matrix[14][125] * vector[14] +matrix[15][125] * vector[15] +matrix[16][125] * vector[16] +matrix[17][125] * vector[17] +matrix[18][125] * vector[18] +matrix[19][125] * vector[19] +matrix[20][125] * vector[20] +matrix[21][125] * vector[21] +matrix[22][125] * vector[22] +matrix[23][125] * vector[23] +matrix[24][125] * vector[24] +matrix[25][125] * vector[25] +matrix[26][125] * vector[26] +matrix[27][125] * vector[27] +matrix[28][125] * vector[28] +matrix[29][125] * vector[29] +matrix[30][125] * vector[30] +matrix[31][125] * vector[31] +matrix[32][125] * vector[32] +matrix[33][125] * vector[33] +matrix[34][125] * vector[34] +matrix[35][125] * vector[35] +matrix[36][125] * vector[36] +matrix[37][125] * vector[37] +matrix[38][125] * vector[38] +matrix[39][125] * vector[39] +matrix[40][125] * vector[40] +matrix[41][125] * vector[41] +matrix[42][125] * vector[42] +matrix[43][125] * vector[43] +matrix[44][125] * vector[44] +matrix[45][125] * vector[45] +matrix[46][125] * vector[46] +matrix[47][125] * vector[47] +matrix[48][125] * vector[48] +matrix[49][125] * vector[49] +matrix[50][125] * vector[50] +matrix[51][125] * vector[51] +matrix[52][125] * vector[52] +matrix[53][125] * vector[53] +matrix[54][125] * vector[54] +matrix[55][125] * vector[55] +matrix[56][125] * vector[56] +matrix[57][125] * vector[57] +matrix[58][125] * vector[58] +matrix[59][125] * vector[59] +matrix[60][125] * vector[60] +matrix[61][125] * vector[61] +matrix[62][125] * vector[62] +matrix[63][125] * vector[63] +matrix[64][125] * vector[64] +matrix[65][125] * vector[65] +matrix[66][125] * vector[66] +matrix[67][125] * vector[67] +matrix[68][125] * vector[68] +matrix[69][125] * vector[69] +matrix[70][125] * vector[70] +matrix[71][125] * vector[71] +matrix[72][125] * vector[72] +matrix[73][125] * vector[73] +matrix[74][125] * vector[74] +matrix[75][125] * vector[75] +matrix[76][125] * vector[76] +matrix[77][125] * vector[77] +matrix[78][125] * vector[78] +matrix[79][125] * vector[79] +matrix[80][125] * vector[80] +matrix[81][125] * vector[81] +matrix[82][125] * vector[82] +matrix[83][125] * vector[83] +matrix[84][125] * vector[84] +matrix[85][125] * vector[85] +matrix[86][125] * vector[86] +matrix[87][125] * vector[87] +matrix[88][125] * vector[88] +matrix[89][125] * vector[89] +matrix[90][125] * vector[90] +matrix[91][125] * vector[91] +matrix[92][125] * vector[92] +matrix[93][125] * vector[93] +matrix[94][125] * vector[94] +matrix[95][125] * vector[95] +matrix[96][125] * vector[96] +matrix[97][125] * vector[97] +matrix[98][125] * vector[98] +matrix[99][125] * vector[99] +b[125];
assign result[126] = matrix[0][126] * vector[0] +matrix[1][126] * vector[1] +matrix[2][126] * vector[2] +matrix[3][126] * vector[3] +matrix[4][126] * vector[4] +matrix[5][126] * vector[5] +matrix[6][126] * vector[6] +matrix[7][126] * vector[7] +matrix[8][126] * vector[8] +matrix[9][126] * vector[9] +matrix[10][126] * vector[10] +matrix[11][126] * vector[11] +matrix[12][126] * vector[12] +matrix[13][126] * vector[13] +matrix[14][126] * vector[14] +matrix[15][126] * vector[15] +matrix[16][126] * vector[16] +matrix[17][126] * vector[17] +matrix[18][126] * vector[18] +matrix[19][126] * vector[19] +matrix[20][126] * vector[20] +matrix[21][126] * vector[21] +matrix[22][126] * vector[22] +matrix[23][126] * vector[23] +matrix[24][126] * vector[24] +matrix[25][126] * vector[25] +matrix[26][126] * vector[26] +matrix[27][126] * vector[27] +matrix[28][126] * vector[28] +matrix[29][126] * vector[29] +matrix[30][126] * vector[30] +matrix[31][126] * vector[31] +matrix[32][126] * vector[32] +matrix[33][126] * vector[33] +matrix[34][126] * vector[34] +matrix[35][126] * vector[35] +matrix[36][126] * vector[36] +matrix[37][126] * vector[37] +matrix[38][126] * vector[38] +matrix[39][126] * vector[39] +matrix[40][126] * vector[40] +matrix[41][126] * vector[41] +matrix[42][126] * vector[42] +matrix[43][126] * vector[43] +matrix[44][126] * vector[44] +matrix[45][126] * vector[45] +matrix[46][126] * vector[46] +matrix[47][126] * vector[47] +matrix[48][126] * vector[48] +matrix[49][126] * vector[49] +matrix[50][126] * vector[50] +matrix[51][126] * vector[51] +matrix[52][126] * vector[52] +matrix[53][126] * vector[53] +matrix[54][126] * vector[54] +matrix[55][126] * vector[55] +matrix[56][126] * vector[56] +matrix[57][126] * vector[57] +matrix[58][126] * vector[58] +matrix[59][126] * vector[59] +matrix[60][126] * vector[60] +matrix[61][126] * vector[61] +matrix[62][126] * vector[62] +matrix[63][126] * vector[63] +matrix[64][126] * vector[64] +matrix[65][126] * vector[65] +matrix[66][126] * vector[66] +matrix[67][126] * vector[67] +matrix[68][126] * vector[68] +matrix[69][126] * vector[69] +matrix[70][126] * vector[70] +matrix[71][126] * vector[71] +matrix[72][126] * vector[72] +matrix[73][126] * vector[73] +matrix[74][126] * vector[74] +matrix[75][126] * vector[75] +matrix[76][126] * vector[76] +matrix[77][126] * vector[77] +matrix[78][126] * vector[78] +matrix[79][126] * vector[79] +matrix[80][126] * vector[80] +matrix[81][126] * vector[81] +matrix[82][126] * vector[82] +matrix[83][126] * vector[83] +matrix[84][126] * vector[84] +matrix[85][126] * vector[85] +matrix[86][126] * vector[86] +matrix[87][126] * vector[87] +matrix[88][126] * vector[88] +matrix[89][126] * vector[89] +matrix[90][126] * vector[90] +matrix[91][126] * vector[91] +matrix[92][126] * vector[92] +matrix[93][126] * vector[93] +matrix[94][126] * vector[94] +matrix[95][126] * vector[95] +matrix[96][126] * vector[96] +matrix[97][126] * vector[97] +matrix[98][126] * vector[98] +matrix[99][126] * vector[99] +b[126];
assign result[127] = matrix[0][127] * vector[0] +matrix[1][127] * vector[1] +matrix[2][127] * vector[2] +matrix[3][127] * vector[3] +matrix[4][127] * vector[4] +matrix[5][127] * vector[5] +matrix[6][127] * vector[6] +matrix[7][127] * vector[7] +matrix[8][127] * vector[8] +matrix[9][127] * vector[9] +matrix[10][127] * vector[10] +matrix[11][127] * vector[11] +matrix[12][127] * vector[12] +matrix[13][127] * vector[13] +matrix[14][127] * vector[14] +matrix[15][127] * vector[15] +matrix[16][127] * vector[16] +matrix[17][127] * vector[17] +matrix[18][127] * vector[18] +matrix[19][127] * vector[19] +matrix[20][127] * vector[20] +matrix[21][127] * vector[21] +matrix[22][127] * vector[22] +matrix[23][127] * vector[23] +matrix[24][127] * vector[24] +matrix[25][127] * vector[25] +matrix[26][127] * vector[26] +matrix[27][127] * vector[27] +matrix[28][127] * vector[28] +matrix[29][127] * vector[29] +matrix[30][127] * vector[30] +matrix[31][127] * vector[31] +matrix[32][127] * vector[32] +matrix[33][127] * vector[33] +matrix[34][127] * vector[34] +matrix[35][127] * vector[35] +matrix[36][127] * vector[36] +matrix[37][127] * vector[37] +matrix[38][127] * vector[38] +matrix[39][127] * vector[39] +matrix[40][127] * vector[40] +matrix[41][127] * vector[41] +matrix[42][127] * vector[42] +matrix[43][127] * vector[43] +matrix[44][127] * vector[44] +matrix[45][127] * vector[45] +matrix[46][127] * vector[46] +matrix[47][127] * vector[47] +matrix[48][127] * vector[48] +matrix[49][127] * vector[49] +matrix[50][127] * vector[50] +matrix[51][127] * vector[51] +matrix[52][127] * vector[52] +matrix[53][127] * vector[53] +matrix[54][127] * vector[54] +matrix[55][127] * vector[55] +matrix[56][127] * vector[56] +matrix[57][127] * vector[57] +matrix[58][127] * vector[58] +matrix[59][127] * vector[59] +matrix[60][127] * vector[60] +matrix[61][127] * vector[61] +matrix[62][127] * vector[62] +matrix[63][127] * vector[63] +matrix[64][127] * vector[64] +matrix[65][127] * vector[65] +matrix[66][127] * vector[66] +matrix[67][127] * vector[67] +matrix[68][127] * vector[68] +matrix[69][127] * vector[69] +matrix[70][127] * vector[70] +matrix[71][127] * vector[71] +matrix[72][127] * vector[72] +matrix[73][127] * vector[73] +matrix[74][127] * vector[74] +matrix[75][127] * vector[75] +matrix[76][127] * vector[76] +matrix[77][127] * vector[77] +matrix[78][127] * vector[78] +matrix[79][127] * vector[79] +matrix[80][127] * vector[80] +matrix[81][127] * vector[81] +matrix[82][127] * vector[82] +matrix[83][127] * vector[83] +matrix[84][127] * vector[84] +matrix[85][127] * vector[85] +matrix[86][127] * vector[86] +matrix[87][127] * vector[87] +matrix[88][127] * vector[88] +matrix[89][127] * vector[89] +matrix[90][127] * vector[90] +matrix[91][127] * vector[91] +matrix[92][127] * vector[92] +matrix[93][127] * vector[93] +matrix[94][127] * vector[94] +matrix[95][127] * vector[95] +matrix[96][127] * vector[96] +matrix[97][127] * vector[97] +matrix[98][127] * vector[98] +matrix[99][127] * vector[99] +b[127];
assign result[128] = matrix[0][128] * vector[0] +matrix[1][128] * vector[1] +matrix[2][128] * vector[2] +matrix[3][128] * vector[3] +matrix[4][128] * vector[4] +matrix[5][128] * vector[5] +matrix[6][128] * vector[6] +matrix[7][128] * vector[7] +matrix[8][128] * vector[8] +matrix[9][128] * vector[9] +matrix[10][128] * vector[10] +matrix[11][128] * vector[11] +matrix[12][128] * vector[12] +matrix[13][128] * vector[13] +matrix[14][128] * vector[14] +matrix[15][128] * vector[15] +matrix[16][128] * vector[16] +matrix[17][128] * vector[17] +matrix[18][128] * vector[18] +matrix[19][128] * vector[19] +matrix[20][128] * vector[20] +matrix[21][128] * vector[21] +matrix[22][128] * vector[22] +matrix[23][128] * vector[23] +matrix[24][128] * vector[24] +matrix[25][128] * vector[25] +matrix[26][128] * vector[26] +matrix[27][128] * vector[27] +matrix[28][128] * vector[28] +matrix[29][128] * vector[29] +matrix[30][128] * vector[30] +matrix[31][128] * vector[31] +matrix[32][128] * vector[32] +matrix[33][128] * vector[33] +matrix[34][128] * vector[34] +matrix[35][128] * vector[35] +matrix[36][128] * vector[36] +matrix[37][128] * vector[37] +matrix[38][128] * vector[38] +matrix[39][128] * vector[39] +matrix[40][128] * vector[40] +matrix[41][128] * vector[41] +matrix[42][128] * vector[42] +matrix[43][128] * vector[43] +matrix[44][128] * vector[44] +matrix[45][128] * vector[45] +matrix[46][128] * vector[46] +matrix[47][128] * vector[47] +matrix[48][128] * vector[48] +matrix[49][128] * vector[49] +matrix[50][128] * vector[50] +matrix[51][128] * vector[51] +matrix[52][128] * vector[52] +matrix[53][128] * vector[53] +matrix[54][128] * vector[54] +matrix[55][128] * vector[55] +matrix[56][128] * vector[56] +matrix[57][128] * vector[57] +matrix[58][128] * vector[58] +matrix[59][128] * vector[59] +matrix[60][128] * vector[60] +matrix[61][128] * vector[61] +matrix[62][128] * vector[62] +matrix[63][128] * vector[63] +matrix[64][128] * vector[64] +matrix[65][128] * vector[65] +matrix[66][128] * vector[66] +matrix[67][128] * vector[67] +matrix[68][128] * vector[68] +matrix[69][128] * vector[69] +matrix[70][128] * vector[70] +matrix[71][128] * vector[71] +matrix[72][128] * vector[72] +matrix[73][128] * vector[73] +matrix[74][128] * vector[74] +matrix[75][128] * vector[75] +matrix[76][128] * vector[76] +matrix[77][128] * vector[77] +matrix[78][128] * vector[78] +matrix[79][128] * vector[79] +matrix[80][128] * vector[80] +matrix[81][128] * vector[81] +matrix[82][128] * vector[82] +matrix[83][128] * vector[83] +matrix[84][128] * vector[84] +matrix[85][128] * vector[85] +matrix[86][128] * vector[86] +matrix[87][128] * vector[87] +matrix[88][128] * vector[88] +matrix[89][128] * vector[89] +matrix[90][128] * vector[90] +matrix[91][128] * vector[91] +matrix[92][128] * vector[92] +matrix[93][128] * vector[93] +matrix[94][128] * vector[94] +matrix[95][128] * vector[95] +matrix[96][128] * vector[96] +matrix[97][128] * vector[97] +matrix[98][128] * vector[98] +matrix[99][128] * vector[99] +b[128];
assign result[129] = matrix[0][129] * vector[0] +matrix[1][129] * vector[1] +matrix[2][129] * vector[2] +matrix[3][129] * vector[3] +matrix[4][129] * vector[4] +matrix[5][129] * vector[5] +matrix[6][129] * vector[6] +matrix[7][129] * vector[7] +matrix[8][129] * vector[8] +matrix[9][129] * vector[9] +matrix[10][129] * vector[10] +matrix[11][129] * vector[11] +matrix[12][129] * vector[12] +matrix[13][129] * vector[13] +matrix[14][129] * vector[14] +matrix[15][129] * vector[15] +matrix[16][129] * vector[16] +matrix[17][129] * vector[17] +matrix[18][129] * vector[18] +matrix[19][129] * vector[19] +matrix[20][129] * vector[20] +matrix[21][129] * vector[21] +matrix[22][129] * vector[22] +matrix[23][129] * vector[23] +matrix[24][129] * vector[24] +matrix[25][129] * vector[25] +matrix[26][129] * vector[26] +matrix[27][129] * vector[27] +matrix[28][129] * vector[28] +matrix[29][129] * vector[29] +matrix[30][129] * vector[30] +matrix[31][129] * vector[31] +matrix[32][129] * vector[32] +matrix[33][129] * vector[33] +matrix[34][129] * vector[34] +matrix[35][129] * vector[35] +matrix[36][129] * vector[36] +matrix[37][129] * vector[37] +matrix[38][129] * vector[38] +matrix[39][129] * vector[39] +matrix[40][129] * vector[40] +matrix[41][129] * vector[41] +matrix[42][129] * vector[42] +matrix[43][129] * vector[43] +matrix[44][129] * vector[44] +matrix[45][129] * vector[45] +matrix[46][129] * vector[46] +matrix[47][129] * vector[47] +matrix[48][129] * vector[48] +matrix[49][129] * vector[49] +matrix[50][129] * vector[50] +matrix[51][129] * vector[51] +matrix[52][129] * vector[52] +matrix[53][129] * vector[53] +matrix[54][129] * vector[54] +matrix[55][129] * vector[55] +matrix[56][129] * vector[56] +matrix[57][129] * vector[57] +matrix[58][129] * vector[58] +matrix[59][129] * vector[59] +matrix[60][129] * vector[60] +matrix[61][129] * vector[61] +matrix[62][129] * vector[62] +matrix[63][129] * vector[63] +matrix[64][129] * vector[64] +matrix[65][129] * vector[65] +matrix[66][129] * vector[66] +matrix[67][129] * vector[67] +matrix[68][129] * vector[68] +matrix[69][129] * vector[69] +matrix[70][129] * vector[70] +matrix[71][129] * vector[71] +matrix[72][129] * vector[72] +matrix[73][129] * vector[73] +matrix[74][129] * vector[74] +matrix[75][129] * vector[75] +matrix[76][129] * vector[76] +matrix[77][129] * vector[77] +matrix[78][129] * vector[78] +matrix[79][129] * vector[79] +matrix[80][129] * vector[80] +matrix[81][129] * vector[81] +matrix[82][129] * vector[82] +matrix[83][129] * vector[83] +matrix[84][129] * vector[84] +matrix[85][129] * vector[85] +matrix[86][129] * vector[86] +matrix[87][129] * vector[87] +matrix[88][129] * vector[88] +matrix[89][129] * vector[89] +matrix[90][129] * vector[90] +matrix[91][129] * vector[91] +matrix[92][129] * vector[92] +matrix[93][129] * vector[93] +matrix[94][129] * vector[94] +matrix[95][129] * vector[95] +matrix[96][129] * vector[96] +matrix[97][129] * vector[97] +matrix[98][129] * vector[98] +matrix[99][129] * vector[99] +b[129];
assign result[130] = matrix[0][130] * vector[0] +matrix[1][130] * vector[1] +matrix[2][130] * vector[2] +matrix[3][130] * vector[3] +matrix[4][130] * vector[4] +matrix[5][130] * vector[5] +matrix[6][130] * vector[6] +matrix[7][130] * vector[7] +matrix[8][130] * vector[8] +matrix[9][130] * vector[9] +matrix[10][130] * vector[10] +matrix[11][130] * vector[11] +matrix[12][130] * vector[12] +matrix[13][130] * vector[13] +matrix[14][130] * vector[14] +matrix[15][130] * vector[15] +matrix[16][130] * vector[16] +matrix[17][130] * vector[17] +matrix[18][130] * vector[18] +matrix[19][130] * vector[19] +matrix[20][130] * vector[20] +matrix[21][130] * vector[21] +matrix[22][130] * vector[22] +matrix[23][130] * vector[23] +matrix[24][130] * vector[24] +matrix[25][130] * vector[25] +matrix[26][130] * vector[26] +matrix[27][130] * vector[27] +matrix[28][130] * vector[28] +matrix[29][130] * vector[29] +matrix[30][130] * vector[30] +matrix[31][130] * vector[31] +matrix[32][130] * vector[32] +matrix[33][130] * vector[33] +matrix[34][130] * vector[34] +matrix[35][130] * vector[35] +matrix[36][130] * vector[36] +matrix[37][130] * vector[37] +matrix[38][130] * vector[38] +matrix[39][130] * vector[39] +matrix[40][130] * vector[40] +matrix[41][130] * vector[41] +matrix[42][130] * vector[42] +matrix[43][130] * vector[43] +matrix[44][130] * vector[44] +matrix[45][130] * vector[45] +matrix[46][130] * vector[46] +matrix[47][130] * vector[47] +matrix[48][130] * vector[48] +matrix[49][130] * vector[49] +matrix[50][130] * vector[50] +matrix[51][130] * vector[51] +matrix[52][130] * vector[52] +matrix[53][130] * vector[53] +matrix[54][130] * vector[54] +matrix[55][130] * vector[55] +matrix[56][130] * vector[56] +matrix[57][130] * vector[57] +matrix[58][130] * vector[58] +matrix[59][130] * vector[59] +matrix[60][130] * vector[60] +matrix[61][130] * vector[61] +matrix[62][130] * vector[62] +matrix[63][130] * vector[63] +matrix[64][130] * vector[64] +matrix[65][130] * vector[65] +matrix[66][130] * vector[66] +matrix[67][130] * vector[67] +matrix[68][130] * vector[68] +matrix[69][130] * vector[69] +matrix[70][130] * vector[70] +matrix[71][130] * vector[71] +matrix[72][130] * vector[72] +matrix[73][130] * vector[73] +matrix[74][130] * vector[74] +matrix[75][130] * vector[75] +matrix[76][130] * vector[76] +matrix[77][130] * vector[77] +matrix[78][130] * vector[78] +matrix[79][130] * vector[79] +matrix[80][130] * vector[80] +matrix[81][130] * vector[81] +matrix[82][130] * vector[82] +matrix[83][130] * vector[83] +matrix[84][130] * vector[84] +matrix[85][130] * vector[85] +matrix[86][130] * vector[86] +matrix[87][130] * vector[87] +matrix[88][130] * vector[88] +matrix[89][130] * vector[89] +matrix[90][130] * vector[90] +matrix[91][130] * vector[91] +matrix[92][130] * vector[92] +matrix[93][130] * vector[93] +matrix[94][130] * vector[94] +matrix[95][130] * vector[95] +matrix[96][130] * vector[96] +matrix[97][130] * vector[97] +matrix[98][130] * vector[98] +matrix[99][130] * vector[99] +b[130];
assign result[131] = matrix[0][131] * vector[0] +matrix[1][131] * vector[1] +matrix[2][131] * vector[2] +matrix[3][131] * vector[3] +matrix[4][131] * vector[4] +matrix[5][131] * vector[5] +matrix[6][131] * vector[6] +matrix[7][131] * vector[7] +matrix[8][131] * vector[8] +matrix[9][131] * vector[9] +matrix[10][131] * vector[10] +matrix[11][131] * vector[11] +matrix[12][131] * vector[12] +matrix[13][131] * vector[13] +matrix[14][131] * vector[14] +matrix[15][131] * vector[15] +matrix[16][131] * vector[16] +matrix[17][131] * vector[17] +matrix[18][131] * vector[18] +matrix[19][131] * vector[19] +matrix[20][131] * vector[20] +matrix[21][131] * vector[21] +matrix[22][131] * vector[22] +matrix[23][131] * vector[23] +matrix[24][131] * vector[24] +matrix[25][131] * vector[25] +matrix[26][131] * vector[26] +matrix[27][131] * vector[27] +matrix[28][131] * vector[28] +matrix[29][131] * vector[29] +matrix[30][131] * vector[30] +matrix[31][131] * vector[31] +matrix[32][131] * vector[32] +matrix[33][131] * vector[33] +matrix[34][131] * vector[34] +matrix[35][131] * vector[35] +matrix[36][131] * vector[36] +matrix[37][131] * vector[37] +matrix[38][131] * vector[38] +matrix[39][131] * vector[39] +matrix[40][131] * vector[40] +matrix[41][131] * vector[41] +matrix[42][131] * vector[42] +matrix[43][131] * vector[43] +matrix[44][131] * vector[44] +matrix[45][131] * vector[45] +matrix[46][131] * vector[46] +matrix[47][131] * vector[47] +matrix[48][131] * vector[48] +matrix[49][131] * vector[49] +matrix[50][131] * vector[50] +matrix[51][131] * vector[51] +matrix[52][131] * vector[52] +matrix[53][131] * vector[53] +matrix[54][131] * vector[54] +matrix[55][131] * vector[55] +matrix[56][131] * vector[56] +matrix[57][131] * vector[57] +matrix[58][131] * vector[58] +matrix[59][131] * vector[59] +matrix[60][131] * vector[60] +matrix[61][131] * vector[61] +matrix[62][131] * vector[62] +matrix[63][131] * vector[63] +matrix[64][131] * vector[64] +matrix[65][131] * vector[65] +matrix[66][131] * vector[66] +matrix[67][131] * vector[67] +matrix[68][131] * vector[68] +matrix[69][131] * vector[69] +matrix[70][131] * vector[70] +matrix[71][131] * vector[71] +matrix[72][131] * vector[72] +matrix[73][131] * vector[73] +matrix[74][131] * vector[74] +matrix[75][131] * vector[75] +matrix[76][131] * vector[76] +matrix[77][131] * vector[77] +matrix[78][131] * vector[78] +matrix[79][131] * vector[79] +matrix[80][131] * vector[80] +matrix[81][131] * vector[81] +matrix[82][131] * vector[82] +matrix[83][131] * vector[83] +matrix[84][131] * vector[84] +matrix[85][131] * vector[85] +matrix[86][131] * vector[86] +matrix[87][131] * vector[87] +matrix[88][131] * vector[88] +matrix[89][131] * vector[89] +matrix[90][131] * vector[90] +matrix[91][131] * vector[91] +matrix[92][131] * vector[92] +matrix[93][131] * vector[93] +matrix[94][131] * vector[94] +matrix[95][131] * vector[95] +matrix[96][131] * vector[96] +matrix[97][131] * vector[97] +matrix[98][131] * vector[98] +matrix[99][131] * vector[99] +b[131];
assign result[132] = matrix[0][132] * vector[0] +matrix[1][132] * vector[1] +matrix[2][132] * vector[2] +matrix[3][132] * vector[3] +matrix[4][132] * vector[4] +matrix[5][132] * vector[5] +matrix[6][132] * vector[6] +matrix[7][132] * vector[7] +matrix[8][132] * vector[8] +matrix[9][132] * vector[9] +matrix[10][132] * vector[10] +matrix[11][132] * vector[11] +matrix[12][132] * vector[12] +matrix[13][132] * vector[13] +matrix[14][132] * vector[14] +matrix[15][132] * vector[15] +matrix[16][132] * vector[16] +matrix[17][132] * vector[17] +matrix[18][132] * vector[18] +matrix[19][132] * vector[19] +matrix[20][132] * vector[20] +matrix[21][132] * vector[21] +matrix[22][132] * vector[22] +matrix[23][132] * vector[23] +matrix[24][132] * vector[24] +matrix[25][132] * vector[25] +matrix[26][132] * vector[26] +matrix[27][132] * vector[27] +matrix[28][132] * vector[28] +matrix[29][132] * vector[29] +matrix[30][132] * vector[30] +matrix[31][132] * vector[31] +matrix[32][132] * vector[32] +matrix[33][132] * vector[33] +matrix[34][132] * vector[34] +matrix[35][132] * vector[35] +matrix[36][132] * vector[36] +matrix[37][132] * vector[37] +matrix[38][132] * vector[38] +matrix[39][132] * vector[39] +matrix[40][132] * vector[40] +matrix[41][132] * vector[41] +matrix[42][132] * vector[42] +matrix[43][132] * vector[43] +matrix[44][132] * vector[44] +matrix[45][132] * vector[45] +matrix[46][132] * vector[46] +matrix[47][132] * vector[47] +matrix[48][132] * vector[48] +matrix[49][132] * vector[49] +matrix[50][132] * vector[50] +matrix[51][132] * vector[51] +matrix[52][132] * vector[52] +matrix[53][132] * vector[53] +matrix[54][132] * vector[54] +matrix[55][132] * vector[55] +matrix[56][132] * vector[56] +matrix[57][132] * vector[57] +matrix[58][132] * vector[58] +matrix[59][132] * vector[59] +matrix[60][132] * vector[60] +matrix[61][132] * vector[61] +matrix[62][132] * vector[62] +matrix[63][132] * vector[63] +matrix[64][132] * vector[64] +matrix[65][132] * vector[65] +matrix[66][132] * vector[66] +matrix[67][132] * vector[67] +matrix[68][132] * vector[68] +matrix[69][132] * vector[69] +matrix[70][132] * vector[70] +matrix[71][132] * vector[71] +matrix[72][132] * vector[72] +matrix[73][132] * vector[73] +matrix[74][132] * vector[74] +matrix[75][132] * vector[75] +matrix[76][132] * vector[76] +matrix[77][132] * vector[77] +matrix[78][132] * vector[78] +matrix[79][132] * vector[79] +matrix[80][132] * vector[80] +matrix[81][132] * vector[81] +matrix[82][132] * vector[82] +matrix[83][132] * vector[83] +matrix[84][132] * vector[84] +matrix[85][132] * vector[85] +matrix[86][132] * vector[86] +matrix[87][132] * vector[87] +matrix[88][132] * vector[88] +matrix[89][132] * vector[89] +matrix[90][132] * vector[90] +matrix[91][132] * vector[91] +matrix[92][132] * vector[92] +matrix[93][132] * vector[93] +matrix[94][132] * vector[94] +matrix[95][132] * vector[95] +matrix[96][132] * vector[96] +matrix[97][132] * vector[97] +matrix[98][132] * vector[98] +matrix[99][132] * vector[99] +b[132];
assign result[133] = matrix[0][133] * vector[0] +matrix[1][133] * vector[1] +matrix[2][133] * vector[2] +matrix[3][133] * vector[3] +matrix[4][133] * vector[4] +matrix[5][133] * vector[5] +matrix[6][133] * vector[6] +matrix[7][133] * vector[7] +matrix[8][133] * vector[8] +matrix[9][133] * vector[9] +matrix[10][133] * vector[10] +matrix[11][133] * vector[11] +matrix[12][133] * vector[12] +matrix[13][133] * vector[13] +matrix[14][133] * vector[14] +matrix[15][133] * vector[15] +matrix[16][133] * vector[16] +matrix[17][133] * vector[17] +matrix[18][133] * vector[18] +matrix[19][133] * vector[19] +matrix[20][133] * vector[20] +matrix[21][133] * vector[21] +matrix[22][133] * vector[22] +matrix[23][133] * vector[23] +matrix[24][133] * vector[24] +matrix[25][133] * vector[25] +matrix[26][133] * vector[26] +matrix[27][133] * vector[27] +matrix[28][133] * vector[28] +matrix[29][133] * vector[29] +matrix[30][133] * vector[30] +matrix[31][133] * vector[31] +matrix[32][133] * vector[32] +matrix[33][133] * vector[33] +matrix[34][133] * vector[34] +matrix[35][133] * vector[35] +matrix[36][133] * vector[36] +matrix[37][133] * vector[37] +matrix[38][133] * vector[38] +matrix[39][133] * vector[39] +matrix[40][133] * vector[40] +matrix[41][133] * vector[41] +matrix[42][133] * vector[42] +matrix[43][133] * vector[43] +matrix[44][133] * vector[44] +matrix[45][133] * vector[45] +matrix[46][133] * vector[46] +matrix[47][133] * vector[47] +matrix[48][133] * vector[48] +matrix[49][133] * vector[49] +matrix[50][133] * vector[50] +matrix[51][133] * vector[51] +matrix[52][133] * vector[52] +matrix[53][133] * vector[53] +matrix[54][133] * vector[54] +matrix[55][133] * vector[55] +matrix[56][133] * vector[56] +matrix[57][133] * vector[57] +matrix[58][133] * vector[58] +matrix[59][133] * vector[59] +matrix[60][133] * vector[60] +matrix[61][133] * vector[61] +matrix[62][133] * vector[62] +matrix[63][133] * vector[63] +matrix[64][133] * vector[64] +matrix[65][133] * vector[65] +matrix[66][133] * vector[66] +matrix[67][133] * vector[67] +matrix[68][133] * vector[68] +matrix[69][133] * vector[69] +matrix[70][133] * vector[70] +matrix[71][133] * vector[71] +matrix[72][133] * vector[72] +matrix[73][133] * vector[73] +matrix[74][133] * vector[74] +matrix[75][133] * vector[75] +matrix[76][133] * vector[76] +matrix[77][133] * vector[77] +matrix[78][133] * vector[78] +matrix[79][133] * vector[79] +matrix[80][133] * vector[80] +matrix[81][133] * vector[81] +matrix[82][133] * vector[82] +matrix[83][133] * vector[83] +matrix[84][133] * vector[84] +matrix[85][133] * vector[85] +matrix[86][133] * vector[86] +matrix[87][133] * vector[87] +matrix[88][133] * vector[88] +matrix[89][133] * vector[89] +matrix[90][133] * vector[90] +matrix[91][133] * vector[91] +matrix[92][133] * vector[92] +matrix[93][133] * vector[93] +matrix[94][133] * vector[94] +matrix[95][133] * vector[95] +matrix[96][133] * vector[96] +matrix[97][133] * vector[97] +matrix[98][133] * vector[98] +matrix[99][133] * vector[99] +b[133];
assign result[134] = matrix[0][134] * vector[0] +matrix[1][134] * vector[1] +matrix[2][134] * vector[2] +matrix[3][134] * vector[3] +matrix[4][134] * vector[4] +matrix[5][134] * vector[5] +matrix[6][134] * vector[6] +matrix[7][134] * vector[7] +matrix[8][134] * vector[8] +matrix[9][134] * vector[9] +matrix[10][134] * vector[10] +matrix[11][134] * vector[11] +matrix[12][134] * vector[12] +matrix[13][134] * vector[13] +matrix[14][134] * vector[14] +matrix[15][134] * vector[15] +matrix[16][134] * vector[16] +matrix[17][134] * vector[17] +matrix[18][134] * vector[18] +matrix[19][134] * vector[19] +matrix[20][134] * vector[20] +matrix[21][134] * vector[21] +matrix[22][134] * vector[22] +matrix[23][134] * vector[23] +matrix[24][134] * vector[24] +matrix[25][134] * vector[25] +matrix[26][134] * vector[26] +matrix[27][134] * vector[27] +matrix[28][134] * vector[28] +matrix[29][134] * vector[29] +matrix[30][134] * vector[30] +matrix[31][134] * vector[31] +matrix[32][134] * vector[32] +matrix[33][134] * vector[33] +matrix[34][134] * vector[34] +matrix[35][134] * vector[35] +matrix[36][134] * vector[36] +matrix[37][134] * vector[37] +matrix[38][134] * vector[38] +matrix[39][134] * vector[39] +matrix[40][134] * vector[40] +matrix[41][134] * vector[41] +matrix[42][134] * vector[42] +matrix[43][134] * vector[43] +matrix[44][134] * vector[44] +matrix[45][134] * vector[45] +matrix[46][134] * vector[46] +matrix[47][134] * vector[47] +matrix[48][134] * vector[48] +matrix[49][134] * vector[49] +matrix[50][134] * vector[50] +matrix[51][134] * vector[51] +matrix[52][134] * vector[52] +matrix[53][134] * vector[53] +matrix[54][134] * vector[54] +matrix[55][134] * vector[55] +matrix[56][134] * vector[56] +matrix[57][134] * vector[57] +matrix[58][134] * vector[58] +matrix[59][134] * vector[59] +matrix[60][134] * vector[60] +matrix[61][134] * vector[61] +matrix[62][134] * vector[62] +matrix[63][134] * vector[63] +matrix[64][134] * vector[64] +matrix[65][134] * vector[65] +matrix[66][134] * vector[66] +matrix[67][134] * vector[67] +matrix[68][134] * vector[68] +matrix[69][134] * vector[69] +matrix[70][134] * vector[70] +matrix[71][134] * vector[71] +matrix[72][134] * vector[72] +matrix[73][134] * vector[73] +matrix[74][134] * vector[74] +matrix[75][134] * vector[75] +matrix[76][134] * vector[76] +matrix[77][134] * vector[77] +matrix[78][134] * vector[78] +matrix[79][134] * vector[79] +matrix[80][134] * vector[80] +matrix[81][134] * vector[81] +matrix[82][134] * vector[82] +matrix[83][134] * vector[83] +matrix[84][134] * vector[84] +matrix[85][134] * vector[85] +matrix[86][134] * vector[86] +matrix[87][134] * vector[87] +matrix[88][134] * vector[88] +matrix[89][134] * vector[89] +matrix[90][134] * vector[90] +matrix[91][134] * vector[91] +matrix[92][134] * vector[92] +matrix[93][134] * vector[93] +matrix[94][134] * vector[94] +matrix[95][134] * vector[95] +matrix[96][134] * vector[96] +matrix[97][134] * vector[97] +matrix[98][134] * vector[98] +matrix[99][134] * vector[99] +b[134];
assign result[135] = matrix[0][135] * vector[0] +matrix[1][135] * vector[1] +matrix[2][135] * vector[2] +matrix[3][135] * vector[3] +matrix[4][135] * vector[4] +matrix[5][135] * vector[5] +matrix[6][135] * vector[6] +matrix[7][135] * vector[7] +matrix[8][135] * vector[8] +matrix[9][135] * vector[9] +matrix[10][135] * vector[10] +matrix[11][135] * vector[11] +matrix[12][135] * vector[12] +matrix[13][135] * vector[13] +matrix[14][135] * vector[14] +matrix[15][135] * vector[15] +matrix[16][135] * vector[16] +matrix[17][135] * vector[17] +matrix[18][135] * vector[18] +matrix[19][135] * vector[19] +matrix[20][135] * vector[20] +matrix[21][135] * vector[21] +matrix[22][135] * vector[22] +matrix[23][135] * vector[23] +matrix[24][135] * vector[24] +matrix[25][135] * vector[25] +matrix[26][135] * vector[26] +matrix[27][135] * vector[27] +matrix[28][135] * vector[28] +matrix[29][135] * vector[29] +matrix[30][135] * vector[30] +matrix[31][135] * vector[31] +matrix[32][135] * vector[32] +matrix[33][135] * vector[33] +matrix[34][135] * vector[34] +matrix[35][135] * vector[35] +matrix[36][135] * vector[36] +matrix[37][135] * vector[37] +matrix[38][135] * vector[38] +matrix[39][135] * vector[39] +matrix[40][135] * vector[40] +matrix[41][135] * vector[41] +matrix[42][135] * vector[42] +matrix[43][135] * vector[43] +matrix[44][135] * vector[44] +matrix[45][135] * vector[45] +matrix[46][135] * vector[46] +matrix[47][135] * vector[47] +matrix[48][135] * vector[48] +matrix[49][135] * vector[49] +matrix[50][135] * vector[50] +matrix[51][135] * vector[51] +matrix[52][135] * vector[52] +matrix[53][135] * vector[53] +matrix[54][135] * vector[54] +matrix[55][135] * vector[55] +matrix[56][135] * vector[56] +matrix[57][135] * vector[57] +matrix[58][135] * vector[58] +matrix[59][135] * vector[59] +matrix[60][135] * vector[60] +matrix[61][135] * vector[61] +matrix[62][135] * vector[62] +matrix[63][135] * vector[63] +matrix[64][135] * vector[64] +matrix[65][135] * vector[65] +matrix[66][135] * vector[66] +matrix[67][135] * vector[67] +matrix[68][135] * vector[68] +matrix[69][135] * vector[69] +matrix[70][135] * vector[70] +matrix[71][135] * vector[71] +matrix[72][135] * vector[72] +matrix[73][135] * vector[73] +matrix[74][135] * vector[74] +matrix[75][135] * vector[75] +matrix[76][135] * vector[76] +matrix[77][135] * vector[77] +matrix[78][135] * vector[78] +matrix[79][135] * vector[79] +matrix[80][135] * vector[80] +matrix[81][135] * vector[81] +matrix[82][135] * vector[82] +matrix[83][135] * vector[83] +matrix[84][135] * vector[84] +matrix[85][135] * vector[85] +matrix[86][135] * vector[86] +matrix[87][135] * vector[87] +matrix[88][135] * vector[88] +matrix[89][135] * vector[89] +matrix[90][135] * vector[90] +matrix[91][135] * vector[91] +matrix[92][135] * vector[92] +matrix[93][135] * vector[93] +matrix[94][135] * vector[94] +matrix[95][135] * vector[95] +matrix[96][135] * vector[96] +matrix[97][135] * vector[97] +matrix[98][135] * vector[98] +matrix[99][135] * vector[99] +b[135];
assign result[136] = matrix[0][136] * vector[0] +matrix[1][136] * vector[1] +matrix[2][136] * vector[2] +matrix[3][136] * vector[3] +matrix[4][136] * vector[4] +matrix[5][136] * vector[5] +matrix[6][136] * vector[6] +matrix[7][136] * vector[7] +matrix[8][136] * vector[8] +matrix[9][136] * vector[9] +matrix[10][136] * vector[10] +matrix[11][136] * vector[11] +matrix[12][136] * vector[12] +matrix[13][136] * vector[13] +matrix[14][136] * vector[14] +matrix[15][136] * vector[15] +matrix[16][136] * vector[16] +matrix[17][136] * vector[17] +matrix[18][136] * vector[18] +matrix[19][136] * vector[19] +matrix[20][136] * vector[20] +matrix[21][136] * vector[21] +matrix[22][136] * vector[22] +matrix[23][136] * vector[23] +matrix[24][136] * vector[24] +matrix[25][136] * vector[25] +matrix[26][136] * vector[26] +matrix[27][136] * vector[27] +matrix[28][136] * vector[28] +matrix[29][136] * vector[29] +matrix[30][136] * vector[30] +matrix[31][136] * vector[31] +matrix[32][136] * vector[32] +matrix[33][136] * vector[33] +matrix[34][136] * vector[34] +matrix[35][136] * vector[35] +matrix[36][136] * vector[36] +matrix[37][136] * vector[37] +matrix[38][136] * vector[38] +matrix[39][136] * vector[39] +matrix[40][136] * vector[40] +matrix[41][136] * vector[41] +matrix[42][136] * vector[42] +matrix[43][136] * vector[43] +matrix[44][136] * vector[44] +matrix[45][136] * vector[45] +matrix[46][136] * vector[46] +matrix[47][136] * vector[47] +matrix[48][136] * vector[48] +matrix[49][136] * vector[49] +matrix[50][136] * vector[50] +matrix[51][136] * vector[51] +matrix[52][136] * vector[52] +matrix[53][136] * vector[53] +matrix[54][136] * vector[54] +matrix[55][136] * vector[55] +matrix[56][136] * vector[56] +matrix[57][136] * vector[57] +matrix[58][136] * vector[58] +matrix[59][136] * vector[59] +matrix[60][136] * vector[60] +matrix[61][136] * vector[61] +matrix[62][136] * vector[62] +matrix[63][136] * vector[63] +matrix[64][136] * vector[64] +matrix[65][136] * vector[65] +matrix[66][136] * vector[66] +matrix[67][136] * vector[67] +matrix[68][136] * vector[68] +matrix[69][136] * vector[69] +matrix[70][136] * vector[70] +matrix[71][136] * vector[71] +matrix[72][136] * vector[72] +matrix[73][136] * vector[73] +matrix[74][136] * vector[74] +matrix[75][136] * vector[75] +matrix[76][136] * vector[76] +matrix[77][136] * vector[77] +matrix[78][136] * vector[78] +matrix[79][136] * vector[79] +matrix[80][136] * vector[80] +matrix[81][136] * vector[81] +matrix[82][136] * vector[82] +matrix[83][136] * vector[83] +matrix[84][136] * vector[84] +matrix[85][136] * vector[85] +matrix[86][136] * vector[86] +matrix[87][136] * vector[87] +matrix[88][136] * vector[88] +matrix[89][136] * vector[89] +matrix[90][136] * vector[90] +matrix[91][136] * vector[91] +matrix[92][136] * vector[92] +matrix[93][136] * vector[93] +matrix[94][136] * vector[94] +matrix[95][136] * vector[95] +matrix[96][136] * vector[96] +matrix[97][136] * vector[97] +matrix[98][136] * vector[98] +matrix[99][136] * vector[99] +b[136];
assign result[137] = matrix[0][137] * vector[0] +matrix[1][137] * vector[1] +matrix[2][137] * vector[2] +matrix[3][137] * vector[3] +matrix[4][137] * vector[4] +matrix[5][137] * vector[5] +matrix[6][137] * vector[6] +matrix[7][137] * vector[7] +matrix[8][137] * vector[8] +matrix[9][137] * vector[9] +matrix[10][137] * vector[10] +matrix[11][137] * vector[11] +matrix[12][137] * vector[12] +matrix[13][137] * vector[13] +matrix[14][137] * vector[14] +matrix[15][137] * vector[15] +matrix[16][137] * vector[16] +matrix[17][137] * vector[17] +matrix[18][137] * vector[18] +matrix[19][137] * vector[19] +matrix[20][137] * vector[20] +matrix[21][137] * vector[21] +matrix[22][137] * vector[22] +matrix[23][137] * vector[23] +matrix[24][137] * vector[24] +matrix[25][137] * vector[25] +matrix[26][137] * vector[26] +matrix[27][137] * vector[27] +matrix[28][137] * vector[28] +matrix[29][137] * vector[29] +matrix[30][137] * vector[30] +matrix[31][137] * vector[31] +matrix[32][137] * vector[32] +matrix[33][137] * vector[33] +matrix[34][137] * vector[34] +matrix[35][137] * vector[35] +matrix[36][137] * vector[36] +matrix[37][137] * vector[37] +matrix[38][137] * vector[38] +matrix[39][137] * vector[39] +matrix[40][137] * vector[40] +matrix[41][137] * vector[41] +matrix[42][137] * vector[42] +matrix[43][137] * vector[43] +matrix[44][137] * vector[44] +matrix[45][137] * vector[45] +matrix[46][137] * vector[46] +matrix[47][137] * vector[47] +matrix[48][137] * vector[48] +matrix[49][137] * vector[49] +matrix[50][137] * vector[50] +matrix[51][137] * vector[51] +matrix[52][137] * vector[52] +matrix[53][137] * vector[53] +matrix[54][137] * vector[54] +matrix[55][137] * vector[55] +matrix[56][137] * vector[56] +matrix[57][137] * vector[57] +matrix[58][137] * vector[58] +matrix[59][137] * vector[59] +matrix[60][137] * vector[60] +matrix[61][137] * vector[61] +matrix[62][137] * vector[62] +matrix[63][137] * vector[63] +matrix[64][137] * vector[64] +matrix[65][137] * vector[65] +matrix[66][137] * vector[66] +matrix[67][137] * vector[67] +matrix[68][137] * vector[68] +matrix[69][137] * vector[69] +matrix[70][137] * vector[70] +matrix[71][137] * vector[71] +matrix[72][137] * vector[72] +matrix[73][137] * vector[73] +matrix[74][137] * vector[74] +matrix[75][137] * vector[75] +matrix[76][137] * vector[76] +matrix[77][137] * vector[77] +matrix[78][137] * vector[78] +matrix[79][137] * vector[79] +matrix[80][137] * vector[80] +matrix[81][137] * vector[81] +matrix[82][137] * vector[82] +matrix[83][137] * vector[83] +matrix[84][137] * vector[84] +matrix[85][137] * vector[85] +matrix[86][137] * vector[86] +matrix[87][137] * vector[87] +matrix[88][137] * vector[88] +matrix[89][137] * vector[89] +matrix[90][137] * vector[90] +matrix[91][137] * vector[91] +matrix[92][137] * vector[92] +matrix[93][137] * vector[93] +matrix[94][137] * vector[94] +matrix[95][137] * vector[95] +matrix[96][137] * vector[96] +matrix[97][137] * vector[97] +matrix[98][137] * vector[98] +matrix[99][137] * vector[99] +b[137];
assign result[138] = matrix[0][138] * vector[0] +matrix[1][138] * vector[1] +matrix[2][138] * vector[2] +matrix[3][138] * vector[3] +matrix[4][138] * vector[4] +matrix[5][138] * vector[5] +matrix[6][138] * vector[6] +matrix[7][138] * vector[7] +matrix[8][138] * vector[8] +matrix[9][138] * vector[9] +matrix[10][138] * vector[10] +matrix[11][138] * vector[11] +matrix[12][138] * vector[12] +matrix[13][138] * vector[13] +matrix[14][138] * vector[14] +matrix[15][138] * vector[15] +matrix[16][138] * vector[16] +matrix[17][138] * vector[17] +matrix[18][138] * vector[18] +matrix[19][138] * vector[19] +matrix[20][138] * vector[20] +matrix[21][138] * vector[21] +matrix[22][138] * vector[22] +matrix[23][138] * vector[23] +matrix[24][138] * vector[24] +matrix[25][138] * vector[25] +matrix[26][138] * vector[26] +matrix[27][138] * vector[27] +matrix[28][138] * vector[28] +matrix[29][138] * vector[29] +matrix[30][138] * vector[30] +matrix[31][138] * vector[31] +matrix[32][138] * vector[32] +matrix[33][138] * vector[33] +matrix[34][138] * vector[34] +matrix[35][138] * vector[35] +matrix[36][138] * vector[36] +matrix[37][138] * vector[37] +matrix[38][138] * vector[38] +matrix[39][138] * vector[39] +matrix[40][138] * vector[40] +matrix[41][138] * vector[41] +matrix[42][138] * vector[42] +matrix[43][138] * vector[43] +matrix[44][138] * vector[44] +matrix[45][138] * vector[45] +matrix[46][138] * vector[46] +matrix[47][138] * vector[47] +matrix[48][138] * vector[48] +matrix[49][138] * vector[49] +matrix[50][138] * vector[50] +matrix[51][138] * vector[51] +matrix[52][138] * vector[52] +matrix[53][138] * vector[53] +matrix[54][138] * vector[54] +matrix[55][138] * vector[55] +matrix[56][138] * vector[56] +matrix[57][138] * vector[57] +matrix[58][138] * vector[58] +matrix[59][138] * vector[59] +matrix[60][138] * vector[60] +matrix[61][138] * vector[61] +matrix[62][138] * vector[62] +matrix[63][138] * vector[63] +matrix[64][138] * vector[64] +matrix[65][138] * vector[65] +matrix[66][138] * vector[66] +matrix[67][138] * vector[67] +matrix[68][138] * vector[68] +matrix[69][138] * vector[69] +matrix[70][138] * vector[70] +matrix[71][138] * vector[71] +matrix[72][138] * vector[72] +matrix[73][138] * vector[73] +matrix[74][138] * vector[74] +matrix[75][138] * vector[75] +matrix[76][138] * vector[76] +matrix[77][138] * vector[77] +matrix[78][138] * vector[78] +matrix[79][138] * vector[79] +matrix[80][138] * vector[80] +matrix[81][138] * vector[81] +matrix[82][138] * vector[82] +matrix[83][138] * vector[83] +matrix[84][138] * vector[84] +matrix[85][138] * vector[85] +matrix[86][138] * vector[86] +matrix[87][138] * vector[87] +matrix[88][138] * vector[88] +matrix[89][138] * vector[89] +matrix[90][138] * vector[90] +matrix[91][138] * vector[91] +matrix[92][138] * vector[92] +matrix[93][138] * vector[93] +matrix[94][138] * vector[94] +matrix[95][138] * vector[95] +matrix[96][138] * vector[96] +matrix[97][138] * vector[97] +matrix[98][138] * vector[98] +matrix[99][138] * vector[99] +b[138];
assign result[139] = matrix[0][139] * vector[0] +matrix[1][139] * vector[1] +matrix[2][139] * vector[2] +matrix[3][139] * vector[3] +matrix[4][139] * vector[4] +matrix[5][139] * vector[5] +matrix[6][139] * vector[6] +matrix[7][139] * vector[7] +matrix[8][139] * vector[8] +matrix[9][139] * vector[9] +matrix[10][139] * vector[10] +matrix[11][139] * vector[11] +matrix[12][139] * vector[12] +matrix[13][139] * vector[13] +matrix[14][139] * vector[14] +matrix[15][139] * vector[15] +matrix[16][139] * vector[16] +matrix[17][139] * vector[17] +matrix[18][139] * vector[18] +matrix[19][139] * vector[19] +matrix[20][139] * vector[20] +matrix[21][139] * vector[21] +matrix[22][139] * vector[22] +matrix[23][139] * vector[23] +matrix[24][139] * vector[24] +matrix[25][139] * vector[25] +matrix[26][139] * vector[26] +matrix[27][139] * vector[27] +matrix[28][139] * vector[28] +matrix[29][139] * vector[29] +matrix[30][139] * vector[30] +matrix[31][139] * vector[31] +matrix[32][139] * vector[32] +matrix[33][139] * vector[33] +matrix[34][139] * vector[34] +matrix[35][139] * vector[35] +matrix[36][139] * vector[36] +matrix[37][139] * vector[37] +matrix[38][139] * vector[38] +matrix[39][139] * vector[39] +matrix[40][139] * vector[40] +matrix[41][139] * vector[41] +matrix[42][139] * vector[42] +matrix[43][139] * vector[43] +matrix[44][139] * vector[44] +matrix[45][139] * vector[45] +matrix[46][139] * vector[46] +matrix[47][139] * vector[47] +matrix[48][139] * vector[48] +matrix[49][139] * vector[49] +matrix[50][139] * vector[50] +matrix[51][139] * vector[51] +matrix[52][139] * vector[52] +matrix[53][139] * vector[53] +matrix[54][139] * vector[54] +matrix[55][139] * vector[55] +matrix[56][139] * vector[56] +matrix[57][139] * vector[57] +matrix[58][139] * vector[58] +matrix[59][139] * vector[59] +matrix[60][139] * vector[60] +matrix[61][139] * vector[61] +matrix[62][139] * vector[62] +matrix[63][139] * vector[63] +matrix[64][139] * vector[64] +matrix[65][139] * vector[65] +matrix[66][139] * vector[66] +matrix[67][139] * vector[67] +matrix[68][139] * vector[68] +matrix[69][139] * vector[69] +matrix[70][139] * vector[70] +matrix[71][139] * vector[71] +matrix[72][139] * vector[72] +matrix[73][139] * vector[73] +matrix[74][139] * vector[74] +matrix[75][139] * vector[75] +matrix[76][139] * vector[76] +matrix[77][139] * vector[77] +matrix[78][139] * vector[78] +matrix[79][139] * vector[79] +matrix[80][139] * vector[80] +matrix[81][139] * vector[81] +matrix[82][139] * vector[82] +matrix[83][139] * vector[83] +matrix[84][139] * vector[84] +matrix[85][139] * vector[85] +matrix[86][139] * vector[86] +matrix[87][139] * vector[87] +matrix[88][139] * vector[88] +matrix[89][139] * vector[89] +matrix[90][139] * vector[90] +matrix[91][139] * vector[91] +matrix[92][139] * vector[92] +matrix[93][139] * vector[93] +matrix[94][139] * vector[94] +matrix[95][139] * vector[95] +matrix[96][139] * vector[96] +matrix[97][139] * vector[97] +matrix[98][139] * vector[98] +matrix[99][139] * vector[99] +b[139];
assign result[140] = matrix[0][140] * vector[0] +matrix[1][140] * vector[1] +matrix[2][140] * vector[2] +matrix[3][140] * vector[3] +matrix[4][140] * vector[4] +matrix[5][140] * vector[5] +matrix[6][140] * vector[6] +matrix[7][140] * vector[7] +matrix[8][140] * vector[8] +matrix[9][140] * vector[9] +matrix[10][140] * vector[10] +matrix[11][140] * vector[11] +matrix[12][140] * vector[12] +matrix[13][140] * vector[13] +matrix[14][140] * vector[14] +matrix[15][140] * vector[15] +matrix[16][140] * vector[16] +matrix[17][140] * vector[17] +matrix[18][140] * vector[18] +matrix[19][140] * vector[19] +matrix[20][140] * vector[20] +matrix[21][140] * vector[21] +matrix[22][140] * vector[22] +matrix[23][140] * vector[23] +matrix[24][140] * vector[24] +matrix[25][140] * vector[25] +matrix[26][140] * vector[26] +matrix[27][140] * vector[27] +matrix[28][140] * vector[28] +matrix[29][140] * vector[29] +matrix[30][140] * vector[30] +matrix[31][140] * vector[31] +matrix[32][140] * vector[32] +matrix[33][140] * vector[33] +matrix[34][140] * vector[34] +matrix[35][140] * vector[35] +matrix[36][140] * vector[36] +matrix[37][140] * vector[37] +matrix[38][140] * vector[38] +matrix[39][140] * vector[39] +matrix[40][140] * vector[40] +matrix[41][140] * vector[41] +matrix[42][140] * vector[42] +matrix[43][140] * vector[43] +matrix[44][140] * vector[44] +matrix[45][140] * vector[45] +matrix[46][140] * vector[46] +matrix[47][140] * vector[47] +matrix[48][140] * vector[48] +matrix[49][140] * vector[49] +matrix[50][140] * vector[50] +matrix[51][140] * vector[51] +matrix[52][140] * vector[52] +matrix[53][140] * vector[53] +matrix[54][140] * vector[54] +matrix[55][140] * vector[55] +matrix[56][140] * vector[56] +matrix[57][140] * vector[57] +matrix[58][140] * vector[58] +matrix[59][140] * vector[59] +matrix[60][140] * vector[60] +matrix[61][140] * vector[61] +matrix[62][140] * vector[62] +matrix[63][140] * vector[63] +matrix[64][140] * vector[64] +matrix[65][140] * vector[65] +matrix[66][140] * vector[66] +matrix[67][140] * vector[67] +matrix[68][140] * vector[68] +matrix[69][140] * vector[69] +matrix[70][140] * vector[70] +matrix[71][140] * vector[71] +matrix[72][140] * vector[72] +matrix[73][140] * vector[73] +matrix[74][140] * vector[74] +matrix[75][140] * vector[75] +matrix[76][140] * vector[76] +matrix[77][140] * vector[77] +matrix[78][140] * vector[78] +matrix[79][140] * vector[79] +matrix[80][140] * vector[80] +matrix[81][140] * vector[81] +matrix[82][140] * vector[82] +matrix[83][140] * vector[83] +matrix[84][140] * vector[84] +matrix[85][140] * vector[85] +matrix[86][140] * vector[86] +matrix[87][140] * vector[87] +matrix[88][140] * vector[88] +matrix[89][140] * vector[89] +matrix[90][140] * vector[90] +matrix[91][140] * vector[91] +matrix[92][140] * vector[92] +matrix[93][140] * vector[93] +matrix[94][140] * vector[94] +matrix[95][140] * vector[95] +matrix[96][140] * vector[96] +matrix[97][140] * vector[97] +matrix[98][140] * vector[98] +matrix[99][140] * vector[99] +b[140];
assign result[141] = matrix[0][141] * vector[0] +matrix[1][141] * vector[1] +matrix[2][141] * vector[2] +matrix[3][141] * vector[3] +matrix[4][141] * vector[4] +matrix[5][141] * vector[5] +matrix[6][141] * vector[6] +matrix[7][141] * vector[7] +matrix[8][141] * vector[8] +matrix[9][141] * vector[9] +matrix[10][141] * vector[10] +matrix[11][141] * vector[11] +matrix[12][141] * vector[12] +matrix[13][141] * vector[13] +matrix[14][141] * vector[14] +matrix[15][141] * vector[15] +matrix[16][141] * vector[16] +matrix[17][141] * vector[17] +matrix[18][141] * vector[18] +matrix[19][141] * vector[19] +matrix[20][141] * vector[20] +matrix[21][141] * vector[21] +matrix[22][141] * vector[22] +matrix[23][141] * vector[23] +matrix[24][141] * vector[24] +matrix[25][141] * vector[25] +matrix[26][141] * vector[26] +matrix[27][141] * vector[27] +matrix[28][141] * vector[28] +matrix[29][141] * vector[29] +matrix[30][141] * vector[30] +matrix[31][141] * vector[31] +matrix[32][141] * vector[32] +matrix[33][141] * vector[33] +matrix[34][141] * vector[34] +matrix[35][141] * vector[35] +matrix[36][141] * vector[36] +matrix[37][141] * vector[37] +matrix[38][141] * vector[38] +matrix[39][141] * vector[39] +matrix[40][141] * vector[40] +matrix[41][141] * vector[41] +matrix[42][141] * vector[42] +matrix[43][141] * vector[43] +matrix[44][141] * vector[44] +matrix[45][141] * vector[45] +matrix[46][141] * vector[46] +matrix[47][141] * vector[47] +matrix[48][141] * vector[48] +matrix[49][141] * vector[49] +matrix[50][141] * vector[50] +matrix[51][141] * vector[51] +matrix[52][141] * vector[52] +matrix[53][141] * vector[53] +matrix[54][141] * vector[54] +matrix[55][141] * vector[55] +matrix[56][141] * vector[56] +matrix[57][141] * vector[57] +matrix[58][141] * vector[58] +matrix[59][141] * vector[59] +matrix[60][141] * vector[60] +matrix[61][141] * vector[61] +matrix[62][141] * vector[62] +matrix[63][141] * vector[63] +matrix[64][141] * vector[64] +matrix[65][141] * vector[65] +matrix[66][141] * vector[66] +matrix[67][141] * vector[67] +matrix[68][141] * vector[68] +matrix[69][141] * vector[69] +matrix[70][141] * vector[70] +matrix[71][141] * vector[71] +matrix[72][141] * vector[72] +matrix[73][141] * vector[73] +matrix[74][141] * vector[74] +matrix[75][141] * vector[75] +matrix[76][141] * vector[76] +matrix[77][141] * vector[77] +matrix[78][141] * vector[78] +matrix[79][141] * vector[79] +matrix[80][141] * vector[80] +matrix[81][141] * vector[81] +matrix[82][141] * vector[82] +matrix[83][141] * vector[83] +matrix[84][141] * vector[84] +matrix[85][141] * vector[85] +matrix[86][141] * vector[86] +matrix[87][141] * vector[87] +matrix[88][141] * vector[88] +matrix[89][141] * vector[89] +matrix[90][141] * vector[90] +matrix[91][141] * vector[91] +matrix[92][141] * vector[92] +matrix[93][141] * vector[93] +matrix[94][141] * vector[94] +matrix[95][141] * vector[95] +matrix[96][141] * vector[96] +matrix[97][141] * vector[97] +matrix[98][141] * vector[98] +matrix[99][141] * vector[99] +b[141];
assign result[142] = matrix[0][142] * vector[0] +matrix[1][142] * vector[1] +matrix[2][142] * vector[2] +matrix[3][142] * vector[3] +matrix[4][142] * vector[4] +matrix[5][142] * vector[5] +matrix[6][142] * vector[6] +matrix[7][142] * vector[7] +matrix[8][142] * vector[8] +matrix[9][142] * vector[9] +matrix[10][142] * vector[10] +matrix[11][142] * vector[11] +matrix[12][142] * vector[12] +matrix[13][142] * vector[13] +matrix[14][142] * vector[14] +matrix[15][142] * vector[15] +matrix[16][142] * vector[16] +matrix[17][142] * vector[17] +matrix[18][142] * vector[18] +matrix[19][142] * vector[19] +matrix[20][142] * vector[20] +matrix[21][142] * vector[21] +matrix[22][142] * vector[22] +matrix[23][142] * vector[23] +matrix[24][142] * vector[24] +matrix[25][142] * vector[25] +matrix[26][142] * vector[26] +matrix[27][142] * vector[27] +matrix[28][142] * vector[28] +matrix[29][142] * vector[29] +matrix[30][142] * vector[30] +matrix[31][142] * vector[31] +matrix[32][142] * vector[32] +matrix[33][142] * vector[33] +matrix[34][142] * vector[34] +matrix[35][142] * vector[35] +matrix[36][142] * vector[36] +matrix[37][142] * vector[37] +matrix[38][142] * vector[38] +matrix[39][142] * vector[39] +matrix[40][142] * vector[40] +matrix[41][142] * vector[41] +matrix[42][142] * vector[42] +matrix[43][142] * vector[43] +matrix[44][142] * vector[44] +matrix[45][142] * vector[45] +matrix[46][142] * vector[46] +matrix[47][142] * vector[47] +matrix[48][142] * vector[48] +matrix[49][142] * vector[49] +matrix[50][142] * vector[50] +matrix[51][142] * vector[51] +matrix[52][142] * vector[52] +matrix[53][142] * vector[53] +matrix[54][142] * vector[54] +matrix[55][142] * vector[55] +matrix[56][142] * vector[56] +matrix[57][142] * vector[57] +matrix[58][142] * vector[58] +matrix[59][142] * vector[59] +matrix[60][142] * vector[60] +matrix[61][142] * vector[61] +matrix[62][142] * vector[62] +matrix[63][142] * vector[63] +matrix[64][142] * vector[64] +matrix[65][142] * vector[65] +matrix[66][142] * vector[66] +matrix[67][142] * vector[67] +matrix[68][142] * vector[68] +matrix[69][142] * vector[69] +matrix[70][142] * vector[70] +matrix[71][142] * vector[71] +matrix[72][142] * vector[72] +matrix[73][142] * vector[73] +matrix[74][142] * vector[74] +matrix[75][142] * vector[75] +matrix[76][142] * vector[76] +matrix[77][142] * vector[77] +matrix[78][142] * vector[78] +matrix[79][142] * vector[79] +matrix[80][142] * vector[80] +matrix[81][142] * vector[81] +matrix[82][142] * vector[82] +matrix[83][142] * vector[83] +matrix[84][142] * vector[84] +matrix[85][142] * vector[85] +matrix[86][142] * vector[86] +matrix[87][142] * vector[87] +matrix[88][142] * vector[88] +matrix[89][142] * vector[89] +matrix[90][142] * vector[90] +matrix[91][142] * vector[91] +matrix[92][142] * vector[92] +matrix[93][142] * vector[93] +matrix[94][142] * vector[94] +matrix[95][142] * vector[95] +matrix[96][142] * vector[96] +matrix[97][142] * vector[97] +matrix[98][142] * vector[98] +matrix[99][142] * vector[99] +b[142];
assign result[143] = matrix[0][143] * vector[0] +matrix[1][143] * vector[1] +matrix[2][143] * vector[2] +matrix[3][143] * vector[3] +matrix[4][143] * vector[4] +matrix[5][143] * vector[5] +matrix[6][143] * vector[6] +matrix[7][143] * vector[7] +matrix[8][143] * vector[8] +matrix[9][143] * vector[9] +matrix[10][143] * vector[10] +matrix[11][143] * vector[11] +matrix[12][143] * vector[12] +matrix[13][143] * vector[13] +matrix[14][143] * vector[14] +matrix[15][143] * vector[15] +matrix[16][143] * vector[16] +matrix[17][143] * vector[17] +matrix[18][143] * vector[18] +matrix[19][143] * vector[19] +matrix[20][143] * vector[20] +matrix[21][143] * vector[21] +matrix[22][143] * vector[22] +matrix[23][143] * vector[23] +matrix[24][143] * vector[24] +matrix[25][143] * vector[25] +matrix[26][143] * vector[26] +matrix[27][143] * vector[27] +matrix[28][143] * vector[28] +matrix[29][143] * vector[29] +matrix[30][143] * vector[30] +matrix[31][143] * vector[31] +matrix[32][143] * vector[32] +matrix[33][143] * vector[33] +matrix[34][143] * vector[34] +matrix[35][143] * vector[35] +matrix[36][143] * vector[36] +matrix[37][143] * vector[37] +matrix[38][143] * vector[38] +matrix[39][143] * vector[39] +matrix[40][143] * vector[40] +matrix[41][143] * vector[41] +matrix[42][143] * vector[42] +matrix[43][143] * vector[43] +matrix[44][143] * vector[44] +matrix[45][143] * vector[45] +matrix[46][143] * vector[46] +matrix[47][143] * vector[47] +matrix[48][143] * vector[48] +matrix[49][143] * vector[49] +matrix[50][143] * vector[50] +matrix[51][143] * vector[51] +matrix[52][143] * vector[52] +matrix[53][143] * vector[53] +matrix[54][143] * vector[54] +matrix[55][143] * vector[55] +matrix[56][143] * vector[56] +matrix[57][143] * vector[57] +matrix[58][143] * vector[58] +matrix[59][143] * vector[59] +matrix[60][143] * vector[60] +matrix[61][143] * vector[61] +matrix[62][143] * vector[62] +matrix[63][143] * vector[63] +matrix[64][143] * vector[64] +matrix[65][143] * vector[65] +matrix[66][143] * vector[66] +matrix[67][143] * vector[67] +matrix[68][143] * vector[68] +matrix[69][143] * vector[69] +matrix[70][143] * vector[70] +matrix[71][143] * vector[71] +matrix[72][143] * vector[72] +matrix[73][143] * vector[73] +matrix[74][143] * vector[74] +matrix[75][143] * vector[75] +matrix[76][143] * vector[76] +matrix[77][143] * vector[77] +matrix[78][143] * vector[78] +matrix[79][143] * vector[79] +matrix[80][143] * vector[80] +matrix[81][143] * vector[81] +matrix[82][143] * vector[82] +matrix[83][143] * vector[83] +matrix[84][143] * vector[84] +matrix[85][143] * vector[85] +matrix[86][143] * vector[86] +matrix[87][143] * vector[87] +matrix[88][143] * vector[88] +matrix[89][143] * vector[89] +matrix[90][143] * vector[90] +matrix[91][143] * vector[91] +matrix[92][143] * vector[92] +matrix[93][143] * vector[93] +matrix[94][143] * vector[94] +matrix[95][143] * vector[95] +matrix[96][143] * vector[96] +matrix[97][143] * vector[97] +matrix[98][143] * vector[98] +matrix[99][143] * vector[99] +b[143];
assign result[144] = matrix[0][144] * vector[0] +matrix[1][144] * vector[1] +matrix[2][144] * vector[2] +matrix[3][144] * vector[3] +matrix[4][144] * vector[4] +matrix[5][144] * vector[5] +matrix[6][144] * vector[6] +matrix[7][144] * vector[7] +matrix[8][144] * vector[8] +matrix[9][144] * vector[9] +matrix[10][144] * vector[10] +matrix[11][144] * vector[11] +matrix[12][144] * vector[12] +matrix[13][144] * vector[13] +matrix[14][144] * vector[14] +matrix[15][144] * vector[15] +matrix[16][144] * vector[16] +matrix[17][144] * vector[17] +matrix[18][144] * vector[18] +matrix[19][144] * vector[19] +matrix[20][144] * vector[20] +matrix[21][144] * vector[21] +matrix[22][144] * vector[22] +matrix[23][144] * vector[23] +matrix[24][144] * vector[24] +matrix[25][144] * vector[25] +matrix[26][144] * vector[26] +matrix[27][144] * vector[27] +matrix[28][144] * vector[28] +matrix[29][144] * vector[29] +matrix[30][144] * vector[30] +matrix[31][144] * vector[31] +matrix[32][144] * vector[32] +matrix[33][144] * vector[33] +matrix[34][144] * vector[34] +matrix[35][144] * vector[35] +matrix[36][144] * vector[36] +matrix[37][144] * vector[37] +matrix[38][144] * vector[38] +matrix[39][144] * vector[39] +matrix[40][144] * vector[40] +matrix[41][144] * vector[41] +matrix[42][144] * vector[42] +matrix[43][144] * vector[43] +matrix[44][144] * vector[44] +matrix[45][144] * vector[45] +matrix[46][144] * vector[46] +matrix[47][144] * vector[47] +matrix[48][144] * vector[48] +matrix[49][144] * vector[49] +matrix[50][144] * vector[50] +matrix[51][144] * vector[51] +matrix[52][144] * vector[52] +matrix[53][144] * vector[53] +matrix[54][144] * vector[54] +matrix[55][144] * vector[55] +matrix[56][144] * vector[56] +matrix[57][144] * vector[57] +matrix[58][144] * vector[58] +matrix[59][144] * vector[59] +matrix[60][144] * vector[60] +matrix[61][144] * vector[61] +matrix[62][144] * vector[62] +matrix[63][144] * vector[63] +matrix[64][144] * vector[64] +matrix[65][144] * vector[65] +matrix[66][144] * vector[66] +matrix[67][144] * vector[67] +matrix[68][144] * vector[68] +matrix[69][144] * vector[69] +matrix[70][144] * vector[70] +matrix[71][144] * vector[71] +matrix[72][144] * vector[72] +matrix[73][144] * vector[73] +matrix[74][144] * vector[74] +matrix[75][144] * vector[75] +matrix[76][144] * vector[76] +matrix[77][144] * vector[77] +matrix[78][144] * vector[78] +matrix[79][144] * vector[79] +matrix[80][144] * vector[80] +matrix[81][144] * vector[81] +matrix[82][144] * vector[82] +matrix[83][144] * vector[83] +matrix[84][144] * vector[84] +matrix[85][144] * vector[85] +matrix[86][144] * vector[86] +matrix[87][144] * vector[87] +matrix[88][144] * vector[88] +matrix[89][144] * vector[89] +matrix[90][144] * vector[90] +matrix[91][144] * vector[91] +matrix[92][144] * vector[92] +matrix[93][144] * vector[93] +matrix[94][144] * vector[94] +matrix[95][144] * vector[95] +matrix[96][144] * vector[96] +matrix[97][144] * vector[97] +matrix[98][144] * vector[98] +matrix[99][144] * vector[99] +b[144];
assign result[145] = matrix[0][145] * vector[0] +matrix[1][145] * vector[1] +matrix[2][145] * vector[2] +matrix[3][145] * vector[3] +matrix[4][145] * vector[4] +matrix[5][145] * vector[5] +matrix[6][145] * vector[6] +matrix[7][145] * vector[7] +matrix[8][145] * vector[8] +matrix[9][145] * vector[9] +matrix[10][145] * vector[10] +matrix[11][145] * vector[11] +matrix[12][145] * vector[12] +matrix[13][145] * vector[13] +matrix[14][145] * vector[14] +matrix[15][145] * vector[15] +matrix[16][145] * vector[16] +matrix[17][145] * vector[17] +matrix[18][145] * vector[18] +matrix[19][145] * vector[19] +matrix[20][145] * vector[20] +matrix[21][145] * vector[21] +matrix[22][145] * vector[22] +matrix[23][145] * vector[23] +matrix[24][145] * vector[24] +matrix[25][145] * vector[25] +matrix[26][145] * vector[26] +matrix[27][145] * vector[27] +matrix[28][145] * vector[28] +matrix[29][145] * vector[29] +matrix[30][145] * vector[30] +matrix[31][145] * vector[31] +matrix[32][145] * vector[32] +matrix[33][145] * vector[33] +matrix[34][145] * vector[34] +matrix[35][145] * vector[35] +matrix[36][145] * vector[36] +matrix[37][145] * vector[37] +matrix[38][145] * vector[38] +matrix[39][145] * vector[39] +matrix[40][145] * vector[40] +matrix[41][145] * vector[41] +matrix[42][145] * vector[42] +matrix[43][145] * vector[43] +matrix[44][145] * vector[44] +matrix[45][145] * vector[45] +matrix[46][145] * vector[46] +matrix[47][145] * vector[47] +matrix[48][145] * vector[48] +matrix[49][145] * vector[49] +matrix[50][145] * vector[50] +matrix[51][145] * vector[51] +matrix[52][145] * vector[52] +matrix[53][145] * vector[53] +matrix[54][145] * vector[54] +matrix[55][145] * vector[55] +matrix[56][145] * vector[56] +matrix[57][145] * vector[57] +matrix[58][145] * vector[58] +matrix[59][145] * vector[59] +matrix[60][145] * vector[60] +matrix[61][145] * vector[61] +matrix[62][145] * vector[62] +matrix[63][145] * vector[63] +matrix[64][145] * vector[64] +matrix[65][145] * vector[65] +matrix[66][145] * vector[66] +matrix[67][145] * vector[67] +matrix[68][145] * vector[68] +matrix[69][145] * vector[69] +matrix[70][145] * vector[70] +matrix[71][145] * vector[71] +matrix[72][145] * vector[72] +matrix[73][145] * vector[73] +matrix[74][145] * vector[74] +matrix[75][145] * vector[75] +matrix[76][145] * vector[76] +matrix[77][145] * vector[77] +matrix[78][145] * vector[78] +matrix[79][145] * vector[79] +matrix[80][145] * vector[80] +matrix[81][145] * vector[81] +matrix[82][145] * vector[82] +matrix[83][145] * vector[83] +matrix[84][145] * vector[84] +matrix[85][145] * vector[85] +matrix[86][145] * vector[86] +matrix[87][145] * vector[87] +matrix[88][145] * vector[88] +matrix[89][145] * vector[89] +matrix[90][145] * vector[90] +matrix[91][145] * vector[91] +matrix[92][145] * vector[92] +matrix[93][145] * vector[93] +matrix[94][145] * vector[94] +matrix[95][145] * vector[95] +matrix[96][145] * vector[96] +matrix[97][145] * vector[97] +matrix[98][145] * vector[98] +matrix[99][145] * vector[99] +b[145];
assign result[146] = matrix[0][146] * vector[0] +matrix[1][146] * vector[1] +matrix[2][146] * vector[2] +matrix[3][146] * vector[3] +matrix[4][146] * vector[4] +matrix[5][146] * vector[5] +matrix[6][146] * vector[6] +matrix[7][146] * vector[7] +matrix[8][146] * vector[8] +matrix[9][146] * vector[9] +matrix[10][146] * vector[10] +matrix[11][146] * vector[11] +matrix[12][146] * vector[12] +matrix[13][146] * vector[13] +matrix[14][146] * vector[14] +matrix[15][146] * vector[15] +matrix[16][146] * vector[16] +matrix[17][146] * vector[17] +matrix[18][146] * vector[18] +matrix[19][146] * vector[19] +matrix[20][146] * vector[20] +matrix[21][146] * vector[21] +matrix[22][146] * vector[22] +matrix[23][146] * vector[23] +matrix[24][146] * vector[24] +matrix[25][146] * vector[25] +matrix[26][146] * vector[26] +matrix[27][146] * vector[27] +matrix[28][146] * vector[28] +matrix[29][146] * vector[29] +matrix[30][146] * vector[30] +matrix[31][146] * vector[31] +matrix[32][146] * vector[32] +matrix[33][146] * vector[33] +matrix[34][146] * vector[34] +matrix[35][146] * vector[35] +matrix[36][146] * vector[36] +matrix[37][146] * vector[37] +matrix[38][146] * vector[38] +matrix[39][146] * vector[39] +matrix[40][146] * vector[40] +matrix[41][146] * vector[41] +matrix[42][146] * vector[42] +matrix[43][146] * vector[43] +matrix[44][146] * vector[44] +matrix[45][146] * vector[45] +matrix[46][146] * vector[46] +matrix[47][146] * vector[47] +matrix[48][146] * vector[48] +matrix[49][146] * vector[49] +matrix[50][146] * vector[50] +matrix[51][146] * vector[51] +matrix[52][146] * vector[52] +matrix[53][146] * vector[53] +matrix[54][146] * vector[54] +matrix[55][146] * vector[55] +matrix[56][146] * vector[56] +matrix[57][146] * vector[57] +matrix[58][146] * vector[58] +matrix[59][146] * vector[59] +matrix[60][146] * vector[60] +matrix[61][146] * vector[61] +matrix[62][146] * vector[62] +matrix[63][146] * vector[63] +matrix[64][146] * vector[64] +matrix[65][146] * vector[65] +matrix[66][146] * vector[66] +matrix[67][146] * vector[67] +matrix[68][146] * vector[68] +matrix[69][146] * vector[69] +matrix[70][146] * vector[70] +matrix[71][146] * vector[71] +matrix[72][146] * vector[72] +matrix[73][146] * vector[73] +matrix[74][146] * vector[74] +matrix[75][146] * vector[75] +matrix[76][146] * vector[76] +matrix[77][146] * vector[77] +matrix[78][146] * vector[78] +matrix[79][146] * vector[79] +matrix[80][146] * vector[80] +matrix[81][146] * vector[81] +matrix[82][146] * vector[82] +matrix[83][146] * vector[83] +matrix[84][146] * vector[84] +matrix[85][146] * vector[85] +matrix[86][146] * vector[86] +matrix[87][146] * vector[87] +matrix[88][146] * vector[88] +matrix[89][146] * vector[89] +matrix[90][146] * vector[90] +matrix[91][146] * vector[91] +matrix[92][146] * vector[92] +matrix[93][146] * vector[93] +matrix[94][146] * vector[94] +matrix[95][146] * vector[95] +matrix[96][146] * vector[96] +matrix[97][146] * vector[97] +matrix[98][146] * vector[98] +matrix[99][146] * vector[99] +b[146];
assign result[147] = matrix[0][147] * vector[0] +matrix[1][147] * vector[1] +matrix[2][147] * vector[2] +matrix[3][147] * vector[3] +matrix[4][147] * vector[4] +matrix[5][147] * vector[5] +matrix[6][147] * vector[6] +matrix[7][147] * vector[7] +matrix[8][147] * vector[8] +matrix[9][147] * vector[9] +matrix[10][147] * vector[10] +matrix[11][147] * vector[11] +matrix[12][147] * vector[12] +matrix[13][147] * vector[13] +matrix[14][147] * vector[14] +matrix[15][147] * vector[15] +matrix[16][147] * vector[16] +matrix[17][147] * vector[17] +matrix[18][147] * vector[18] +matrix[19][147] * vector[19] +matrix[20][147] * vector[20] +matrix[21][147] * vector[21] +matrix[22][147] * vector[22] +matrix[23][147] * vector[23] +matrix[24][147] * vector[24] +matrix[25][147] * vector[25] +matrix[26][147] * vector[26] +matrix[27][147] * vector[27] +matrix[28][147] * vector[28] +matrix[29][147] * vector[29] +matrix[30][147] * vector[30] +matrix[31][147] * vector[31] +matrix[32][147] * vector[32] +matrix[33][147] * vector[33] +matrix[34][147] * vector[34] +matrix[35][147] * vector[35] +matrix[36][147] * vector[36] +matrix[37][147] * vector[37] +matrix[38][147] * vector[38] +matrix[39][147] * vector[39] +matrix[40][147] * vector[40] +matrix[41][147] * vector[41] +matrix[42][147] * vector[42] +matrix[43][147] * vector[43] +matrix[44][147] * vector[44] +matrix[45][147] * vector[45] +matrix[46][147] * vector[46] +matrix[47][147] * vector[47] +matrix[48][147] * vector[48] +matrix[49][147] * vector[49] +matrix[50][147] * vector[50] +matrix[51][147] * vector[51] +matrix[52][147] * vector[52] +matrix[53][147] * vector[53] +matrix[54][147] * vector[54] +matrix[55][147] * vector[55] +matrix[56][147] * vector[56] +matrix[57][147] * vector[57] +matrix[58][147] * vector[58] +matrix[59][147] * vector[59] +matrix[60][147] * vector[60] +matrix[61][147] * vector[61] +matrix[62][147] * vector[62] +matrix[63][147] * vector[63] +matrix[64][147] * vector[64] +matrix[65][147] * vector[65] +matrix[66][147] * vector[66] +matrix[67][147] * vector[67] +matrix[68][147] * vector[68] +matrix[69][147] * vector[69] +matrix[70][147] * vector[70] +matrix[71][147] * vector[71] +matrix[72][147] * vector[72] +matrix[73][147] * vector[73] +matrix[74][147] * vector[74] +matrix[75][147] * vector[75] +matrix[76][147] * vector[76] +matrix[77][147] * vector[77] +matrix[78][147] * vector[78] +matrix[79][147] * vector[79] +matrix[80][147] * vector[80] +matrix[81][147] * vector[81] +matrix[82][147] * vector[82] +matrix[83][147] * vector[83] +matrix[84][147] * vector[84] +matrix[85][147] * vector[85] +matrix[86][147] * vector[86] +matrix[87][147] * vector[87] +matrix[88][147] * vector[88] +matrix[89][147] * vector[89] +matrix[90][147] * vector[90] +matrix[91][147] * vector[91] +matrix[92][147] * vector[92] +matrix[93][147] * vector[93] +matrix[94][147] * vector[94] +matrix[95][147] * vector[95] +matrix[96][147] * vector[96] +matrix[97][147] * vector[97] +matrix[98][147] * vector[98] +matrix[99][147] * vector[99] +b[147];
assign result[148] = matrix[0][148] * vector[0] +matrix[1][148] * vector[1] +matrix[2][148] * vector[2] +matrix[3][148] * vector[3] +matrix[4][148] * vector[4] +matrix[5][148] * vector[5] +matrix[6][148] * vector[6] +matrix[7][148] * vector[7] +matrix[8][148] * vector[8] +matrix[9][148] * vector[9] +matrix[10][148] * vector[10] +matrix[11][148] * vector[11] +matrix[12][148] * vector[12] +matrix[13][148] * vector[13] +matrix[14][148] * vector[14] +matrix[15][148] * vector[15] +matrix[16][148] * vector[16] +matrix[17][148] * vector[17] +matrix[18][148] * vector[18] +matrix[19][148] * vector[19] +matrix[20][148] * vector[20] +matrix[21][148] * vector[21] +matrix[22][148] * vector[22] +matrix[23][148] * vector[23] +matrix[24][148] * vector[24] +matrix[25][148] * vector[25] +matrix[26][148] * vector[26] +matrix[27][148] * vector[27] +matrix[28][148] * vector[28] +matrix[29][148] * vector[29] +matrix[30][148] * vector[30] +matrix[31][148] * vector[31] +matrix[32][148] * vector[32] +matrix[33][148] * vector[33] +matrix[34][148] * vector[34] +matrix[35][148] * vector[35] +matrix[36][148] * vector[36] +matrix[37][148] * vector[37] +matrix[38][148] * vector[38] +matrix[39][148] * vector[39] +matrix[40][148] * vector[40] +matrix[41][148] * vector[41] +matrix[42][148] * vector[42] +matrix[43][148] * vector[43] +matrix[44][148] * vector[44] +matrix[45][148] * vector[45] +matrix[46][148] * vector[46] +matrix[47][148] * vector[47] +matrix[48][148] * vector[48] +matrix[49][148] * vector[49] +matrix[50][148] * vector[50] +matrix[51][148] * vector[51] +matrix[52][148] * vector[52] +matrix[53][148] * vector[53] +matrix[54][148] * vector[54] +matrix[55][148] * vector[55] +matrix[56][148] * vector[56] +matrix[57][148] * vector[57] +matrix[58][148] * vector[58] +matrix[59][148] * vector[59] +matrix[60][148] * vector[60] +matrix[61][148] * vector[61] +matrix[62][148] * vector[62] +matrix[63][148] * vector[63] +matrix[64][148] * vector[64] +matrix[65][148] * vector[65] +matrix[66][148] * vector[66] +matrix[67][148] * vector[67] +matrix[68][148] * vector[68] +matrix[69][148] * vector[69] +matrix[70][148] * vector[70] +matrix[71][148] * vector[71] +matrix[72][148] * vector[72] +matrix[73][148] * vector[73] +matrix[74][148] * vector[74] +matrix[75][148] * vector[75] +matrix[76][148] * vector[76] +matrix[77][148] * vector[77] +matrix[78][148] * vector[78] +matrix[79][148] * vector[79] +matrix[80][148] * vector[80] +matrix[81][148] * vector[81] +matrix[82][148] * vector[82] +matrix[83][148] * vector[83] +matrix[84][148] * vector[84] +matrix[85][148] * vector[85] +matrix[86][148] * vector[86] +matrix[87][148] * vector[87] +matrix[88][148] * vector[88] +matrix[89][148] * vector[89] +matrix[90][148] * vector[90] +matrix[91][148] * vector[91] +matrix[92][148] * vector[92] +matrix[93][148] * vector[93] +matrix[94][148] * vector[94] +matrix[95][148] * vector[95] +matrix[96][148] * vector[96] +matrix[97][148] * vector[97] +matrix[98][148] * vector[98] +matrix[99][148] * vector[99] +b[148];
assign result[149] = matrix[0][149] * vector[0] +matrix[1][149] * vector[1] +matrix[2][149] * vector[2] +matrix[3][149] * vector[3] +matrix[4][149] * vector[4] +matrix[5][149] * vector[5] +matrix[6][149] * vector[6] +matrix[7][149] * vector[7] +matrix[8][149] * vector[8] +matrix[9][149] * vector[9] +matrix[10][149] * vector[10] +matrix[11][149] * vector[11] +matrix[12][149] * vector[12] +matrix[13][149] * vector[13] +matrix[14][149] * vector[14] +matrix[15][149] * vector[15] +matrix[16][149] * vector[16] +matrix[17][149] * vector[17] +matrix[18][149] * vector[18] +matrix[19][149] * vector[19] +matrix[20][149] * vector[20] +matrix[21][149] * vector[21] +matrix[22][149] * vector[22] +matrix[23][149] * vector[23] +matrix[24][149] * vector[24] +matrix[25][149] * vector[25] +matrix[26][149] * vector[26] +matrix[27][149] * vector[27] +matrix[28][149] * vector[28] +matrix[29][149] * vector[29] +matrix[30][149] * vector[30] +matrix[31][149] * vector[31] +matrix[32][149] * vector[32] +matrix[33][149] * vector[33] +matrix[34][149] * vector[34] +matrix[35][149] * vector[35] +matrix[36][149] * vector[36] +matrix[37][149] * vector[37] +matrix[38][149] * vector[38] +matrix[39][149] * vector[39] +matrix[40][149] * vector[40] +matrix[41][149] * vector[41] +matrix[42][149] * vector[42] +matrix[43][149] * vector[43] +matrix[44][149] * vector[44] +matrix[45][149] * vector[45] +matrix[46][149] * vector[46] +matrix[47][149] * vector[47] +matrix[48][149] * vector[48] +matrix[49][149] * vector[49] +matrix[50][149] * vector[50] +matrix[51][149] * vector[51] +matrix[52][149] * vector[52] +matrix[53][149] * vector[53] +matrix[54][149] * vector[54] +matrix[55][149] * vector[55] +matrix[56][149] * vector[56] +matrix[57][149] * vector[57] +matrix[58][149] * vector[58] +matrix[59][149] * vector[59] +matrix[60][149] * vector[60] +matrix[61][149] * vector[61] +matrix[62][149] * vector[62] +matrix[63][149] * vector[63] +matrix[64][149] * vector[64] +matrix[65][149] * vector[65] +matrix[66][149] * vector[66] +matrix[67][149] * vector[67] +matrix[68][149] * vector[68] +matrix[69][149] * vector[69] +matrix[70][149] * vector[70] +matrix[71][149] * vector[71] +matrix[72][149] * vector[72] +matrix[73][149] * vector[73] +matrix[74][149] * vector[74] +matrix[75][149] * vector[75] +matrix[76][149] * vector[76] +matrix[77][149] * vector[77] +matrix[78][149] * vector[78] +matrix[79][149] * vector[79] +matrix[80][149] * vector[80] +matrix[81][149] * vector[81] +matrix[82][149] * vector[82] +matrix[83][149] * vector[83] +matrix[84][149] * vector[84] +matrix[85][149] * vector[85] +matrix[86][149] * vector[86] +matrix[87][149] * vector[87] +matrix[88][149] * vector[88] +matrix[89][149] * vector[89] +matrix[90][149] * vector[90] +matrix[91][149] * vector[91] +matrix[92][149] * vector[92] +matrix[93][149] * vector[93] +matrix[94][149] * vector[94] +matrix[95][149] * vector[95] +matrix[96][149] * vector[96] +matrix[97][149] * vector[97] +matrix[98][149] * vector[98] +matrix[99][149] * vector[99] +b[149];
assign result[150] = matrix[0][150] * vector[0] +matrix[1][150] * vector[1] +matrix[2][150] * vector[2] +matrix[3][150] * vector[3] +matrix[4][150] * vector[4] +matrix[5][150] * vector[5] +matrix[6][150] * vector[6] +matrix[7][150] * vector[7] +matrix[8][150] * vector[8] +matrix[9][150] * vector[9] +matrix[10][150] * vector[10] +matrix[11][150] * vector[11] +matrix[12][150] * vector[12] +matrix[13][150] * vector[13] +matrix[14][150] * vector[14] +matrix[15][150] * vector[15] +matrix[16][150] * vector[16] +matrix[17][150] * vector[17] +matrix[18][150] * vector[18] +matrix[19][150] * vector[19] +matrix[20][150] * vector[20] +matrix[21][150] * vector[21] +matrix[22][150] * vector[22] +matrix[23][150] * vector[23] +matrix[24][150] * vector[24] +matrix[25][150] * vector[25] +matrix[26][150] * vector[26] +matrix[27][150] * vector[27] +matrix[28][150] * vector[28] +matrix[29][150] * vector[29] +matrix[30][150] * vector[30] +matrix[31][150] * vector[31] +matrix[32][150] * vector[32] +matrix[33][150] * vector[33] +matrix[34][150] * vector[34] +matrix[35][150] * vector[35] +matrix[36][150] * vector[36] +matrix[37][150] * vector[37] +matrix[38][150] * vector[38] +matrix[39][150] * vector[39] +matrix[40][150] * vector[40] +matrix[41][150] * vector[41] +matrix[42][150] * vector[42] +matrix[43][150] * vector[43] +matrix[44][150] * vector[44] +matrix[45][150] * vector[45] +matrix[46][150] * vector[46] +matrix[47][150] * vector[47] +matrix[48][150] * vector[48] +matrix[49][150] * vector[49] +matrix[50][150] * vector[50] +matrix[51][150] * vector[51] +matrix[52][150] * vector[52] +matrix[53][150] * vector[53] +matrix[54][150] * vector[54] +matrix[55][150] * vector[55] +matrix[56][150] * vector[56] +matrix[57][150] * vector[57] +matrix[58][150] * vector[58] +matrix[59][150] * vector[59] +matrix[60][150] * vector[60] +matrix[61][150] * vector[61] +matrix[62][150] * vector[62] +matrix[63][150] * vector[63] +matrix[64][150] * vector[64] +matrix[65][150] * vector[65] +matrix[66][150] * vector[66] +matrix[67][150] * vector[67] +matrix[68][150] * vector[68] +matrix[69][150] * vector[69] +matrix[70][150] * vector[70] +matrix[71][150] * vector[71] +matrix[72][150] * vector[72] +matrix[73][150] * vector[73] +matrix[74][150] * vector[74] +matrix[75][150] * vector[75] +matrix[76][150] * vector[76] +matrix[77][150] * vector[77] +matrix[78][150] * vector[78] +matrix[79][150] * vector[79] +matrix[80][150] * vector[80] +matrix[81][150] * vector[81] +matrix[82][150] * vector[82] +matrix[83][150] * vector[83] +matrix[84][150] * vector[84] +matrix[85][150] * vector[85] +matrix[86][150] * vector[86] +matrix[87][150] * vector[87] +matrix[88][150] * vector[88] +matrix[89][150] * vector[89] +matrix[90][150] * vector[90] +matrix[91][150] * vector[91] +matrix[92][150] * vector[92] +matrix[93][150] * vector[93] +matrix[94][150] * vector[94] +matrix[95][150] * vector[95] +matrix[96][150] * vector[96] +matrix[97][150] * vector[97] +matrix[98][150] * vector[98] +matrix[99][150] * vector[99] +b[150];
assign result[151] = matrix[0][151] * vector[0] +matrix[1][151] * vector[1] +matrix[2][151] * vector[2] +matrix[3][151] * vector[3] +matrix[4][151] * vector[4] +matrix[5][151] * vector[5] +matrix[6][151] * vector[6] +matrix[7][151] * vector[7] +matrix[8][151] * vector[8] +matrix[9][151] * vector[9] +matrix[10][151] * vector[10] +matrix[11][151] * vector[11] +matrix[12][151] * vector[12] +matrix[13][151] * vector[13] +matrix[14][151] * vector[14] +matrix[15][151] * vector[15] +matrix[16][151] * vector[16] +matrix[17][151] * vector[17] +matrix[18][151] * vector[18] +matrix[19][151] * vector[19] +matrix[20][151] * vector[20] +matrix[21][151] * vector[21] +matrix[22][151] * vector[22] +matrix[23][151] * vector[23] +matrix[24][151] * vector[24] +matrix[25][151] * vector[25] +matrix[26][151] * vector[26] +matrix[27][151] * vector[27] +matrix[28][151] * vector[28] +matrix[29][151] * vector[29] +matrix[30][151] * vector[30] +matrix[31][151] * vector[31] +matrix[32][151] * vector[32] +matrix[33][151] * vector[33] +matrix[34][151] * vector[34] +matrix[35][151] * vector[35] +matrix[36][151] * vector[36] +matrix[37][151] * vector[37] +matrix[38][151] * vector[38] +matrix[39][151] * vector[39] +matrix[40][151] * vector[40] +matrix[41][151] * vector[41] +matrix[42][151] * vector[42] +matrix[43][151] * vector[43] +matrix[44][151] * vector[44] +matrix[45][151] * vector[45] +matrix[46][151] * vector[46] +matrix[47][151] * vector[47] +matrix[48][151] * vector[48] +matrix[49][151] * vector[49] +matrix[50][151] * vector[50] +matrix[51][151] * vector[51] +matrix[52][151] * vector[52] +matrix[53][151] * vector[53] +matrix[54][151] * vector[54] +matrix[55][151] * vector[55] +matrix[56][151] * vector[56] +matrix[57][151] * vector[57] +matrix[58][151] * vector[58] +matrix[59][151] * vector[59] +matrix[60][151] * vector[60] +matrix[61][151] * vector[61] +matrix[62][151] * vector[62] +matrix[63][151] * vector[63] +matrix[64][151] * vector[64] +matrix[65][151] * vector[65] +matrix[66][151] * vector[66] +matrix[67][151] * vector[67] +matrix[68][151] * vector[68] +matrix[69][151] * vector[69] +matrix[70][151] * vector[70] +matrix[71][151] * vector[71] +matrix[72][151] * vector[72] +matrix[73][151] * vector[73] +matrix[74][151] * vector[74] +matrix[75][151] * vector[75] +matrix[76][151] * vector[76] +matrix[77][151] * vector[77] +matrix[78][151] * vector[78] +matrix[79][151] * vector[79] +matrix[80][151] * vector[80] +matrix[81][151] * vector[81] +matrix[82][151] * vector[82] +matrix[83][151] * vector[83] +matrix[84][151] * vector[84] +matrix[85][151] * vector[85] +matrix[86][151] * vector[86] +matrix[87][151] * vector[87] +matrix[88][151] * vector[88] +matrix[89][151] * vector[89] +matrix[90][151] * vector[90] +matrix[91][151] * vector[91] +matrix[92][151] * vector[92] +matrix[93][151] * vector[93] +matrix[94][151] * vector[94] +matrix[95][151] * vector[95] +matrix[96][151] * vector[96] +matrix[97][151] * vector[97] +matrix[98][151] * vector[98] +matrix[99][151] * vector[99] +b[151];
assign result[152] = matrix[0][152] * vector[0] +matrix[1][152] * vector[1] +matrix[2][152] * vector[2] +matrix[3][152] * vector[3] +matrix[4][152] * vector[4] +matrix[5][152] * vector[5] +matrix[6][152] * vector[6] +matrix[7][152] * vector[7] +matrix[8][152] * vector[8] +matrix[9][152] * vector[9] +matrix[10][152] * vector[10] +matrix[11][152] * vector[11] +matrix[12][152] * vector[12] +matrix[13][152] * vector[13] +matrix[14][152] * vector[14] +matrix[15][152] * vector[15] +matrix[16][152] * vector[16] +matrix[17][152] * vector[17] +matrix[18][152] * vector[18] +matrix[19][152] * vector[19] +matrix[20][152] * vector[20] +matrix[21][152] * vector[21] +matrix[22][152] * vector[22] +matrix[23][152] * vector[23] +matrix[24][152] * vector[24] +matrix[25][152] * vector[25] +matrix[26][152] * vector[26] +matrix[27][152] * vector[27] +matrix[28][152] * vector[28] +matrix[29][152] * vector[29] +matrix[30][152] * vector[30] +matrix[31][152] * vector[31] +matrix[32][152] * vector[32] +matrix[33][152] * vector[33] +matrix[34][152] * vector[34] +matrix[35][152] * vector[35] +matrix[36][152] * vector[36] +matrix[37][152] * vector[37] +matrix[38][152] * vector[38] +matrix[39][152] * vector[39] +matrix[40][152] * vector[40] +matrix[41][152] * vector[41] +matrix[42][152] * vector[42] +matrix[43][152] * vector[43] +matrix[44][152] * vector[44] +matrix[45][152] * vector[45] +matrix[46][152] * vector[46] +matrix[47][152] * vector[47] +matrix[48][152] * vector[48] +matrix[49][152] * vector[49] +matrix[50][152] * vector[50] +matrix[51][152] * vector[51] +matrix[52][152] * vector[52] +matrix[53][152] * vector[53] +matrix[54][152] * vector[54] +matrix[55][152] * vector[55] +matrix[56][152] * vector[56] +matrix[57][152] * vector[57] +matrix[58][152] * vector[58] +matrix[59][152] * vector[59] +matrix[60][152] * vector[60] +matrix[61][152] * vector[61] +matrix[62][152] * vector[62] +matrix[63][152] * vector[63] +matrix[64][152] * vector[64] +matrix[65][152] * vector[65] +matrix[66][152] * vector[66] +matrix[67][152] * vector[67] +matrix[68][152] * vector[68] +matrix[69][152] * vector[69] +matrix[70][152] * vector[70] +matrix[71][152] * vector[71] +matrix[72][152] * vector[72] +matrix[73][152] * vector[73] +matrix[74][152] * vector[74] +matrix[75][152] * vector[75] +matrix[76][152] * vector[76] +matrix[77][152] * vector[77] +matrix[78][152] * vector[78] +matrix[79][152] * vector[79] +matrix[80][152] * vector[80] +matrix[81][152] * vector[81] +matrix[82][152] * vector[82] +matrix[83][152] * vector[83] +matrix[84][152] * vector[84] +matrix[85][152] * vector[85] +matrix[86][152] * vector[86] +matrix[87][152] * vector[87] +matrix[88][152] * vector[88] +matrix[89][152] * vector[89] +matrix[90][152] * vector[90] +matrix[91][152] * vector[91] +matrix[92][152] * vector[92] +matrix[93][152] * vector[93] +matrix[94][152] * vector[94] +matrix[95][152] * vector[95] +matrix[96][152] * vector[96] +matrix[97][152] * vector[97] +matrix[98][152] * vector[98] +matrix[99][152] * vector[99] +b[152];
assign result[153] = matrix[0][153] * vector[0] +matrix[1][153] * vector[1] +matrix[2][153] * vector[2] +matrix[3][153] * vector[3] +matrix[4][153] * vector[4] +matrix[5][153] * vector[5] +matrix[6][153] * vector[6] +matrix[7][153] * vector[7] +matrix[8][153] * vector[8] +matrix[9][153] * vector[9] +matrix[10][153] * vector[10] +matrix[11][153] * vector[11] +matrix[12][153] * vector[12] +matrix[13][153] * vector[13] +matrix[14][153] * vector[14] +matrix[15][153] * vector[15] +matrix[16][153] * vector[16] +matrix[17][153] * vector[17] +matrix[18][153] * vector[18] +matrix[19][153] * vector[19] +matrix[20][153] * vector[20] +matrix[21][153] * vector[21] +matrix[22][153] * vector[22] +matrix[23][153] * vector[23] +matrix[24][153] * vector[24] +matrix[25][153] * vector[25] +matrix[26][153] * vector[26] +matrix[27][153] * vector[27] +matrix[28][153] * vector[28] +matrix[29][153] * vector[29] +matrix[30][153] * vector[30] +matrix[31][153] * vector[31] +matrix[32][153] * vector[32] +matrix[33][153] * vector[33] +matrix[34][153] * vector[34] +matrix[35][153] * vector[35] +matrix[36][153] * vector[36] +matrix[37][153] * vector[37] +matrix[38][153] * vector[38] +matrix[39][153] * vector[39] +matrix[40][153] * vector[40] +matrix[41][153] * vector[41] +matrix[42][153] * vector[42] +matrix[43][153] * vector[43] +matrix[44][153] * vector[44] +matrix[45][153] * vector[45] +matrix[46][153] * vector[46] +matrix[47][153] * vector[47] +matrix[48][153] * vector[48] +matrix[49][153] * vector[49] +matrix[50][153] * vector[50] +matrix[51][153] * vector[51] +matrix[52][153] * vector[52] +matrix[53][153] * vector[53] +matrix[54][153] * vector[54] +matrix[55][153] * vector[55] +matrix[56][153] * vector[56] +matrix[57][153] * vector[57] +matrix[58][153] * vector[58] +matrix[59][153] * vector[59] +matrix[60][153] * vector[60] +matrix[61][153] * vector[61] +matrix[62][153] * vector[62] +matrix[63][153] * vector[63] +matrix[64][153] * vector[64] +matrix[65][153] * vector[65] +matrix[66][153] * vector[66] +matrix[67][153] * vector[67] +matrix[68][153] * vector[68] +matrix[69][153] * vector[69] +matrix[70][153] * vector[70] +matrix[71][153] * vector[71] +matrix[72][153] * vector[72] +matrix[73][153] * vector[73] +matrix[74][153] * vector[74] +matrix[75][153] * vector[75] +matrix[76][153] * vector[76] +matrix[77][153] * vector[77] +matrix[78][153] * vector[78] +matrix[79][153] * vector[79] +matrix[80][153] * vector[80] +matrix[81][153] * vector[81] +matrix[82][153] * vector[82] +matrix[83][153] * vector[83] +matrix[84][153] * vector[84] +matrix[85][153] * vector[85] +matrix[86][153] * vector[86] +matrix[87][153] * vector[87] +matrix[88][153] * vector[88] +matrix[89][153] * vector[89] +matrix[90][153] * vector[90] +matrix[91][153] * vector[91] +matrix[92][153] * vector[92] +matrix[93][153] * vector[93] +matrix[94][153] * vector[94] +matrix[95][153] * vector[95] +matrix[96][153] * vector[96] +matrix[97][153] * vector[97] +matrix[98][153] * vector[98] +matrix[99][153] * vector[99] +b[153];
assign result[154] = matrix[0][154] * vector[0] +matrix[1][154] * vector[1] +matrix[2][154] * vector[2] +matrix[3][154] * vector[3] +matrix[4][154] * vector[4] +matrix[5][154] * vector[5] +matrix[6][154] * vector[6] +matrix[7][154] * vector[7] +matrix[8][154] * vector[8] +matrix[9][154] * vector[9] +matrix[10][154] * vector[10] +matrix[11][154] * vector[11] +matrix[12][154] * vector[12] +matrix[13][154] * vector[13] +matrix[14][154] * vector[14] +matrix[15][154] * vector[15] +matrix[16][154] * vector[16] +matrix[17][154] * vector[17] +matrix[18][154] * vector[18] +matrix[19][154] * vector[19] +matrix[20][154] * vector[20] +matrix[21][154] * vector[21] +matrix[22][154] * vector[22] +matrix[23][154] * vector[23] +matrix[24][154] * vector[24] +matrix[25][154] * vector[25] +matrix[26][154] * vector[26] +matrix[27][154] * vector[27] +matrix[28][154] * vector[28] +matrix[29][154] * vector[29] +matrix[30][154] * vector[30] +matrix[31][154] * vector[31] +matrix[32][154] * vector[32] +matrix[33][154] * vector[33] +matrix[34][154] * vector[34] +matrix[35][154] * vector[35] +matrix[36][154] * vector[36] +matrix[37][154] * vector[37] +matrix[38][154] * vector[38] +matrix[39][154] * vector[39] +matrix[40][154] * vector[40] +matrix[41][154] * vector[41] +matrix[42][154] * vector[42] +matrix[43][154] * vector[43] +matrix[44][154] * vector[44] +matrix[45][154] * vector[45] +matrix[46][154] * vector[46] +matrix[47][154] * vector[47] +matrix[48][154] * vector[48] +matrix[49][154] * vector[49] +matrix[50][154] * vector[50] +matrix[51][154] * vector[51] +matrix[52][154] * vector[52] +matrix[53][154] * vector[53] +matrix[54][154] * vector[54] +matrix[55][154] * vector[55] +matrix[56][154] * vector[56] +matrix[57][154] * vector[57] +matrix[58][154] * vector[58] +matrix[59][154] * vector[59] +matrix[60][154] * vector[60] +matrix[61][154] * vector[61] +matrix[62][154] * vector[62] +matrix[63][154] * vector[63] +matrix[64][154] * vector[64] +matrix[65][154] * vector[65] +matrix[66][154] * vector[66] +matrix[67][154] * vector[67] +matrix[68][154] * vector[68] +matrix[69][154] * vector[69] +matrix[70][154] * vector[70] +matrix[71][154] * vector[71] +matrix[72][154] * vector[72] +matrix[73][154] * vector[73] +matrix[74][154] * vector[74] +matrix[75][154] * vector[75] +matrix[76][154] * vector[76] +matrix[77][154] * vector[77] +matrix[78][154] * vector[78] +matrix[79][154] * vector[79] +matrix[80][154] * vector[80] +matrix[81][154] * vector[81] +matrix[82][154] * vector[82] +matrix[83][154] * vector[83] +matrix[84][154] * vector[84] +matrix[85][154] * vector[85] +matrix[86][154] * vector[86] +matrix[87][154] * vector[87] +matrix[88][154] * vector[88] +matrix[89][154] * vector[89] +matrix[90][154] * vector[90] +matrix[91][154] * vector[91] +matrix[92][154] * vector[92] +matrix[93][154] * vector[93] +matrix[94][154] * vector[94] +matrix[95][154] * vector[95] +matrix[96][154] * vector[96] +matrix[97][154] * vector[97] +matrix[98][154] * vector[98] +matrix[99][154] * vector[99] +b[154];
assign result[155] = matrix[0][155] * vector[0] +matrix[1][155] * vector[1] +matrix[2][155] * vector[2] +matrix[3][155] * vector[3] +matrix[4][155] * vector[4] +matrix[5][155] * vector[5] +matrix[6][155] * vector[6] +matrix[7][155] * vector[7] +matrix[8][155] * vector[8] +matrix[9][155] * vector[9] +matrix[10][155] * vector[10] +matrix[11][155] * vector[11] +matrix[12][155] * vector[12] +matrix[13][155] * vector[13] +matrix[14][155] * vector[14] +matrix[15][155] * vector[15] +matrix[16][155] * vector[16] +matrix[17][155] * vector[17] +matrix[18][155] * vector[18] +matrix[19][155] * vector[19] +matrix[20][155] * vector[20] +matrix[21][155] * vector[21] +matrix[22][155] * vector[22] +matrix[23][155] * vector[23] +matrix[24][155] * vector[24] +matrix[25][155] * vector[25] +matrix[26][155] * vector[26] +matrix[27][155] * vector[27] +matrix[28][155] * vector[28] +matrix[29][155] * vector[29] +matrix[30][155] * vector[30] +matrix[31][155] * vector[31] +matrix[32][155] * vector[32] +matrix[33][155] * vector[33] +matrix[34][155] * vector[34] +matrix[35][155] * vector[35] +matrix[36][155] * vector[36] +matrix[37][155] * vector[37] +matrix[38][155] * vector[38] +matrix[39][155] * vector[39] +matrix[40][155] * vector[40] +matrix[41][155] * vector[41] +matrix[42][155] * vector[42] +matrix[43][155] * vector[43] +matrix[44][155] * vector[44] +matrix[45][155] * vector[45] +matrix[46][155] * vector[46] +matrix[47][155] * vector[47] +matrix[48][155] * vector[48] +matrix[49][155] * vector[49] +matrix[50][155] * vector[50] +matrix[51][155] * vector[51] +matrix[52][155] * vector[52] +matrix[53][155] * vector[53] +matrix[54][155] * vector[54] +matrix[55][155] * vector[55] +matrix[56][155] * vector[56] +matrix[57][155] * vector[57] +matrix[58][155] * vector[58] +matrix[59][155] * vector[59] +matrix[60][155] * vector[60] +matrix[61][155] * vector[61] +matrix[62][155] * vector[62] +matrix[63][155] * vector[63] +matrix[64][155] * vector[64] +matrix[65][155] * vector[65] +matrix[66][155] * vector[66] +matrix[67][155] * vector[67] +matrix[68][155] * vector[68] +matrix[69][155] * vector[69] +matrix[70][155] * vector[70] +matrix[71][155] * vector[71] +matrix[72][155] * vector[72] +matrix[73][155] * vector[73] +matrix[74][155] * vector[74] +matrix[75][155] * vector[75] +matrix[76][155] * vector[76] +matrix[77][155] * vector[77] +matrix[78][155] * vector[78] +matrix[79][155] * vector[79] +matrix[80][155] * vector[80] +matrix[81][155] * vector[81] +matrix[82][155] * vector[82] +matrix[83][155] * vector[83] +matrix[84][155] * vector[84] +matrix[85][155] * vector[85] +matrix[86][155] * vector[86] +matrix[87][155] * vector[87] +matrix[88][155] * vector[88] +matrix[89][155] * vector[89] +matrix[90][155] * vector[90] +matrix[91][155] * vector[91] +matrix[92][155] * vector[92] +matrix[93][155] * vector[93] +matrix[94][155] * vector[94] +matrix[95][155] * vector[95] +matrix[96][155] * vector[96] +matrix[97][155] * vector[97] +matrix[98][155] * vector[98] +matrix[99][155] * vector[99] +b[155];
assign result[156] = matrix[0][156] * vector[0] +matrix[1][156] * vector[1] +matrix[2][156] * vector[2] +matrix[3][156] * vector[3] +matrix[4][156] * vector[4] +matrix[5][156] * vector[5] +matrix[6][156] * vector[6] +matrix[7][156] * vector[7] +matrix[8][156] * vector[8] +matrix[9][156] * vector[9] +matrix[10][156] * vector[10] +matrix[11][156] * vector[11] +matrix[12][156] * vector[12] +matrix[13][156] * vector[13] +matrix[14][156] * vector[14] +matrix[15][156] * vector[15] +matrix[16][156] * vector[16] +matrix[17][156] * vector[17] +matrix[18][156] * vector[18] +matrix[19][156] * vector[19] +matrix[20][156] * vector[20] +matrix[21][156] * vector[21] +matrix[22][156] * vector[22] +matrix[23][156] * vector[23] +matrix[24][156] * vector[24] +matrix[25][156] * vector[25] +matrix[26][156] * vector[26] +matrix[27][156] * vector[27] +matrix[28][156] * vector[28] +matrix[29][156] * vector[29] +matrix[30][156] * vector[30] +matrix[31][156] * vector[31] +matrix[32][156] * vector[32] +matrix[33][156] * vector[33] +matrix[34][156] * vector[34] +matrix[35][156] * vector[35] +matrix[36][156] * vector[36] +matrix[37][156] * vector[37] +matrix[38][156] * vector[38] +matrix[39][156] * vector[39] +matrix[40][156] * vector[40] +matrix[41][156] * vector[41] +matrix[42][156] * vector[42] +matrix[43][156] * vector[43] +matrix[44][156] * vector[44] +matrix[45][156] * vector[45] +matrix[46][156] * vector[46] +matrix[47][156] * vector[47] +matrix[48][156] * vector[48] +matrix[49][156] * vector[49] +matrix[50][156] * vector[50] +matrix[51][156] * vector[51] +matrix[52][156] * vector[52] +matrix[53][156] * vector[53] +matrix[54][156] * vector[54] +matrix[55][156] * vector[55] +matrix[56][156] * vector[56] +matrix[57][156] * vector[57] +matrix[58][156] * vector[58] +matrix[59][156] * vector[59] +matrix[60][156] * vector[60] +matrix[61][156] * vector[61] +matrix[62][156] * vector[62] +matrix[63][156] * vector[63] +matrix[64][156] * vector[64] +matrix[65][156] * vector[65] +matrix[66][156] * vector[66] +matrix[67][156] * vector[67] +matrix[68][156] * vector[68] +matrix[69][156] * vector[69] +matrix[70][156] * vector[70] +matrix[71][156] * vector[71] +matrix[72][156] * vector[72] +matrix[73][156] * vector[73] +matrix[74][156] * vector[74] +matrix[75][156] * vector[75] +matrix[76][156] * vector[76] +matrix[77][156] * vector[77] +matrix[78][156] * vector[78] +matrix[79][156] * vector[79] +matrix[80][156] * vector[80] +matrix[81][156] * vector[81] +matrix[82][156] * vector[82] +matrix[83][156] * vector[83] +matrix[84][156] * vector[84] +matrix[85][156] * vector[85] +matrix[86][156] * vector[86] +matrix[87][156] * vector[87] +matrix[88][156] * vector[88] +matrix[89][156] * vector[89] +matrix[90][156] * vector[90] +matrix[91][156] * vector[91] +matrix[92][156] * vector[92] +matrix[93][156] * vector[93] +matrix[94][156] * vector[94] +matrix[95][156] * vector[95] +matrix[96][156] * vector[96] +matrix[97][156] * vector[97] +matrix[98][156] * vector[98] +matrix[99][156] * vector[99] +b[156];
assign result[157] = matrix[0][157] * vector[0] +matrix[1][157] * vector[1] +matrix[2][157] * vector[2] +matrix[3][157] * vector[3] +matrix[4][157] * vector[4] +matrix[5][157] * vector[5] +matrix[6][157] * vector[6] +matrix[7][157] * vector[7] +matrix[8][157] * vector[8] +matrix[9][157] * vector[9] +matrix[10][157] * vector[10] +matrix[11][157] * vector[11] +matrix[12][157] * vector[12] +matrix[13][157] * vector[13] +matrix[14][157] * vector[14] +matrix[15][157] * vector[15] +matrix[16][157] * vector[16] +matrix[17][157] * vector[17] +matrix[18][157] * vector[18] +matrix[19][157] * vector[19] +matrix[20][157] * vector[20] +matrix[21][157] * vector[21] +matrix[22][157] * vector[22] +matrix[23][157] * vector[23] +matrix[24][157] * vector[24] +matrix[25][157] * vector[25] +matrix[26][157] * vector[26] +matrix[27][157] * vector[27] +matrix[28][157] * vector[28] +matrix[29][157] * vector[29] +matrix[30][157] * vector[30] +matrix[31][157] * vector[31] +matrix[32][157] * vector[32] +matrix[33][157] * vector[33] +matrix[34][157] * vector[34] +matrix[35][157] * vector[35] +matrix[36][157] * vector[36] +matrix[37][157] * vector[37] +matrix[38][157] * vector[38] +matrix[39][157] * vector[39] +matrix[40][157] * vector[40] +matrix[41][157] * vector[41] +matrix[42][157] * vector[42] +matrix[43][157] * vector[43] +matrix[44][157] * vector[44] +matrix[45][157] * vector[45] +matrix[46][157] * vector[46] +matrix[47][157] * vector[47] +matrix[48][157] * vector[48] +matrix[49][157] * vector[49] +matrix[50][157] * vector[50] +matrix[51][157] * vector[51] +matrix[52][157] * vector[52] +matrix[53][157] * vector[53] +matrix[54][157] * vector[54] +matrix[55][157] * vector[55] +matrix[56][157] * vector[56] +matrix[57][157] * vector[57] +matrix[58][157] * vector[58] +matrix[59][157] * vector[59] +matrix[60][157] * vector[60] +matrix[61][157] * vector[61] +matrix[62][157] * vector[62] +matrix[63][157] * vector[63] +matrix[64][157] * vector[64] +matrix[65][157] * vector[65] +matrix[66][157] * vector[66] +matrix[67][157] * vector[67] +matrix[68][157] * vector[68] +matrix[69][157] * vector[69] +matrix[70][157] * vector[70] +matrix[71][157] * vector[71] +matrix[72][157] * vector[72] +matrix[73][157] * vector[73] +matrix[74][157] * vector[74] +matrix[75][157] * vector[75] +matrix[76][157] * vector[76] +matrix[77][157] * vector[77] +matrix[78][157] * vector[78] +matrix[79][157] * vector[79] +matrix[80][157] * vector[80] +matrix[81][157] * vector[81] +matrix[82][157] * vector[82] +matrix[83][157] * vector[83] +matrix[84][157] * vector[84] +matrix[85][157] * vector[85] +matrix[86][157] * vector[86] +matrix[87][157] * vector[87] +matrix[88][157] * vector[88] +matrix[89][157] * vector[89] +matrix[90][157] * vector[90] +matrix[91][157] * vector[91] +matrix[92][157] * vector[92] +matrix[93][157] * vector[93] +matrix[94][157] * vector[94] +matrix[95][157] * vector[95] +matrix[96][157] * vector[96] +matrix[97][157] * vector[97] +matrix[98][157] * vector[98] +matrix[99][157] * vector[99] +b[157];
assign result[158] = matrix[0][158] * vector[0] +matrix[1][158] * vector[1] +matrix[2][158] * vector[2] +matrix[3][158] * vector[3] +matrix[4][158] * vector[4] +matrix[5][158] * vector[5] +matrix[6][158] * vector[6] +matrix[7][158] * vector[7] +matrix[8][158] * vector[8] +matrix[9][158] * vector[9] +matrix[10][158] * vector[10] +matrix[11][158] * vector[11] +matrix[12][158] * vector[12] +matrix[13][158] * vector[13] +matrix[14][158] * vector[14] +matrix[15][158] * vector[15] +matrix[16][158] * vector[16] +matrix[17][158] * vector[17] +matrix[18][158] * vector[18] +matrix[19][158] * vector[19] +matrix[20][158] * vector[20] +matrix[21][158] * vector[21] +matrix[22][158] * vector[22] +matrix[23][158] * vector[23] +matrix[24][158] * vector[24] +matrix[25][158] * vector[25] +matrix[26][158] * vector[26] +matrix[27][158] * vector[27] +matrix[28][158] * vector[28] +matrix[29][158] * vector[29] +matrix[30][158] * vector[30] +matrix[31][158] * vector[31] +matrix[32][158] * vector[32] +matrix[33][158] * vector[33] +matrix[34][158] * vector[34] +matrix[35][158] * vector[35] +matrix[36][158] * vector[36] +matrix[37][158] * vector[37] +matrix[38][158] * vector[38] +matrix[39][158] * vector[39] +matrix[40][158] * vector[40] +matrix[41][158] * vector[41] +matrix[42][158] * vector[42] +matrix[43][158] * vector[43] +matrix[44][158] * vector[44] +matrix[45][158] * vector[45] +matrix[46][158] * vector[46] +matrix[47][158] * vector[47] +matrix[48][158] * vector[48] +matrix[49][158] * vector[49] +matrix[50][158] * vector[50] +matrix[51][158] * vector[51] +matrix[52][158] * vector[52] +matrix[53][158] * vector[53] +matrix[54][158] * vector[54] +matrix[55][158] * vector[55] +matrix[56][158] * vector[56] +matrix[57][158] * vector[57] +matrix[58][158] * vector[58] +matrix[59][158] * vector[59] +matrix[60][158] * vector[60] +matrix[61][158] * vector[61] +matrix[62][158] * vector[62] +matrix[63][158] * vector[63] +matrix[64][158] * vector[64] +matrix[65][158] * vector[65] +matrix[66][158] * vector[66] +matrix[67][158] * vector[67] +matrix[68][158] * vector[68] +matrix[69][158] * vector[69] +matrix[70][158] * vector[70] +matrix[71][158] * vector[71] +matrix[72][158] * vector[72] +matrix[73][158] * vector[73] +matrix[74][158] * vector[74] +matrix[75][158] * vector[75] +matrix[76][158] * vector[76] +matrix[77][158] * vector[77] +matrix[78][158] * vector[78] +matrix[79][158] * vector[79] +matrix[80][158] * vector[80] +matrix[81][158] * vector[81] +matrix[82][158] * vector[82] +matrix[83][158] * vector[83] +matrix[84][158] * vector[84] +matrix[85][158] * vector[85] +matrix[86][158] * vector[86] +matrix[87][158] * vector[87] +matrix[88][158] * vector[88] +matrix[89][158] * vector[89] +matrix[90][158] * vector[90] +matrix[91][158] * vector[91] +matrix[92][158] * vector[92] +matrix[93][158] * vector[93] +matrix[94][158] * vector[94] +matrix[95][158] * vector[95] +matrix[96][158] * vector[96] +matrix[97][158] * vector[97] +matrix[98][158] * vector[98] +matrix[99][158] * vector[99] +b[158];
assign result[159] = matrix[0][159] * vector[0] +matrix[1][159] * vector[1] +matrix[2][159] * vector[2] +matrix[3][159] * vector[3] +matrix[4][159] * vector[4] +matrix[5][159] * vector[5] +matrix[6][159] * vector[6] +matrix[7][159] * vector[7] +matrix[8][159] * vector[8] +matrix[9][159] * vector[9] +matrix[10][159] * vector[10] +matrix[11][159] * vector[11] +matrix[12][159] * vector[12] +matrix[13][159] * vector[13] +matrix[14][159] * vector[14] +matrix[15][159] * vector[15] +matrix[16][159] * vector[16] +matrix[17][159] * vector[17] +matrix[18][159] * vector[18] +matrix[19][159] * vector[19] +matrix[20][159] * vector[20] +matrix[21][159] * vector[21] +matrix[22][159] * vector[22] +matrix[23][159] * vector[23] +matrix[24][159] * vector[24] +matrix[25][159] * vector[25] +matrix[26][159] * vector[26] +matrix[27][159] * vector[27] +matrix[28][159] * vector[28] +matrix[29][159] * vector[29] +matrix[30][159] * vector[30] +matrix[31][159] * vector[31] +matrix[32][159] * vector[32] +matrix[33][159] * vector[33] +matrix[34][159] * vector[34] +matrix[35][159] * vector[35] +matrix[36][159] * vector[36] +matrix[37][159] * vector[37] +matrix[38][159] * vector[38] +matrix[39][159] * vector[39] +matrix[40][159] * vector[40] +matrix[41][159] * vector[41] +matrix[42][159] * vector[42] +matrix[43][159] * vector[43] +matrix[44][159] * vector[44] +matrix[45][159] * vector[45] +matrix[46][159] * vector[46] +matrix[47][159] * vector[47] +matrix[48][159] * vector[48] +matrix[49][159] * vector[49] +matrix[50][159] * vector[50] +matrix[51][159] * vector[51] +matrix[52][159] * vector[52] +matrix[53][159] * vector[53] +matrix[54][159] * vector[54] +matrix[55][159] * vector[55] +matrix[56][159] * vector[56] +matrix[57][159] * vector[57] +matrix[58][159] * vector[58] +matrix[59][159] * vector[59] +matrix[60][159] * vector[60] +matrix[61][159] * vector[61] +matrix[62][159] * vector[62] +matrix[63][159] * vector[63] +matrix[64][159] * vector[64] +matrix[65][159] * vector[65] +matrix[66][159] * vector[66] +matrix[67][159] * vector[67] +matrix[68][159] * vector[68] +matrix[69][159] * vector[69] +matrix[70][159] * vector[70] +matrix[71][159] * vector[71] +matrix[72][159] * vector[72] +matrix[73][159] * vector[73] +matrix[74][159] * vector[74] +matrix[75][159] * vector[75] +matrix[76][159] * vector[76] +matrix[77][159] * vector[77] +matrix[78][159] * vector[78] +matrix[79][159] * vector[79] +matrix[80][159] * vector[80] +matrix[81][159] * vector[81] +matrix[82][159] * vector[82] +matrix[83][159] * vector[83] +matrix[84][159] * vector[84] +matrix[85][159] * vector[85] +matrix[86][159] * vector[86] +matrix[87][159] * vector[87] +matrix[88][159] * vector[88] +matrix[89][159] * vector[89] +matrix[90][159] * vector[90] +matrix[91][159] * vector[91] +matrix[92][159] * vector[92] +matrix[93][159] * vector[93] +matrix[94][159] * vector[94] +matrix[95][159] * vector[95] +matrix[96][159] * vector[96] +matrix[97][159] * vector[97] +matrix[98][159] * vector[98] +matrix[99][159] * vector[99] +b[159];
assign result[160] = matrix[0][160] * vector[0] +matrix[1][160] * vector[1] +matrix[2][160] * vector[2] +matrix[3][160] * vector[3] +matrix[4][160] * vector[4] +matrix[5][160] * vector[5] +matrix[6][160] * vector[6] +matrix[7][160] * vector[7] +matrix[8][160] * vector[8] +matrix[9][160] * vector[9] +matrix[10][160] * vector[10] +matrix[11][160] * vector[11] +matrix[12][160] * vector[12] +matrix[13][160] * vector[13] +matrix[14][160] * vector[14] +matrix[15][160] * vector[15] +matrix[16][160] * vector[16] +matrix[17][160] * vector[17] +matrix[18][160] * vector[18] +matrix[19][160] * vector[19] +matrix[20][160] * vector[20] +matrix[21][160] * vector[21] +matrix[22][160] * vector[22] +matrix[23][160] * vector[23] +matrix[24][160] * vector[24] +matrix[25][160] * vector[25] +matrix[26][160] * vector[26] +matrix[27][160] * vector[27] +matrix[28][160] * vector[28] +matrix[29][160] * vector[29] +matrix[30][160] * vector[30] +matrix[31][160] * vector[31] +matrix[32][160] * vector[32] +matrix[33][160] * vector[33] +matrix[34][160] * vector[34] +matrix[35][160] * vector[35] +matrix[36][160] * vector[36] +matrix[37][160] * vector[37] +matrix[38][160] * vector[38] +matrix[39][160] * vector[39] +matrix[40][160] * vector[40] +matrix[41][160] * vector[41] +matrix[42][160] * vector[42] +matrix[43][160] * vector[43] +matrix[44][160] * vector[44] +matrix[45][160] * vector[45] +matrix[46][160] * vector[46] +matrix[47][160] * vector[47] +matrix[48][160] * vector[48] +matrix[49][160] * vector[49] +matrix[50][160] * vector[50] +matrix[51][160] * vector[51] +matrix[52][160] * vector[52] +matrix[53][160] * vector[53] +matrix[54][160] * vector[54] +matrix[55][160] * vector[55] +matrix[56][160] * vector[56] +matrix[57][160] * vector[57] +matrix[58][160] * vector[58] +matrix[59][160] * vector[59] +matrix[60][160] * vector[60] +matrix[61][160] * vector[61] +matrix[62][160] * vector[62] +matrix[63][160] * vector[63] +matrix[64][160] * vector[64] +matrix[65][160] * vector[65] +matrix[66][160] * vector[66] +matrix[67][160] * vector[67] +matrix[68][160] * vector[68] +matrix[69][160] * vector[69] +matrix[70][160] * vector[70] +matrix[71][160] * vector[71] +matrix[72][160] * vector[72] +matrix[73][160] * vector[73] +matrix[74][160] * vector[74] +matrix[75][160] * vector[75] +matrix[76][160] * vector[76] +matrix[77][160] * vector[77] +matrix[78][160] * vector[78] +matrix[79][160] * vector[79] +matrix[80][160] * vector[80] +matrix[81][160] * vector[81] +matrix[82][160] * vector[82] +matrix[83][160] * vector[83] +matrix[84][160] * vector[84] +matrix[85][160] * vector[85] +matrix[86][160] * vector[86] +matrix[87][160] * vector[87] +matrix[88][160] * vector[88] +matrix[89][160] * vector[89] +matrix[90][160] * vector[90] +matrix[91][160] * vector[91] +matrix[92][160] * vector[92] +matrix[93][160] * vector[93] +matrix[94][160] * vector[94] +matrix[95][160] * vector[95] +matrix[96][160] * vector[96] +matrix[97][160] * vector[97] +matrix[98][160] * vector[98] +matrix[99][160] * vector[99] +b[160];
assign result[161] = matrix[0][161] * vector[0] +matrix[1][161] * vector[1] +matrix[2][161] * vector[2] +matrix[3][161] * vector[3] +matrix[4][161] * vector[4] +matrix[5][161] * vector[5] +matrix[6][161] * vector[6] +matrix[7][161] * vector[7] +matrix[8][161] * vector[8] +matrix[9][161] * vector[9] +matrix[10][161] * vector[10] +matrix[11][161] * vector[11] +matrix[12][161] * vector[12] +matrix[13][161] * vector[13] +matrix[14][161] * vector[14] +matrix[15][161] * vector[15] +matrix[16][161] * vector[16] +matrix[17][161] * vector[17] +matrix[18][161] * vector[18] +matrix[19][161] * vector[19] +matrix[20][161] * vector[20] +matrix[21][161] * vector[21] +matrix[22][161] * vector[22] +matrix[23][161] * vector[23] +matrix[24][161] * vector[24] +matrix[25][161] * vector[25] +matrix[26][161] * vector[26] +matrix[27][161] * vector[27] +matrix[28][161] * vector[28] +matrix[29][161] * vector[29] +matrix[30][161] * vector[30] +matrix[31][161] * vector[31] +matrix[32][161] * vector[32] +matrix[33][161] * vector[33] +matrix[34][161] * vector[34] +matrix[35][161] * vector[35] +matrix[36][161] * vector[36] +matrix[37][161] * vector[37] +matrix[38][161] * vector[38] +matrix[39][161] * vector[39] +matrix[40][161] * vector[40] +matrix[41][161] * vector[41] +matrix[42][161] * vector[42] +matrix[43][161] * vector[43] +matrix[44][161] * vector[44] +matrix[45][161] * vector[45] +matrix[46][161] * vector[46] +matrix[47][161] * vector[47] +matrix[48][161] * vector[48] +matrix[49][161] * vector[49] +matrix[50][161] * vector[50] +matrix[51][161] * vector[51] +matrix[52][161] * vector[52] +matrix[53][161] * vector[53] +matrix[54][161] * vector[54] +matrix[55][161] * vector[55] +matrix[56][161] * vector[56] +matrix[57][161] * vector[57] +matrix[58][161] * vector[58] +matrix[59][161] * vector[59] +matrix[60][161] * vector[60] +matrix[61][161] * vector[61] +matrix[62][161] * vector[62] +matrix[63][161] * vector[63] +matrix[64][161] * vector[64] +matrix[65][161] * vector[65] +matrix[66][161] * vector[66] +matrix[67][161] * vector[67] +matrix[68][161] * vector[68] +matrix[69][161] * vector[69] +matrix[70][161] * vector[70] +matrix[71][161] * vector[71] +matrix[72][161] * vector[72] +matrix[73][161] * vector[73] +matrix[74][161] * vector[74] +matrix[75][161] * vector[75] +matrix[76][161] * vector[76] +matrix[77][161] * vector[77] +matrix[78][161] * vector[78] +matrix[79][161] * vector[79] +matrix[80][161] * vector[80] +matrix[81][161] * vector[81] +matrix[82][161] * vector[82] +matrix[83][161] * vector[83] +matrix[84][161] * vector[84] +matrix[85][161] * vector[85] +matrix[86][161] * vector[86] +matrix[87][161] * vector[87] +matrix[88][161] * vector[88] +matrix[89][161] * vector[89] +matrix[90][161] * vector[90] +matrix[91][161] * vector[91] +matrix[92][161] * vector[92] +matrix[93][161] * vector[93] +matrix[94][161] * vector[94] +matrix[95][161] * vector[95] +matrix[96][161] * vector[96] +matrix[97][161] * vector[97] +matrix[98][161] * vector[98] +matrix[99][161] * vector[99] +b[161];
assign result[162] = matrix[0][162] * vector[0] +matrix[1][162] * vector[1] +matrix[2][162] * vector[2] +matrix[3][162] * vector[3] +matrix[4][162] * vector[4] +matrix[5][162] * vector[5] +matrix[6][162] * vector[6] +matrix[7][162] * vector[7] +matrix[8][162] * vector[8] +matrix[9][162] * vector[9] +matrix[10][162] * vector[10] +matrix[11][162] * vector[11] +matrix[12][162] * vector[12] +matrix[13][162] * vector[13] +matrix[14][162] * vector[14] +matrix[15][162] * vector[15] +matrix[16][162] * vector[16] +matrix[17][162] * vector[17] +matrix[18][162] * vector[18] +matrix[19][162] * vector[19] +matrix[20][162] * vector[20] +matrix[21][162] * vector[21] +matrix[22][162] * vector[22] +matrix[23][162] * vector[23] +matrix[24][162] * vector[24] +matrix[25][162] * vector[25] +matrix[26][162] * vector[26] +matrix[27][162] * vector[27] +matrix[28][162] * vector[28] +matrix[29][162] * vector[29] +matrix[30][162] * vector[30] +matrix[31][162] * vector[31] +matrix[32][162] * vector[32] +matrix[33][162] * vector[33] +matrix[34][162] * vector[34] +matrix[35][162] * vector[35] +matrix[36][162] * vector[36] +matrix[37][162] * vector[37] +matrix[38][162] * vector[38] +matrix[39][162] * vector[39] +matrix[40][162] * vector[40] +matrix[41][162] * vector[41] +matrix[42][162] * vector[42] +matrix[43][162] * vector[43] +matrix[44][162] * vector[44] +matrix[45][162] * vector[45] +matrix[46][162] * vector[46] +matrix[47][162] * vector[47] +matrix[48][162] * vector[48] +matrix[49][162] * vector[49] +matrix[50][162] * vector[50] +matrix[51][162] * vector[51] +matrix[52][162] * vector[52] +matrix[53][162] * vector[53] +matrix[54][162] * vector[54] +matrix[55][162] * vector[55] +matrix[56][162] * vector[56] +matrix[57][162] * vector[57] +matrix[58][162] * vector[58] +matrix[59][162] * vector[59] +matrix[60][162] * vector[60] +matrix[61][162] * vector[61] +matrix[62][162] * vector[62] +matrix[63][162] * vector[63] +matrix[64][162] * vector[64] +matrix[65][162] * vector[65] +matrix[66][162] * vector[66] +matrix[67][162] * vector[67] +matrix[68][162] * vector[68] +matrix[69][162] * vector[69] +matrix[70][162] * vector[70] +matrix[71][162] * vector[71] +matrix[72][162] * vector[72] +matrix[73][162] * vector[73] +matrix[74][162] * vector[74] +matrix[75][162] * vector[75] +matrix[76][162] * vector[76] +matrix[77][162] * vector[77] +matrix[78][162] * vector[78] +matrix[79][162] * vector[79] +matrix[80][162] * vector[80] +matrix[81][162] * vector[81] +matrix[82][162] * vector[82] +matrix[83][162] * vector[83] +matrix[84][162] * vector[84] +matrix[85][162] * vector[85] +matrix[86][162] * vector[86] +matrix[87][162] * vector[87] +matrix[88][162] * vector[88] +matrix[89][162] * vector[89] +matrix[90][162] * vector[90] +matrix[91][162] * vector[91] +matrix[92][162] * vector[92] +matrix[93][162] * vector[93] +matrix[94][162] * vector[94] +matrix[95][162] * vector[95] +matrix[96][162] * vector[96] +matrix[97][162] * vector[97] +matrix[98][162] * vector[98] +matrix[99][162] * vector[99] +b[162];
assign result[163] = matrix[0][163] * vector[0] +matrix[1][163] * vector[1] +matrix[2][163] * vector[2] +matrix[3][163] * vector[3] +matrix[4][163] * vector[4] +matrix[5][163] * vector[5] +matrix[6][163] * vector[6] +matrix[7][163] * vector[7] +matrix[8][163] * vector[8] +matrix[9][163] * vector[9] +matrix[10][163] * vector[10] +matrix[11][163] * vector[11] +matrix[12][163] * vector[12] +matrix[13][163] * vector[13] +matrix[14][163] * vector[14] +matrix[15][163] * vector[15] +matrix[16][163] * vector[16] +matrix[17][163] * vector[17] +matrix[18][163] * vector[18] +matrix[19][163] * vector[19] +matrix[20][163] * vector[20] +matrix[21][163] * vector[21] +matrix[22][163] * vector[22] +matrix[23][163] * vector[23] +matrix[24][163] * vector[24] +matrix[25][163] * vector[25] +matrix[26][163] * vector[26] +matrix[27][163] * vector[27] +matrix[28][163] * vector[28] +matrix[29][163] * vector[29] +matrix[30][163] * vector[30] +matrix[31][163] * vector[31] +matrix[32][163] * vector[32] +matrix[33][163] * vector[33] +matrix[34][163] * vector[34] +matrix[35][163] * vector[35] +matrix[36][163] * vector[36] +matrix[37][163] * vector[37] +matrix[38][163] * vector[38] +matrix[39][163] * vector[39] +matrix[40][163] * vector[40] +matrix[41][163] * vector[41] +matrix[42][163] * vector[42] +matrix[43][163] * vector[43] +matrix[44][163] * vector[44] +matrix[45][163] * vector[45] +matrix[46][163] * vector[46] +matrix[47][163] * vector[47] +matrix[48][163] * vector[48] +matrix[49][163] * vector[49] +matrix[50][163] * vector[50] +matrix[51][163] * vector[51] +matrix[52][163] * vector[52] +matrix[53][163] * vector[53] +matrix[54][163] * vector[54] +matrix[55][163] * vector[55] +matrix[56][163] * vector[56] +matrix[57][163] * vector[57] +matrix[58][163] * vector[58] +matrix[59][163] * vector[59] +matrix[60][163] * vector[60] +matrix[61][163] * vector[61] +matrix[62][163] * vector[62] +matrix[63][163] * vector[63] +matrix[64][163] * vector[64] +matrix[65][163] * vector[65] +matrix[66][163] * vector[66] +matrix[67][163] * vector[67] +matrix[68][163] * vector[68] +matrix[69][163] * vector[69] +matrix[70][163] * vector[70] +matrix[71][163] * vector[71] +matrix[72][163] * vector[72] +matrix[73][163] * vector[73] +matrix[74][163] * vector[74] +matrix[75][163] * vector[75] +matrix[76][163] * vector[76] +matrix[77][163] * vector[77] +matrix[78][163] * vector[78] +matrix[79][163] * vector[79] +matrix[80][163] * vector[80] +matrix[81][163] * vector[81] +matrix[82][163] * vector[82] +matrix[83][163] * vector[83] +matrix[84][163] * vector[84] +matrix[85][163] * vector[85] +matrix[86][163] * vector[86] +matrix[87][163] * vector[87] +matrix[88][163] * vector[88] +matrix[89][163] * vector[89] +matrix[90][163] * vector[90] +matrix[91][163] * vector[91] +matrix[92][163] * vector[92] +matrix[93][163] * vector[93] +matrix[94][163] * vector[94] +matrix[95][163] * vector[95] +matrix[96][163] * vector[96] +matrix[97][163] * vector[97] +matrix[98][163] * vector[98] +matrix[99][163] * vector[99] +b[163];
assign result[164] = matrix[0][164] * vector[0] +matrix[1][164] * vector[1] +matrix[2][164] * vector[2] +matrix[3][164] * vector[3] +matrix[4][164] * vector[4] +matrix[5][164] * vector[5] +matrix[6][164] * vector[6] +matrix[7][164] * vector[7] +matrix[8][164] * vector[8] +matrix[9][164] * vector[9] +matrix[10][164] * vector[10] +matrix[11][164] * vector[11] +matrix[12][164] * vector[12] +matrix[13][164] * vector[13] +matrix[14][164] * vector[14] +matrix[15][164] * vector[15] +matrix[16][164] * vector[16] +matrix[17][164] * vector[17] +matrix[18][164] * vector[18] +matrix[19][164] * vector[19] +matrix[20][164] * vector[20] +matrix[21][164] * vector[21] +matrix[22][164] * vector[22] +matrix[23][164] * vector[23] +matrix[24][164] * vector[24] +matrix[25][164] * vector[25] +matrix[26][164] * vector[26] +matrix[27][164] * vector[27] +matrix[28][164] * vector[28] +matrix[29][164] * vector[29] +matrix[30][164] * vector[30] +matrix[31][164] * vector[31] +matrix[32][164] * vector[32] +matrix[33][164] * vector[33] +matrix[34][164] * vector[34] +matrix[35][164] * vector[35] +matrix[36][164] * vector[36] +matrix[37][164] * vector[37] +matrix[38][164] * vector[38] +matrix[39][164] * vector[39] +matrix[40][164] * vector[40] +matrix[41][164] * vector[41] +matrix[42][164] * vector[42] +matrix[43][164] * vector[43] +matrix[44][164] * vector[44] +matrix[45][164] * vector[45] +matrix[46][164] * vector[46] +matrix[47][164] * vector[47] +matrix[48][164] * vector[48] +matrix[49][164] * vector[49] +matrix[50][164] * vector[50] +matrix[51][164] * vector[51] +matrix[52][164] * vector[52] +matrix[53][164] * vector[53] +matrix[54][164] * vector[54] +matrix[55][164] * vector[55] +matrix[56][164] * vector[56] +matrix[57][164] * vector[57] +matrix[58][164] * vector[58] +matrix[59][164] * vector[59] +matrix[60][164] * vector[60] +matrix[61][164] * vector[61] +matrix[62][164] * vector[62] +matrix[63][164] * vector[63] +matrix[64][164] * vector[64] +matrix[65][164] * vector[65] +matrix[66][164] * vector[66] +matrix[67][164] * vector[67] +matrix[68][164] * vector[68] +matrix[69][164] * vector[69] +matrix[70][164] * vector[70] +matrix[71][164] * vector[71] +matrix[72][164] * vector[72] +matrix[73][164] * vector[73] +matrix[74][164] * vector[74] +matrix[75][164] * vector[75] +matrix[76][164] * vector[76] +matrix[77][164] * vector[77] +matrix[78][164] * vector[78] +matrix[79][164] * vector[79] +matrix[80][164] * vector[80] +matrix[81][164] * vector[81] +matrix[82][164] * vector[82] +matrix[83][164] * vector[83] +matrix[84][164] * vector[84] +matrix[85][164] * vector[85] +matrix[86][164] * vector[86] +matrix[87][164] * vector[87] +matrix[88][164] * vector[88] +matrix[89][164] * vector[89] +matrix[90][164] * vector[90] +matrix[91][164] * vector[91] +matrix[92][164] * vector[92] +matrix[93][164] * vector[93] +matrix[94][164] * vector[94] +matrix[95][164] * vector[95] +matrix[96][164] * vector[96] +matrix[97][164] * vector[97] +matrix[98][164] * vector[98] +matrix[99][164] * vector[99] +b[164];
assign result[165] = matrix[0][165] * vector[0] +matrix[1][165] * vector[1] +matrix[2][165] * vector[2] +matrix[3][165] * vector[3] +matrix[4][165] * vector[4] +matrix[5][165] * vector[5] +matrix[6][165] * vector[6] +matrix[7][165] * vector[7] +matrix[8][165] * vector[8] +matrix[9][165] * vector[9] +matrix[10][165] * vector[10] +matrix[11][165] * vector[11] +matrix[12][165] * vector[12] +matrix[13][165] * vector[13] +matrix[14][165] * vector[14] +matrix[15][165] * vector[15] +matrix[16][165] * vector[16] +matrix[17][165] * vector[17] +matrix[18][165] * vector[18] +matrix[19][165] * vector[19] +matrix[20][165] * vector[20] +matrix[21][165] * vector[21] +matrix[22][165] * vector[22] +matrix[23][165] * vector[23] +matrix[24][165] * vector[24] +matrix[25][165] * vector[25] +matrix[26][165] * vector[26] +matrix[27][165] * vector[27] +matrix[28][165] * vector[28] +matrix[29][165] * vector[29] +matrix[30][165] * vector[30] +matrix[31][165] * vector[31] +matrix[32][165] * vector[32] +matrix[33][165] * vector[33] +matrix[34][165] * vector[34] +matrix[35][165] * vector[35] +matrix[36][165] * vector[36] +matrix[37][165] * vector[37] +matrix[38][165] * vector[38] +matrix[39][165] * vector[39] +matrix[40][165] * vector[40] +matrix[41][165] * vector[41] +matrix[42][165] * vector[42] +matrix[43][165] * vector[43] +matrix[44][165] * vector[44] +matrix[45][165] * vector[45] +matrix[46][165] * vector[46] +matrix[47][165] * vector[47] +matrix[48][165] * vector[48] +matrix[49][165] * vector[49] +matrix[50][165] * vector[50] +matrix[51][165] * vector[51] +matrix[52][165] * vector[52] +matrix[53][165] * vector[53] +matrix[54][165] * vector[54] +matrix[55][165] * vector[55] +matrix[56][165] * vector[56] +matrix[57][165] * vector[57] +matrix[58][165] * vector[58] +matrix[59][165] * vector[59] +matrix[60][165] * vector[60] +matrix[61][165] * vector[61] +matrix[62][165] * vector[62] +matrix[63][165] * vector[63] +matrix[64][165] * vector[64] +matrix[65][165] * vector[65] +matrix[66][165] * vector[66] +matrix[67][165] * vector[67] +matrix[68][165] * vector[68] +matrix[69][165] * vector[69] +matrix[70][165] * vector[70] +matrix[71][165] * vector[71] +matrix[72][165] * vector[72] +matrix[73][165] * vector[73] +matrix[74][165] * vector[74] +matrix[75][165] * vector[75] +matrix[76][165] * vector[76] +matrix[77][165] * vector[77] +matrix[78][165] * vector[78] +matrix[79][165] * vector[79] +matrix[80][165] * vector[80] +matrix[81][165] * vector[81] +matrix[82][165] * vector[82] +matrix[83][165] * vector[83] +matrix[84][165] * vector[84] +matrix[85][165] * vector[85] +matrix[86][165] * vector[86] +matrix[87][165] * vector[87] +matrix[88][165] * vector[88] +matrix[89][165] * vector[89] +matrix[90][165] * vector[90] +matrix[91][165] * vector[91] +matrix[92][165] * vector[92] +matrix[93][165] * vector[93] +matrix[94][165] * vector[94] +matrix[95][165] * vector[95] +matrix[96][165] * vector[96] +matrix[97][165] * vector[97] +matrix[98][165] * vector[98] +matrix[99][165] * vector[99] +b[165];
assign result[166] = matrix[0][166] * vector[0] +matrix[1][166] * vector[1] +matrix[2][166] * vector[2] +matrix[3][166] * vector[3] +matrix[4][166] * vector[4] +matrix[5][166] * vector[5] +matrix[6][166] * vector[6] +matrix[7][166] * vector[7] +matrix[8][166] * vector[8] +matrix[9][166] * vector[9] +matrix[10][166] * vector[10] +matrix[11][166] * vector[11] +matrix[12][166] * vector[12] +matrix[13][166] * vector[13] +matrix[14][166] * vector[14] +matrix[15][166] * vector[15] +matrix[16][166] * vector[16] +matrix[17][166] * vector[17] +matrix[18][166] * vector[18] +matrix[19][166] * vector[19] +matrix[20][166] * vector[20] +matrix[21][166] * vector[21] +matrix[22][166] * vector[22] +matrix[23][166] * vector[23] +matrix[24][166] * vector[24] +matrix[25][166] * vector[25] +matrix[26][166] * vector[26] +matrix[27][166] * vector[27] +matrix[28][166] * vector[28] +matrix[29][166] * vector[29] +matrix[30][166] * vector[30] +matrix[31][166] * vector[31] +matrix[32][166] * vector[32] +matrix[33][166] * vector[33] +matrix[34][166] * vector[34] +matrix[35][166] * vector[35] +matrix[36][166] * vector[36] +matrix[37][166] * vector[37] +matrix[38][166] * vector[38] +matrix[39][166] * vector[39] +matrix[40][166] * vector[40] +matrix[41][166] * vector[41] +matrix[42][166] * vector[42] +matrix[43][166] * vector[43] +matrix[44][166] * vector[44] +matrix[45][166] * vector[45] +matrix[46][166] * vector[46] +matrix[47][166] * vector[47] +matrix[48][166] * vector[48] +matrix[49][166] * vector[49] +matrix[50][166] * vector[50] +matrix[51][166] * vector[51] +matrix[52][166] * vector[52] +matrix[53][166] * vector[53] +matrix[54][166] * vector[54] +matrix[55][166] * vector[55] +matrix[56][166] * vector[56] +matrix[57][166] * vector[57] +matrix[58][166] * vector[58] +matrix[59][166] * vector[59] +matrix[60][166] * vector[60] +matrix[61][166] * vector[61] +matrix[62][166] * vector[62] +matrix[63][166] * vector[63] +matrix[64][166] * vector[64] +matrix[65][166] * vector[65] +matrix[66][166] * vector[66] +matrix[67][166] * vector[67] +matrix[68][166] * vector[68] +matrix[69][166] * vector[69] +matrix[70][166] * vector[70] +matrix[71][166] * vector[71] +matrix[72][166] * vector[72] +matrix[73][166] * vector[73] +matrix[74][166] * vector[74] +matrix[75][166] * vector[75] +matrix[76][166] * vector[76] +matrix[77][166] * vector[77] +matrix[78][166] * vector[78] +matrix[79][166] * vector[79] +matrix[80][166] * vector[80] +matrix[81][166] * vector[81] +matrix[82][166] * vector[82] +matrix[83][166] * vector[83] +matrix[84][166] * vector[84] +matrix[85][166] * vector[85] +matrix[86][166] * vector[86] +matrix[87][166] * vector[87] +matrix[88][166] * vector[88] +matrix[89][166] * vector[89] +matrix[90][166] * vector[90] +matrix[91][166] * vector[91] +matrix[92][166] * vector[92] +matrix[93][166] * vector[93] +matrix[94][166] * vector[94] +matrix[95][166] * vector[95] +matrix[96][166] * vector[96] +matrix[97][166] * vector[97] +matrix[98][166] * vector[98] +matrix[99][166] * vector[99] +b[166];
assign result[167] = matrix[0][167] * vector[0] +matrix[1][167] * vector[1] +matrix[2][167] * vector[2] +matrix[3][167] * vector[3] +matrix[4][167] * vector[4] +matrix[5][167] * vector[5] +matrix[6][167] * vector[6] +matrix[7][167] * vector[7] +matrix[8][167] * vector[8] +matrix[9][167] * vector[9] +matrix[10][167] * vector[10] +matrix[11][167] * vector[11] +matrix[12][167] * vector[12] +matrix[13][167] * vector[13] +matrix[14][167] * vector[14] +matrix[15][167] * vector[15] +matrix[16][167] * vector[16] +matrix[17][167] * vector[17] +matrix[18][167] * vector[18] +matrix[19][167] * vector[19] +matrix[20][167] * vector[20] +matrix[21][167] * vector[21] +matrix[22][167] * vector[22] +matrix[23][167] * vector[23] +matrix[24][167] * vector[24] +matrix[25][167] * vector[25] +matrix[26][167] * vector[26] +matrix[27][167] * vector[27] +matrix[28][167] * vector[28] +matrix[29][167] * vector[29] +matrix[30][167] * vector[30] +matrix[31][167] * vector[31] +matrix[32][167] * vector[32] +matrix[33][167] * vector[33] +matrix[34][167] * vector[34] +matrix[35][167] * vector[35] +matrix[36][167] * vector[36] +matrix[37][167] * vector[37] +matrix[38][167] * vector[38] +matrix[39][167] * vector[39] +matrix[40][167] * vector[40] +matrix[41][167] * vector[41] +matrix[42][167] * vector[42] +matrix[43][167] * vector[43] +matrix[44][167] * vector[44] +matrix[45][167] * vector[45] +matrix[46][167] * vector[46] +matrix[47][167] * vector[47] +matrix[48][167] * vector[48] +matrix[49][167] * vector[49] +matrix[50][167] * vector[50] +matrix[51][167] * vector[51] +matrix[52][167] * vector[52] +matrix[53][167] * vector[53] +matrix[54][167] * vector[54] +matrix[55][167] * vector[55] +matrix[56][167] * vector[56] +matrix[57][167] * vector[57] +matrix[58][167] * vector[58] +matrix[59][167] * vector[59] +matrix[60][167] * vector[60] +matrix[61][167] * vector[61] +matrix[62][167] * vector[62] +matrix[63][167] * vector[63] +matrix[64][167] * vector[64] +matrix[65][167] * vector[65] +matrix[66][167] * vector[66] +matrix[67][167] * vector[67] +matrix[68][167] * vector[68] +matrix[69][167] * vector[69] +matrix[70][167] * vector[70] +matrix[71][167] * vector[71] +matrix[72][167] * vector[72] +matrix[73][167] * vector[73] +matrix[74][167] * vector[74] +matrix[75][167] * vector[75] +matrix[76][167] * vector[76] +matrix[77][167] * vector[77] +matrix[78][167] * vector[78] +matrix[79][167] * vector[79] +matrix[80][167] * vector[80] +matrix[81][167] * vector[81] +matrix[82][167] * vector[82] +matrix[83][167] * vector[83] +matrix[84][167] * vector[84] +matrix[85][167] * vector[85] +matrix[86][167] * vector[86] +matrix[87][167] * vector[87] +matrix[88][167] * vector[88] +matrix[89][167] * vector[89] +matrix[90][167] * vector[90] +matrix[91][167] * vector[91] +matrix[92][167] * vector[92] +matrix[93][167] * vector[93] +matrix[94][167] * vector[94] +matrix[95][167] * vector[95] +matrix[96][167] * vector[96] +matrix[97][167] * vector[97] +matrix[98][167] * vector[98] +matrix[99][167] * vector[99] +b[167];
assign result[168] = matrix[0][168] * vector[0] +matrix[1][168] * vector[1] +matrix[2][168] * vector[2] +matrix[3][168] * vector[3] +matrix[4][168] * vector[4] +matrix[5][168] * vector[5] +matrix[6][168] * vector[6] +matrix[7][168] * vector[7] +matrix[8][168] * vector[8] +matrix[9][168] * vector[9] +matrix[10][168] * vector[10] +matrix[11][168] * vector[11] +matrix[12][168] * vector[12] +matrix[13][168] * vector[13] +matrix[14][168] * vector[14] +matrix[15][168] * vector[15] +matrix[16][168] * vector[16] +matrix[17][168] * vector[17] +matrix[18][168] * vector[18] +matrix[19][168] * vector[19] +matrix[20][168] * vector[20] +matrix[21][168] * vector[21] +matrix[22][168] * vector[22] +matrix[23][168] * vector[23] +matrix[24][168] * vector[24] +matrix[25][168] * vector[25] +matrix[26][168] * vector[26] +matrix[27][168] * vector[27] +matrix[28][168] * vector[28] +matrix[29][168] * vector[29] +matrix[30][168] * vector[30] +matrix[31][168] * vector[31] +matrix[32][168] * vector[32] +matrix[33][168] * vector[33] +matrix[34][168] * vector[34] +matrix[35][168] * vector[35] +matrix[36][168] * vector[36] +matrix[37][168] * vector[37] +matrix[38][168] * vector[38] +matrix[39][168] * vector[39] +matrix[40][168] * vector[40] +matrix[41][168] * vector[41] +matrix[42][168] * vector[42] +matrix[43][168] * vector[43] +matrix[44][168] * vector[44] +matrix[45][168] * vector[45] +matrix[46][168] * vector[46] +matrix[47][168] * vector[47] +matrix[48][168] * vector[48] +matrix[49][168] * vector[49] +matrix[50][168] * vector[50] +matrix[51][168] * vector[51] +matrix[52][168] * vector[52] +matrix[53][168] * vector[53] +matrix[54][168] * vector[54] +matrix[55][168] * vector[55] +matrix[56][168] * vector[56] +matrix[57][168] * vector[57] +matrix[58][168] * vector[58] +matrix[59][168] * vector[59] +matrix[60][168] * vector[60] +matrix[61][168] * vector[61] +matrix[62][168] * vector[62] +matrix[63][168] * vector[63] +matrix[64][168] * vector[64] +matrix[65][168] * vector[65] +matrix[66][168] * vector[66] +matrix[67][168] * vector[67] +matrix[68][168] * vector[68] +matrix[69][168] * vector[69] +matrix[70][168] * vector[70] +matrix[71][168] * vector[71] +matrix[72][168] * vector[72] +matrix[73][168] * vector[73] +matrix[74][168] * vector[74] +matrix[75][168] * vector[75] +matrix[76][168] * vector[76] +matrix[77][168] * vector[77] +matrix[78][168] * vector[78] +matrix[79][168] * vector[79] +matrix[80][168] * vector[80] +matrix[81][168] * vector[81] +matrix[82][168] * vector[82] +matrix[83][168] * vector[83] +matrix[84][168] * vector[84] +matrix[85][168] * vector[85] +matrix[86][168] * vector[86] +matrix[87][168] * vector[87] +matrix[88][168] * vector[88] +matrix[89][168] * vector[89] +matrix[90][168] * vector[90] +matrix[91][168] * vector[91] +matrix[92][168] * vector[92] +matrix[93][168] * vector[93] +matrix[94][168] * vector[94] +matrix[95][168] * vector[95] +matrix[96][168] * vector[96] +matrix[97][168] * vector[97] +matrix[98][168] * vector[98] +matrix[99][168] * vector[99] +b[168];
assign result[169] = matrix[0][169] * vector[0] +matrix[1][169] * vector[1] +matrix[2][169] * vector[2] +matrix[3][169] * vector[3] +matrix[4][169] * vector[4] +matrix[5][169] * vector[5] +matrix[6][169] * vector[6] +matrix[7][169] * vector[7] +matrix[8][169] * vector[8] +matrix[9][169] * vector[9] +matrix[10][169] * vector[10] +matrix[11][169] * vector[11] +matrix[12][169] * vector[12] +matrix[13][169] * vector[13] +matrix[14][169] * vector[14] +matrix[15][169] * vector[15] +matrix[16][169] * vector[16] +matrix[17][169] * vector[17] +matrix[18][169] * vector[18] +matrix[19][169] * vector[19] +matrix[20][169] * vector[20] +matrix[21][169] * vector[21] +matrix[22][169] * vector[22] +matrix[23][169] * vector[23] +matrix[24][169] * vector[24] +matrix[25][169] * vector[25] +matrix[26][169] * vector[26] +matrix[27][169] * vector[27] +matrix[28][169] * vector[28] +matrix[29][169] * vector[29] +matrix[30][169] * vector[30] +matrix[31][169] * vector[31] +matrix[32][169] * vector[32] +matrix[33][169] * vector[33] +matrix[34][169] * vector[34] +matrix[35][169] * vector[35] +matrix[36][169] * vector[36] +matrix[37][169] * vector[37] +matrix[38][169] * vector[38] +matrix[39][169] * vector[39] +matrix[40][169] * vector[40] +matrix[41][169] * vector[41] +matrix[42][169] * vector[42] +matrix[43][169] * vector[43] +matrix[44][169] * vector[44] +matrix[45][169] * vector[45] +matrix[46][169] * vector[46] +matrix[47][169] * vector[47] +matrix[48][169] * vector[48] +matrix[49][169] * vector[49] +matrix[50][169] * vector[50] +matrix[51][169] * vector[51] +matrix[52][169] * vector[52] +matrix[53][169] * vector[53] +matrix[54][169] * vector[54] +matrix[55][169] * vector[55] +matrix[56][169] * vector[56] +matrix[57][169] * vector[57] +matrix[58][169] * vector[58] +matrix[59][169] * vector[59] +matrix[60][169] * vector[60] +matrix[61][169] * vector[61] +matrix[62][169] * vector[62] +matrix[63][169] * vector[63] +matrix[64][169] * vector[64] +matrix[65][169] * vector[65] +matrix[66][169] * vector[66] +matrix[67][169] * vector[67] +matrix[68][169] * vector[68] +matrix[69][169] * vector[69] +matrix[70][169] * vector[70] +matrix[71][169] * vector[71] +matrix[72][169] * vector[72] +matrix[73][169] * vector[73] +matrix[74][169] * vector[74] +matrix[75][169] * vector[75] +matrix[76][169] * vector[76] +matrix[77][169] * vector[77] +matrix[78][169] * vector[78] +matrix[79][169] * vector[79] +matrix[80][169] * vector[80] +matrix[81][169] * vector[81] +matrix[82][169] * vector[82] +matrix[83][169] * vector[83] +matrix[84][169] * vector[84] +matrix[85][169] * vector[85] +matrix[86][169] * vector[86] +matrix[87][169] * vector[87] +matrix[88][169] * vector[88] +matrix[89][169] * vector[89] +matrix[90][169] * vector[90] +matrix[91][169] * vector[91] +matrix[92][169] * vector[92] +matrix[93][169] * vector[93] +matrix[94][169] * vector[94] +matrix[95][169] * vector[95] +matrix[96][169] * vector[96] +matrix[97][169] * vector[97] +matrix[98][169] * vector[98] +matrix[99][169] * vector[99] +b[169];
assign result[170] = matrix[0][170] * vector[0] +matrix[1][170] * vector[1] +matrix[2][170] * vector[2] +matrix[3][170] * vector[3] +matrix[4][170] * vector[4] +matrix[5][170] * vector[5] +matrix[6][170] * vector[6] +matrix[7][170] * vector[7] +matrix[8][170] * vector[8] +matrix[9][170] * vector[9] +matrix[10][170] * vector[10] +matrix[11][170] * vector[11] +matrix[12][170] * vector[12] +matrix[13][170] * vector[13] +matrix[14][170] * vector[14] +matrix[15][170] * vector[15] +matrix[16][170] * vector[16] +matrix[17][170] * vector[17] +matrix[18][170] * vector[18] +matrix[19][170] * vector[19] +matrix[20][170] * vector[20] +matrix[21][170] * vector[21] +matrix[22][170] * vector[22] +matrix[23][170] * vector[23] +matrix[24][170] * vector[24] +matrix[25][170] * vector[25] +matrix[26][170] * vector[26] +matrix[27][170] * vector[27] +matrix[28][170] * vector[28] +matrix[29][170] * vector[29] +matrix[30][170] * vector[30] +matrix[31][170] * vector[31] +matrix[32][170] * vector[32] +matrix[33][170] * vector[33] +matrix[34][170] * vector[34] +matrix[35][170] * vector[35] +matrix[36][170] * vector[36] +matrix[37][170] * vector[37] +matrix[38][170] * vector[38] +matrix[39][170] * vector[39] +matrix[40][170] * vector[40] +matrix[41][170] * vector[41] +matrix[42][170] * vector[42] +matrix[43][170] * vector[43] +matrix[44][170] * vector[44] +matrix[45][170] * vector[45] +matrix[46][170] * vector[46] +matrix[47][170] * vector[47] +matrix[48][170] * vector[48] +matrix[49][170] * vector[49] +matrix[50][170] * vector[50] +matrix[51][170] * vector[51] +matrix[52][170] * vector[52] +matrix[53][170] * vector[53] +matrix[54][170] * vector[54] +matrix[55][170] * vector[55] +matrix[56][170] * vector[56] +matrix[57][170] * vector[57] +matrix[58][170] * vector[58] +matrix[59][170] * vector[59] +matrix[60][170] * vector[60] +matrix[61][170] * vector[61] +matrix[62][170] * vector[62] +matrix[63][170] * vector[63] +matrix[64][170] * vector[64] +matrix[65][170] * vector[65] +matrix[66][170] * vector[66] +matrix[67][170] * vector[67] +matrix[68][170] * vector[68] +matrix[69][170] * vector[69] +matrix[70][170] * vector[70] +matrix[71][170] * vector[71] +matrix[72][170] * vector[72] +matrix[73][170] * vector[73] +matrix[74][170] * vector[74] +matrix[75][170] * vector[75] +matrix[76][170] * vector[76] +matrix[77][170] * vector[77] +matrix[78][170] * vector[78] +matrix[79][170] * vector[79] +matrix[80][170] * vector[80] +matrix[81][170] * vector[81] +matrix[82][170] * vector[82] +matrix[83][170] * vector[83] +matrix[84][170] * vector[84] +matrix[85][170] * vector[85] +matrix[86][170] * vector[86] +matrix[87][170] * vector[87] +matrix[88][170] * vector[88] +matrix[89][170] * vector[89] +matrix[90][170] * vector[90] +matrix[91][170] * vector[91] +matrix[92][170] * vector[92] +matrix[93][170] * vector[93] +matrix[94][170] * vector[94] +matrix[95][170] * vector[95] +matrix[96][170] * vector[96] +matrix[97][170] * vector[97] +matrix[98][170] * vector[98] +matrix[99][170] * vector[99] +b[170];
assign result[171] = matrix[0][171] * vector[0] +matrix[1][171] * vector[1] +matrix[2][171] * vector[2] +matrix[3][171] * vector[3] +matrix[4][171] * vector[4] +matrix[5][171] * vector[5] +matrix[6][171] * vector[6] +matrix[7][171] * vector[7] +matrix[8][171] * vector[8] +matrix[9][171] * vector[9] +matrix[10][171] * vector[10] +matrix[11][171] * vector[11] +matrix[12][171] * vector[12] +matrix[13][171] * vector[13] +matrix[14][171] * vector[14] +matrix[15][171] * vector[15] +matrix[16][171] * vector[16] +matrix[17][171] * vector[17] +matrix[18][171] * vector[18] +matrix[19][171] * vector[19] +matrix[20][171] * vector[20] +matrix[21][171] * vector[21] +matrix[22][171] * vector[22] +matrix[23][171] * vector[23] +matrix[24][171] * vector[24] +matrix[25][171] * vector[25] +matrix[26][171] * vector[26] +matrix[27][171] * vector[27] +matrix[28][171] * vector[28] +matrix[29][171] * vector[29] +matrix[30][171] * vector[30] +matrix[31][171] * vector[31] +matrix[32][171] * vector[32] +matrix[33][171] * vector[33] +matrix[34][171] * vector[34] +matrix[35][171] * vector[35] +matrix[36][171] * vector[36] +matrix[37][171] * vector[37] +matrix[38][171] * vector[38] +matrix[39][171] * vector[39] +matrix[40][171] * vector[40] +matrix[41][171] * vector[41] +matrix[42][171] * vector[42] +matrix[43][171] * vector[43] +matrix[44][171] * vector[44] +matrix[45][171] * vector[45] +matrix[46][171] * vector[46] +matrix[47][171] * vector[47] +matrix[48][171] * vector[48] +matrix[49][171] * vector[49] +matrix[50][171] * vector[50] +matrix[51][171] * vector[51] +matrix[52][171] * vector[52] +matrix[53][171] * vector[53] +matrix[54][171] * vector[54] +matrix[55][171] * vector[55] +matrix[56][171] * vector[56] +matrix[57][171] * vector[57] +matrix[58][171] * vector[58] +matrix[59][171] * vector[59] +matrix[60][171] * vector[60] +matrix[61][171] * vector[61] +matrix[62][171] * vector[62] +matrix[63][171] * vector[63] +matrix[64][171] * vector[64] +matrix[65][171] * vector[65] +matrix[66][171] * vector[66] +matrix[67][171] * vector[67] +matrix[68][171] * vector[68] +matrix[69][171] * vector[69] +matrix[70][171] * vector[70] +matrix[71][171] * vector[71] +matrix[72][171] * vector[72] +matrix[73][171] * vector[73] +matrix[74][171] * vector[74] +matrix[75][171] * vector[75] +matrix[76][171] * vector[76] +matrix[77][171] * vector[77] +matrix[78][171] * vector[78] +matrix[79][171] * vector[79] +matrix[80][171] * vector[80] +matrix[81][171] * vector[81] +matrix[82][171] * vector[82] +matrix[83][171] * vector[83] +matrix[84][171] * vector[84] +matrix[85][171] * vector[85] +matrix[86][171] * vector[86] +matrix[87][171] * vector[87] +matrix[88][171] * vector[88] +matrix[89][171] * vector[89] +matrix[90][171] * vector[90] +matrix[91][171] * vector[91] +matrix[92][171] * vector[92] +matrix[93][171] * vector[93] +matrix[94][171] * vector[94] +matrix[95][171] * vector[95] +matrix[96][171] * vector[96] +matrix[97][171] * vector[97] +matrix[98][171] * vector[98] +matrix[99][171] * vector[99] +b[171];
assign result[172] = matrix[0][172] * vector[0] +matrix[1][172] * vector[1] +matrix[2][172] * vector[2] +matrix[3][172] * vector[3] +matrix[4][172] * vector[4] +matrix[5][172] * vector[5] +matrix[6][172] * vector[6] +matrix[7][172] * vector[7] +matrix[8][172] * vector[8] +matrix[9][172] * vector[9] +matrix[10][172] * vector[10] +matrix[11][172] * vector[11] +matrix[12][172] * vector[12] +matrix[13][172] * vector[13] +matrix[14][172] * vector[14] +matrix[15][172] * vector[15] +matrix[16][172] * vector[16] +matrix[17][172] * vector[17] +matrix[18][172] * vector[18] +matrix[19][172] * vector[19] +matrix[20][172] * vector[20] +matrix[21][172] * vector[21] +matrix[22][172] * vector[22] +matrix[23][172] * vector[23] +matrix[24][172] * vector[24] +matrix[25][172] * vector[25] +matrix[26][172] * vector[26] +matrix[27][172] * vector[27] +matrix[28][172] * vector[28] +matrix[29][172] * vector[29] +matrix[30][172] * vector[30] +matrix[31][172] * vector[31] +matrix[32][172] * vector[32] +matrix[33][172] * vector[33] +matrix[34][172] * vector[34] +matrix[35][172] * vector[35] +matrix[36][172] * vector[36] +matrix[37][172] * vector[37] +matrix[38][172] * vector[38] +matrix[39][172] * vector[39] +matrix[40][172] * vector[40] +matrix[41][172] * vector[41] +matrix[42][172] * vector[42] +matrix[43][172] * vector[43] +matrix[44][172] * vector[44] +matrix[45][172] * vector[45] +matrix[46][172] * vector[46] +matrix[47][172] * vector[47] +matrix[48][172] * vector[48] +matrix[49][172] * vector[49] +matrix[50][172] * vector[50] +matrix[51][172] * vector[51] +matrix[52][172] * vector[52] +matrix[53][172] * vector[53] +matrix[54][172] * vector[54] +matrix[55][172] * vector[55] +matrix[56][172] * vector[56] +matrix[57][172] * vector[57] +matrix[58][172] * vector[58] +matrix[59][172] * vector[59] +matrix[60][172] * vector[60] +matrix[61][172] * vector[61] +matrix[62][172] * vector[62] +matrix[63][172] * vector[63] +matrix[64][172] * vector[64] +matrix[65][172] * vector[65] +matrix[66][172] * vector[66] +matrix[67][172] * vector[67] +matrix[68][172] * vector[68] +matrix[69][172] * vector[69] +matrix[70][172] * vector[70] +matrix[71][172] * vector[71] +matrix[72][172] * vector[72] +matrix[73][172] * vector[73] +matrix[74][172] * vector[74] +matrix[75][172] * vector[75] +matrix[76][172] * vector[76] +matrix[77][172] * vector[77] +matrix[78][172] * vector[78] +matrix[79][172] * vector[79] +matrix[80][172] * vector[80] +matrix[81][172] * vector[81] +matrix[82][172] * vector[82] +matrix[83][172] * vector[83] +matrix[84][172] * vector[84] +matrix[85][172] * vector[85] +matrix[86][172] * vector[86] +matrix[87][172] * vector[87] +matrix[88][172] * vector[88] +matrix[89][172] * vector[89] +matrix[90][172] * vector[90] +matrix[91][172] * vector[91] +matrix[92][172] * vector[92] +matrix[93][172] * vector[93] +matrix[94][172] * vector[94] +matrix[95][172] * vector[95] +matrix[96][172] * vector[96] +matrix[97][172] * vector[97] +matrix[98][172] * vector[98] +matrix[99][172] * vector[99] +b[172];
assign result[173] = matrix[0][173] * vector[0] +matrix[1][173] * vector[1] +matrix[2][173] * vector[2] +matrix[3][173] * vector[3] +matrix[4][173] * vector[4] +matrix[5][173] * vector[5] +matrix[6][173] * vector[6] +matrix[7][173] * vector[7] +matrix[8][173] * vector[8] +matrix[9][173] * vector[9] +matrix[10][173] * vector[10] +matrix[11][173] * vector[11] +matrix[12][173] * vector[12] +matrix[13][173] * vector[13] +matrix[14][173] * vector[14] +matrix[15][173] * vector[15] +matrix[16][173] * vector[16] +matrix[17][173] * vector[17] +matrix[18][173] * vector[18] +matrix[19][173] * vector[19] +matrix[20][173] * vector[20] +matrix[21][173] * vector[21] +matrix[22][173] * vector[22] +matrix[23][173] * vector[23] +matrix[24][173] * vector[24] +matrix[25][173] * vector[25] +matrix[26][173] * vector[26] +matrix[27][173] * vector[27] +matrix[28][173] * vector[28] +matrix[29][173] * vector[29] +matrix[30][173] * vector[30] +matrix[31][173] * vector[31] +matrix[32][173] * vector[32] +matrix[33][173] * vector[33] +matrix[34][173] * vector[34] +matrix[35][173] * vector[35] +matrix[36][173] * vector[36] +matrix[37][173] * vector[37] +matrix[38][173] * vector[38] +matrix[39][173] * vector[39] +matrix[40][173] * vector[40] +matrix[41][173] * vector[41] +matrix[42][173] * vector[42] +matrix[43][173] * vector[43] +matrix[44][173] * vector[44] +matrix[45][173] * vector[45] +matrix[46][173] * vector[46] +matrix[47][173] * vector[47] +matrix[48][173] * vector[48] +matrix[49][173] * vector[49] +matrix[50][173] * vector[50] +matrix[51][173] * vector[51] +matrix[52][173] * vector[52] +matrix[53][173] * vector[53] +matrix[54][173] * vector[54] +matrix[55][173] * vector[55] +matrix[56][173] * vector[56] +matrix[57][173] * vector[57] +matrix[58][173] * vector[58] +matrix[59][173] * vector[59] +matrix[60][173] * vector[60] +matrix[61][173] * vector[61] +matrix[62][173] * vector[62] +matrix[63][173] * vector[63] +matrix[64][173] * vector[64] +matrix[65][173] * vector[65] +matrix[66][173] * vector[66] +matrix[67][173] * vector[67] +matrix[68][173] * vector[68] +matrix[69][173] * vector[69] +matrix[70][173] * vector[70] +matrix[71][173] * vector[71] +matrix[72][173] * vector[72] +matrix[73][173] * vector[73] +matrix[74][173] * vector[74] +matrix[75][173] * vector[75] +matrix[76][173] * vector[76] +matrix[77][173] * vector[77] +matrix[78][173] * vector[78] +matrix[79][173] * vector[79] +matrix[80][173] * vector[80] +matrix[81][173] * vector[81] +matrix[82][173] * vector[82] +matrix[83][173] * vector[83] +matrix[84][173] * vector[84] +matrix[85][173] * vector[85] +matrix[86][173] * vector[86] +matrix[87][173] * vector[87] +matrix[88][173] * vector[88] +matrix[89][173] * vector[89] +matrix[90][173] * vector[90] +matrix[91][173] * vector[91] +matrix[92][173] * vector[92] +matrix[93][173] * vector[93] +matrix[94][173] * vector[94] +matrix[95][173] * vector[95] +matrix[96][173] * vector[96] +matrix[97][173] * vector[97] +matrix[98][173] * vector[98] +matrix[99][173] * vector[99] +b[173];
assign result[174] = matrix[0][174] * vector[0] +matrix[1][174] * vector[1] +matrix[2][174] * vector[2] +matrix[3][174] * vector[3] +matrix[4][174] * vector[4] +matrix[5][174] * vector[5] +matrix[6][174] * vector[6] +matrix[7][174] * vector[7] +matrix[8][174] * vector[8] +matrix[9][174] * vector[9] +matrix[10][174] * vector[10] +matrix[11][174] * vector[11] +matrix[12][174] * vector[12] +matrix[13][174] * vector[13] +matrix[14][174] * vector[14] +matrix[15][174] * vector[15] +matrix[16][174] * vector[16] +matrix[17][174] * vector[17] +matrix[18][174] * vector[18] +matrix[19][174] * vector[19] +matrix[20][174] * vector[20] +matrix[21][174] * vector[21] +matrix[22][174] * vector[22] +matrix[23][174] * vector[23] +matrix[24][174] * vector[24] +matrix[25][174] * vector[25] +matrix[26][174] * vector[26] +matrix[27][174] * vector[27] +matrix[28][174] * vector[28] +matrix[29][174] * vector[29] +matrix[30][174] * vector[30] +matrix[31][174] * vector[31] +matrix[32][174] * vector[32] +matrix[33][174] * vector[33] +matrix[34][174] * vector[34] +matrix[35][174] * vector[35] +matrix[36][174] * vector[36] +matrix[37][174] * vector[37] +matrix[38][174] * vector[38] +matrix[39][174] * vector[39] +matrix[40][174] * vector[40] +matrix[41][174] * vector[41] +matrix[42][174] * vector[42] +matrix[43][174] * vector[43] +matrix[44][174] * vector[44] +matrix[45][174] * vector[45] +matrix[46][174] * vector[46] +matrix[47][174] * vector[47] +matrix[48][174] * vector[48] +matrix[49][174] * vector[49] +matrix[50][174] * vector[50] +matrix[51][174] * vector[51] +matrix[52][174] * vector[52] +matrix[53][174] * vector[53] +matrix[54][174] * vector[54] +matrix[55][174] * vector[55] +matrix[56][174] * vector[56] +matrix[57][174] * vector[57] +matrix[58][174] * vector[58] +matrix[59][174] * vector[59] +matrix[60][174] * vector[60] +matrix[61][174] * vector[61] +matrix[62][174] * vector[62] +matrix[63][174] * vector[63] +matrix[64][174] * vector[64] +matrix[65][174] * vector[65] +matrix[66][174] * vector[66] +matrix[67][174] * vector[67] +matrix[68][174] * vector[68] +matrix[69][174] * vector[69] +matrix[70][174] * vector[70] +matrix[71][174] * vector[71] +matrix[72][174] * vector[72] +matrix[73][174] * vector[73] +matrix[74][174] * vector[74] +matrix[75][174] * vector[75] +matrix[76][174] * vector[76] +matrix[77][174] * vector[77] +matrix[78][174] * vector[78] +matrix[79][174] * vector[79] +matrix[80][174] * vector[80] +matrix[81][174] * vector[81] +matrix[82][174] * vector[82] +matrix[83][174] * vector[83] +matrix[84][174] * vector[84] +matrix[85][174] * vector[85] +matrix[86][174] * vector[86] +matrix[87][174] * vector[87] +matrix[88][174] * vector[88] +matrix[89][174] * vector[89] +matrix[90][174] * vector[90] +matrix[91][174] * vector[91] +matrix[92][174] * vector[92] +matrix[93][174] * vector[93] +matrix[94][174] * vector[94] +matrix[95][174] * vector[95] +matrix[96][174] * vector[96] +matrix[97][174] * vector[97] +matrix[98][174] * vector[98] +matrix[99][174] * vector[99] +b[174];
assign result[175] = matrix[0][175] * vector[0] +matrix[1][175] * vector[1] +matrix[2][175] * vector[2] +matrix[3][175] * vector[3] +matrix[4][175] * vector[4] +matrix[5][175] * vector[5] +matrix[6][175] * vector[6] +matrix[7][175] * vector[7] +matrix[8][175] * vector[8] +matrix[9][175] * vector[9] +matrix[10][175] * vector[10] +matrix[11][175] * vector[11] +matrix[12][175] * vector[12] +matrix[13][175] * vector[13] +matrix[14][175] * vector[14] +matrix[15][175] * vector[15] +matrix[16][175] * vector[16] +matrix[17][175] * vector[17] +matrix[18][175] * vector[18] +matrix[19][175] * vector[19] +matrix[20][175] * vector[20] +matrix[21][175] * vector[21] +matrix[22][175] * vector[22] +matrix[23][175] * vector[23] +matrix[24][175] * vector[24] +matrix[25][175] * vector[25] +matrix[26][175] * vector[26] +matrix[27][175] * vector[27] +matrix[28][175] * vector[28] +matrix[29][175] * vector[29] +matrix[30][175] * vector[30] +matrix[31][175] * vector[31] +matrix[32][175] * vector[32] +matrix[33][175] * vector[33] +matrix[34][175] * vector[34] +matrix[35][175] * vector[35] +matrix[36][175] * vector[36] +matrix[37][175] * vector[37] +matrix[38][175] * vector[38] +matrix[39][175] * vector[39] +matrix[40][175] * vector[40] +matrix[41][175] * vector[41] +matrix[42][175] * vector[42] +matrix[43][175] * vector[43] +matrix[44][175] * vector[44] +matrix[45][175] * vector[45] +matrix[46][175] * vector[46] +matrix[47][175] * vector[47] +matrix[48][175] * vector[48] +matrix[49][175] * vector[49] +matrix[50][175] * vector[50] +matrix[51][175] * vector[51] +matrix[52][175] * vector[52] +matrix[53][175] * vector[53] +matrix[54][175] * vector[54] +matrix[55][175] * vector[55] +matrix[56][175] * vector[56] +matrix[57][175] * vector[57] +matrix[58][175] * vector[58] +matrix[59][175] * vector[59] +matrix[60][175] * vector[60] +matrix[61][175] * vector[61] +matrix[62][175] * vector[62] +matrix[63][175] * vector[63] +matrix[64][175] * vector[64] +matrix[65][175] * vector[65] +matrix[66][175] * vector[66] +matrix[67][175] * vector[67] +matrix[68][175] * vector[68] +matrix[69][175] * vector[69] +matrix[70][175] * vector[70] +matrix[71][175] * vector[71] +matrix[72][175] * vector[72] +matrix[73][175] * vector[73] +matrix[74][175] * vector[74] +matrix[75][175] * vector[75] +matrix[76][175] * vector[76] +matrix[77][175] * vector[77] +matrix[78][175] * vector[78] +matrix[79][175] * vector[79] +matrix[80][175] * vector[80] +matrix[81][175] * vector[81] +matrix[82][175] * vector[82] +matrix[83][175] * vector[83] +matrix[84][175] * vector[84] +matrix[85][175] * vector[85] +matrix[86][175] * vector[86] +matrix[87][175] * vector[87] +matrix[88][175] * vector[88] +matrix[89][175] * vector[89] +matrix[90][175] * vector[90] +matrix[91][175] * vector[91] +matrix[92][175] * vector[92] +matrix[93][175] * vector[93] +matrix[94][175] * vector[94] +matrix[95][175] * vector[95] +matrix[96][175] * vector[96] +matrix[97][175] * vector[97] +matrix[98][175] * vector[98] +matrix[99][175] * vector[99] +b[175];
assign result[176] = matrix[0][176] * vector[0] +matrix[1][176] * vector[1] +matrix[2][176] * vector[2] +matrix[3][176] * vector[3] +matrix[4][176] * vector[4] +matrix[5][176] * vector[5] +matrix[6][176] * vector[6] +matrix[7][176] * vector[7] +matrix[8][176] * vector[8] +matrix[9][176] * vector[9] +matrix[10][176] * vector[10] +matrix[11][176] * vector[11] +matrix[12][176] * vector[12] +matrix[13][176] * vector[13] +matrix[14][176] * vector[14] +matrix[15][176] * vector[15] +matrix[16][176] * vector[16] +matrix[17][176] * vector[17] +matrix[18][176] * vector[18] +matrix[19][176] * vector[19] +matrix[20][176] * vector[20] +matrix[21][176] * vector[21] +matrix[22][176] * vector[22] +matrix[23][176] * vector[23] +matrix[24][176] * vector[24] +matrix[25][176] * vector[25] +matrix[26][176] * vector[26] +matrix[27][176] * vector[27] +matrix[28][176] * vector[28] +matrix[29][176] * vector[29] +matrix[30][176] * vector[30] +matrix[31][176] * vector[31] +matrix[32][176] * vector[32] +matrix[33][176] * vector[33] +matrix[34][176] * vector[34] +matrix[35][176] * vector[35] +matrix[36][176] * vector[36] +matrix[37][176] * vector[37] +matrix[38][176] * vector[38] +matrix[39][176] * vector[39] +matrix[40][176] * vector[40] +matrix[41][176] * vector[41] +matrix[42][176] * vector[42] +matrix[43][176] * vector[43] +matrix[44][176] * vector[44] +matrix[45][176] * vector[45] +matrix[46][176] * vector[46] +matrix[47][176] * vector[47] +matrix[48][176] * vector[48] +matrix[49][176] * vector[49] +matrix[50][176] * vector[50] +matrix[51][176] * vector[51] +matrix[52][176] * vector[52] +matrix[53][176] * vector[53] +matrix[54][176] * vector[54] +matrix[55][176] * vector[55] +matrix[56][176] * vector[56] +matrix[57][176] * vector[57] +matrix[58][176] * vector[58] +matrix[59][176] * vector[59] +matrix[60][176] * vector[60] +matrix[61][176] * vector[61] +matrix[62][176] * vector[62] +matrix[63][176] * vector[63] +matrix[64][176] * vector[64] +matrix[65][176] * vector[65] +matrix[66][176] * vector[66] +matrix[67][176] * vector[67] +matrix[68][176] * vector[68] +matrix[69][176] * vector[69] +matrix[70][176] * vector[70] +matrix[71][176] * vector[71] +matrix[72][176] * vector[72] +matrix[73][176] * vector[73] +matrix[74][176] * vector[74] +matrix[75][176] * vector[75] +matrix[76][176] * vector[76] +matrix[77][176] * vector[77] +matrix[78][176] * vector[78] +matrix[79][176] * vector[79] +matrix[80][176] * vector[80] +matrix[81][176] * vector[81] +matrix[82][176] * vector[82] +matrix[83][176] * vector[83] +matrix[84][176] * vector[84] +matrix[85][176] * vector[85] +matrix[86][176] * vector[86] +matrix[87][176] * vector[87] +matrix[88][176] * vector[88] +matrix[89][176] * vector[89] +matrix[90][176] * vector[90] +matrix[91][176] * vector[91] +matrix[92][176] * vector[92] +matrix[93][176] * vector[93] +matrix[94][176] * vector[94] +matrix[95][176] * vector[95] +matrix[96][176] * vector[96] +matrix[97][176] * vector[97] +matrix[98][176] * vector[98] +matrix[99][176] * vector[99] +b[176];
assign result[177] = matrix[0][177] * vector[0] +matrix[1][177] * vector[1] +matrix[2][177] * vector[2] +matrix[3][177] * vector[3] +matrix[4][177] * vector[4] +matrix[5][177] * vector[5] +matrix[6][177] * vector[6] +matrix[7][177] * vector[7] +matrix[8][177] * vector[8] +matrix[9][177] * vector[9] +matrix[10][177] * vector[10] +matrix[11][177] * vector[11] +matrix[12][177] * vector[12] +matrix[13][177] * vector[13] +matrix[14][177] * vector[14] +matrix[15][177] * vector[15] +matrix[16][177] * vector[16] +matrix[17][177] * vector[17] +matrix[18][177] * vector[18] +matrix[19][177] * vector[19] +matrix[20][177] * vector[20] +matrix[21][177] * vector[21] +matrix[22][177] * vector[22] +matrix[23][177] * vector[23] +matrix[24][177] * vector[24] +matrix[25][177] * vector[25] +matrix[26][177] * vector[26] +matrix[27][177] * vector[27] +matrix[28][177] * vector[28] +matrix[29][177] * vector[29] +matrix[30][177] * vector[30] +matrix[31][177] * vector[31] +matrix[32][177] * vector[32] +matrix[33][177] * vector[33] +matrix[34][177] * vector[34] +matrix[35][177] * vector[35] +matrix[36][177] * vector[36] +matrix[37][177] * vector[37] +matrix[38][177] * vector[38] +matrix[39][177] * vector[39] +matrix[40][177] * vector[40] +matrix[41][177] * vector[41] +matrix[42][177] * vector[42] +matrix[43][177] * vector[43] +matrix[44][177] * vector[44] +matrix[45][177] * vector[45] +matrix[46][177] * vector[46] +matrix[47][177] * vector[47] +matrix[48][177] * vector[48] +matrix[49][177] * vector[49] +matrix[50][177] * vector[50] +matrix[51][177] * vector[51] +matrix[52][177] * vector[52] +matrix[53][177] * vector[53] +matrix[54][177] * vector[54] +matrix[55][177] * vector[55] +matrix[56][177] * vector[56] +matrix[57][177] * vector[57] +matrix[58][177] * vector[58] +matrix[59][177] * vector[59] +matrix[60][177] * vector[60] +matrix[61][177] * vector[61] +matrix[62][177] * vector[62] +matrix[63][177] * vector[63] +matrix[64][177] * vector[64] +matrix[65][177] * vector[65] +matrix[66][177] * vector[66] +matrix[67][177] * vector[67] +matrix[68][177] * vector[68] +matrix[69][177] * vector[69] +matrix[70][177] * vector[70] +matrix[71][177] * vector[71] +matrix[72][177] * vector[72] +matrix[73][177] * vector[73] +matrix[74][177] * vector[74] +matrix[75][177] * vector[75] +matrix[76][177] * vector[76] +matrix[77][177] * vector[77] +matrix[78][177] * vector[78] +matrix[79][177] * vector[79] +matrix[80][177] * vector[80] +matrix[81][177] * vector[81] +matrix[82][177] * vector[82] +matrix[83][177] * vector[83] +matrix[84][177] * vector[84] +matrix[85][177] * vector[85] +matrix[86][177] * vector[86] +matrix[87][177] * vector[87] +matrix[88][177] * vector[88] +matrix[89][177] * vector[89] +matrix[90][177] * vector[90] +matrix[91][177] * vector[91] +matrix[92][177] * vector[92] +matrix[93][177] * vector[93] +matrix[94][177] * vector[94] +matrix[95][177] * vector[95] +matrix[96][177] * vector[96] +matrix[97][177] * vector[97] +matrix[98][177] * vector[98] +matrix[99][177] * vector[99] +b[177];
assign result[178] = matrix[0][178] * vector[0] +matrix[1][178] * vector[1] +matrix[2][178] * vector[2] +matrix[3][178] * vector[3] +matrix[4][178] * vector[4] +matrix[5][178] * vector[5] +matrix[6][178] * vector[6] +matrix[7][178] * vector[7] +matrix[8][178] * vector[8] +matrix[9][178] * vector[9] +matrix[10][178] * vector[10] +matrix[11][178] * vector[11] +matrix[12][178] * vector[12] +matrix[13][178] * vector[13] +matrix[14][178] * vector[14] +matrix[15][178] * vector[15] +matrix[16][178] * vector[16] +matrix[17][178] * vector[17] +matrix[18][178] * vector[18] +matrix[19][178] * vector[19] +matrix[20][178] * vector[20] +matrix[21][178] * vector[21] +matrix[22][178] * vector[22] +matrix[23][178] * vector[23] +matrix[24][178] * vector[24] +matrix[25][178] * vector[25] +matrix[26][178] * vector[26] +matrix[27][178] * vector[27] +matrix[28][178] * vector[28] +matrix[29][178] * vector[29] +matrix[30][178] * vector[30] +matrix[31][178] * vector[31] +matrix[32][178] * vector[32] +matrix[33][178] * vector[33] +matrix[34][178] * vector[34] +matrix[35][178] * vector[35] +matrix[36][178] * vector[36] +matrix[37][178] * vector[37] +matrix[38][178] * vector[38] +matrix[39][178] * vector[39] +matrix[40][178] * vector[40] +matrix[41][178] * vector[41] +matrix[42][178] * vector[42] +matrix[43][178] * vector[43] +matrix[44][178] * vector[44] +matrix[45][178] * vector[45] +matrix[46][178] * vector[46] +matrix[47][178] * vector[47] +matrix[48][178] * vector[48] +matrix[49][178] * vector[49] +matrix[50][178] * vector[50] +matrix[51][178] * vector[51] +matrix[52][178] * vector[52] +matrix[53][178] * vector[53] +matrix[54][178] * vector[54] +matrix[55][178] * vector[55] +matrix[56][178] * vector[56] +matrix[57][178] * vector[57] +matrix[58][178] * vector[58] +matrix[59][178] * vector[59] +matrix[60][178] * vector[60] +matrix[61][178] * vector[61] +matrix[62][178] * vector[62] +matrix[63][178] * vector[63] +matrix[64][178] * vector[64] +matrix[65][178] * vector[65] +matrix[66][178] * vector[66] +matrix[67][178] * vector[67] +matrix[68][178] * vector[68] +matrix[69][178] * vector[69] +matrix[70][178] * vector[70] +matrix[71][178] * vector[71] +matrix[72][178] * vector[72] +matrix[73][178] * vector[73] +matrix[74][178] * vector[74] +matrix[75][178] * vector[75] +matrix[76][178] * vector[76] +matrix[77][178] * vector[77] +matrix[78][178] * vector[78] +matrix[79][178] * vector[79] +matrix[80][178] * vector[80] +matrix[81][178] * vector[81] +matrix[82][178] * vector[82] +matrix[83][178] * vector[83] +matrix[84][178] * vector[84] +matrix[85][178] * vector[85] +matrix[86][178] * vector[86] +matrix[87][178] * vector[87] +matrix[88][178] * vector[88] +matrix[89][178] * vector[89] +matrix[90][178] * vector[90] +matrix[91][178] * vector[91] +matrix[92][178] * vector[92] +matrix[93][178] * vector[93] +matrix[94][178] * vector[94] +matrix[95][178] * vector[95] +matrix[96][178] * vector[96] +matrix[97][178] * vector[97] +matrix[98][178] * vector[98] +matrix[99][178] * vector[99] +b[178];
assign result[179] = matrix[0][179] * vector[0] +matrix[1][179] * vector[1] +matrix[2][179] * vector[2] +matrix[3][179] * vector[3] +matrix[4][179] * vector[4] +matrix[5][179] * vector[5] +matrix[6][179] * vector[6] +matrix[7][179] * vector[7] +matrix[8][179] * vector[8] +matrix[9][179] * vector[9] +matrix[10][179] * vector[10] +matrix[11][179] * vector[11] +matrix[12][179] * vector[12] +matrix[13][179] * vector[13] +matrix[14][179] * vector[14] +matrix[15][179] * vector[15] +matrix[16][179] * vector[16] +matrix[17][179] * vector[17] +matrix[18][179] * vector[18] +matrix[19][179] * vector[19] +matrix[20][179] * vector[20] +matrix[21][179] * vector[21] +matrix[22][179] * vector[22] +matrix[23][179] * vector[23] +matrix[24][179] * vector[24] +matrix[25][179] * vector[25] +matrix[26][179] * vector[26] +matrix[27][179] * vector[27] +matrix[28][179] * vector[28] +matrix[29][179] * vector[29] +matrix[30][179] * vector[30] +matrix[31][179] * vector[31] +matrix[32][179] * vector[32] +matrix[33][179] * vector[33] +matrix[34][179] * vector[34] +matrix[35][179] * vector[35] +matrix[36][179] * vector[36] +matrix[37][179] * vector[37] +matrix[38][179] * vector[38] +matrix[39][179] * vector[39] +matrix[40][179] * vector[40] +matrix[41][179] * vector[41] +matrix[42][179] * vector[42] +matrix[43][179] * vector[43] +matrix[44][179] * vector[44] +matrix[45][179] * vector[45] +matrix[46][179] * vector[46] +matrix[47][179] * vector[47] +matrix[48][179] * vector[48] +matrix[49][179] * vector[49] +matrix[50][179] * vector[50] +matrix[51][179] * vector[51] +matrix[52][179] * vector[52] +matrix[53][179] * vector[53] +matrix[54][179] * vector[54] +matrix[55][179] * vector[55] +matrix[56][179] * vector[56] +matrix[57][179] * vector[57] +matrix[58][179] * vector[58] +matrix[59][179] * vector[59] +matrix[60][179] * vector[60] +matrix[61][179] * vector[61] +matrix[62][179] * vector[62] +matrix[63][179] * vector[63] +matrix[64][179] * vector[64] +matrix[65][179] * vector[65] +matrix[66][179] * vector[66] +matrix[67][179] * vector[67] +matrix[68][179] * vector[68] +matrix[69][179] * vector[69] +matrix[70][179] * vector[70] +matrix[71][179] * vector[71] +matrix[72][179] * vector[72] +matrix[73][179] * vector[73] +matrix[74][179] * vector[74] +matrix[75][179] * vector[75] +matrix[76][179] * vector[76] +matrix[77][179] * vector[77] +matrix[78][179] * vector[78] +matrix[79][179] * vector[79] +matrix[80][179] * vector[80] +matrix[81][179] * vector[81] +matrix[82][179] * vector[82] +matrix[83][179] * vector[83] +matrix[84][179] * vector[84] +matrix[85][179] * vector[85] +matrix[86][179] * vector[86] +matrix[87][179] * vector[87] +matrix[88][179] * vector[88] +matrix[89][179] * vector[89] +matrix[90][179] * vector[90] +matrix[91][179] * vector[91] +matrix[92][179] * vector[92] +matrix[93][179] * vector[93] +matrix[94][179] * vector[94] +matrix[95][179] * vector[95] +matrix[96][179] * vector[96] +matrix[97][179] * vector[97] +matrix[98][179] * vector[98] +matrix[99][179] * vector[99] +b[179];
assign result[180] = matrix[0][180] * vector[0] +matrix[1][180] * vector[1] +matrix[2][180] * vector[2] +matrix[3][180] * vector[3] +matrix[4][180] * vector[4] +matrix[5][180] * vector[5] +matrix[6][180] * vector[6] +matrix[7][180] * vector[7] +matrix[8][180] * vector[8] +matrix[9][180] * vector[9] +matrix[10][180] * vector[10] +matrix[11][180] * vector[11] +matrix[12][180] * vector[12] +matrix[13][180] * vector[13] +matrix[14][180] * vector[14] +matrix[15][180] * vector[15] +matrix[16][180] * vector[16] +matrix[17][180] * vector[17] +matrix[18][180] * vector[18] +matrix[19][180] * vector[19] +matrix[20][180] * vector[20] +matrix[21][180] * vector[21] +matrix[22][180] * vector[22] +matrix[23][180] * vector[23] +matrix[24][180] * vector[24] +matrix[25][180] * vector[25] +matrix[26][180] * vector[26] +matrix[27][180] * vector[27] +matrix[28][180] * vector[28] +matrix[29][180] * vector[29] +matrix[30][180] * vector[30] +matrix[31][180] * vector[31] +matrix[32][180] * vector[32] +matrix[33][180] * vector[33] +matrix[34][180] * vector[34] +matrix[35][180] * vector[35] +matrix[36][180] * vector[36] +matrix[37][180] * vector[37] +matrix[38][180] * vector[38] +matrix[39][180] * vector[39] +matrix[40][180] * vector[40] +matrix[41][180] * vector[41] +matrix[42][180] * vector[42] +matrix[43][180] * vector[43] +matrix[44][180] * vector[44] +matrix[45][180] * vector[45] +matrix[46][180] * vector[46] +matrix[47][180] * vector[47] +matrix[48][180] * vector[48] +matrix[49][180] * vector[49] +matrix[50][180] * vector[50] +matrix[51][180] * vector[51] +matrix[52][180] * vector[52] +matrix[53][180] * vector[53] +matrix[54][180] * vector[54] +matrix[55][180] * vector[55] +matrix[56][180] * vector[56] +matrix[57][180] * vector[57] +matrix[58][180] * vector[58] +matrix[59][180] * vector[59] +matrix[60][180] * vector[60] +matrix[61][180] * vector[61] +matrix[62][180] * vector[62] +matrix[63][180] * vector[63] +matrix[64][180] * vector[64] +matrix[65][180] * vector[65] +matrix[66][180] * vector[66] +matrix[67][180] * vector[67] +matrix[68][180] * vector[68] +matrix[69][180] * vector[69] +matrix[70][180] * vector[70] +matrix[71][180] * vector[71] +matrix[72][180] * vector[72] +matrix[73][180] * vector[73] +matrix[74][180] * vector[74] +matrix[75][180] * vector[75] +matrix[76][180] * vector[76] +matrix[77][180] * vector[77] +matrix[78][180] * vector[78] +matrix[79][180] * vector[79] +matrix[80][180] * vector[80] +matrix[81][180] * vector[81] +matrix[82][180] * vector[82] +matrix[83][180] * vector[83] +matrix[84][180] * vector[84] +matrix[85][180] * vector[85] +matrix[86][180] * vector[86] +matrix[87][180] * vector[87] +matrix[88][180] * vector[88] +matrix[89][180] * vector[89] +matrix[90][180] * vector[90] +matrix[91][180] * vector[91] +matrix[92][180] * vector[92] +matrix[93][180] * vector[93] +matrix[94][180] * vector[94] +matrix[95][180] * vector[95] +matrix[96][180] * vector[96] +matrix[97][180] * vector[97] +matrix[98][180] * vector[98] +matrix[99][180] * vector[99] +b[180];
assign result[181] = matrix[0][181] * vector[0] +matrix[1][181] * vector[1] +matrix[2][181] * vector[2] +matrix[3][181] * vector[3] +matrix[4][181] * vector[4] +matrix[5][181] * vector[5] +matrix[6][181] * vector[6] +matrix[7][181] * vector[7] +matrix[8][181] * vector[8] +matrix[9][181] * vector[9] +matrix[10][181] * vector[10] +matrix[11][181] * vector[11] +matrix[12][181] * vector[12] +matrix[13][181] * vector[13] +matrix[14][181] * vector[14] +matrix[15][181] * vector[15] +matrix[16][181] * vector[16] +matrix[17][181] * vector[17] +matrix[18][181] * vector[18] +matrix[19][181] * vector[19] +matrix[20][181] * vector[20] +matrix[21][181] * vector[21] +matrix[22][181] * vector[22] +matrix[23][181] * vector[23] +matrix[24][181] * vector[24] +matrix[25][181] * vector[25] +matrix[26][181] * vector[26] +matrix[27][181] * vector[27] +matrix[28][181] * vector[28] +matrix[29][181] * vector[29] +matrix[30][181] * vector[30] +matrix[31][181] * vector[31] +matrix[32][181] * vector[32] +matrix[33][181] * vector[33] +matrix[34][181] * vector[34] +matrix[35][181] * vector[35] +matrix[36][181] * vector[36] +matrix[37][181] * vector[37] +matrix[38][181] * vector[38] +matrix[39][181] * vector[39] +matrix[40][181] * vector[40] +matrix[41][181] * vector[41] +matrix[42][181] * vector[42] +matrix[43][181] * vector[43] +matrix[44][181] * vector[44] +matrix[45][181] * vector[45] +matrix[46][181] * vector[46] +matrix[47][181] * vector[47] +matrix[48][181] * vector[48] +matrix[49][181] * vector[49] +matrix[50][181] * vector[50] +matrix[51][181] * vector[51] +matrix[52][181] * vector[52] +matrix[53][181] * vector[53] +matrix[54][181] * vector[54] +matrix[55][181] * vector[55] +matrix[56][181] * vector[56] +matrix[57][181] * vector[57] +matrix[58][181] * vector[58] +matrix[59][181] * vector[59] +matrix[60][181] * vector[60] +matrix[61][181] * vector[61] +matrix[62][181] * vector[62] +matrix[63][181] * vector[63] +matrix[64][181] * vector[64] +matrix[65][181] * vector[65] +matrix[66][181] * vector[66] +matrix[67][181] * vector[67] +matrix[68][181] * vector[68] +matrix[69][181] * vector[69] +matrix[70][181] * vector[70] +matrix[71][181] * vector[71] +matrix[72][181] * vector[72] +matrix[73][181] * vector[73] +matrix[74][181] * vector[74] +matrix[75][181] * vector[75] +matrix[76][181] * vector[76] +matrix[77][181] * vector[77] +matrix[78][181] * vector[78] +matrix[79][181] * vector[79] +matrix[80][181] * vector[80] +matrix[81][181] * vector[81] +matrix[82][181] * vector[82] +matrix[83][181] * vector[83] +matrix[84][181] * vector[84] +matrix[85][181] * vector[85] +matrix[86][181] * vector[86] +matrix[87][181] * vector[87] +matrix[88][181] * vector[88] +matrix[89][181] * vector[89] +matrix[90][181] * vector[90] +matrix[91][181] * vector[91] +matrix[92][181] * vector[92] +matrix[93][181] * vector[93] +matrix[94][181] * vector[94] +matrix[95][181] * vector[95] +matrix[96][181] * vector[96] +matrix[97][181] * vector[97] +matrix[98][181] * vector[98] +matrix[99][181] * vector[99] +b[181];
assign result[182] = matrix[0][182] * vector[0] +matrix[1][182] * vector[1] +matrix[2][182] * vector[2] +matrix[3][182] * vector[3] +matrix[4][182] * vector[4] +matrix[5][182] * vector[5] +matrix[6][182] * vector[6] +matrix[7][182] * vector[7] +matrix[8][182] * vector[8] +matrix[9][182] * vector[9] +matrix[10][182] * vector[10] +matrix[11][182] * vector[11] +matrix[12][182] * vector[12] +matrix[13][182] * vector[13] +matrix[14][182] * vector[14] +matrix[15][182] * vector[15] +matrix[16][182] * vector[16] +matrix[17][182] * vector[17] +matrix[18][182] * vector[18] +matrix[19][182] * vector[19] +matrix[20][182] * vector[20] +matrix[21][182] * vector[21] +matrix[22][182] * vector[22] +matrix[23][182] * vector[23] +matrix[24][182] * vector[24] +matrix[25][182] * vector[25] +matrix[26][182] * vector[26] +matrix[27][182] * vector[27] +matrix[28][182] * vector[28] +matrix[29][182] * vector[29] +matrix[30][182] * vector[30] +matrix[31][182] * vector[31] +matrix[32][182] * vector[32] +matrix[33][182] * vector[33] +matrix[34][182] * vector[34] +matrix[35][182] * vector[35] +matrix[36][182] * vector[36] +matrix[37][182] * vector[37] +matrix[38][182] * vector[38] +matrix[39][182] * vector[39] +matrix[40][182] * vector[40] +matrix[41][182] * vector[41] +matrix[42][182] * vector[42] +matrix[43][182] * vector[43] +matrix[44][182] * vector[44] +matrix[45][182] * vector[45] +matrix[46][182] * vector[46] +matrix[47][182] * vector[47] +matrix[48][182] * vector[48] +matrix[49][182] * vector[49] +matrix[50][182] * vector[50] +matrix[51][182] * vector[51] +matrix[52][182] * vector[52] +matrix[53][182] * vector[53] +matrix[54][182] * vector[54] +matrix[55][182] * vector[55] +matrix[56][182] * vector[56] +matrix[57][182] * vector[57] +matrix[58][182] * vector[58] +matrix[59][182] * vector[59] +matrix[60][182] * vector[60] +matrix[61][182] * vector[61] +matrix[62][182] * vector[62] +matrix[63][182] * vector[63] +matrix[64][182] * vector[64] +matrix[65][182] * vector[65] +matrix[66][182] * vector[66] +matrix[67][182] * vector[67] +matrix[68][182] * vector[68] +matrix[69][182] * vector[69] +matrix[70][182] * vector[70] +matrix[71][182] * vector[71] +matrix[72][182] * vector[72] +matrix[73][182] * vector[73] +matrix[74][182] * vector[74] +matrix[75][182] * vector[75] +matrix[76][182] * vector[76] +matrix[77][182] * vector[77] +matrix[78][182] * vector[78] +matrix[79][182] * vector[79] +matrix[80][182] * vector[80] +matrix[81][182] * vector[81] +matrix[82][182] * vector[82] +matrix[83][182] * vector[83] +matrix[84][182] * vector[84] +matrix[85][182] * vector[85] +matrix[86][182] * vector[86] +matrix[87][182] * vector[87] +matrix[88][182] * vector[88] +matrix[89][182] * vector[89] +matrix[90][182] * vector[90] +matrix[91][182] * vector[91] +matrix[92][182] * vector[92] +matrix[93][182] * vector[93] +matrix[94][182] * vector[94] +matrix[95][182] * vector[95] +matrix[96][182] * vector[96] +matrix[97][182] * vector[97] +matrix[98][182] * vector[98] +matrix[99][182] * vector[99] +b[182];
assign result[183] = matrix[0][183] * vector[0] +matrix[1][183] * vector[1] +matrix[2][183] * vector[2] +matrix[3][183] * vector[3] +matrix[4][183] * vector[4] +matrix[5][183] * vector[5] +matrix[6][183] * vector[6] +matrix[7][183] * vector[7] +matrix[8][183] * vector[8] +matrix[9][183] * vector[9] +matrix[10][183] * vector[10] +matrix[11][183] * vector[11] +matrix[12][183] * vector[12] +matrix[13][183] * vector[13] +matrix[14][183] * vector[14] +matrix[15][183] * vector[15] +matrix[16][183] * vector[16] +matrix[17][183] * vector[17] +matrix[18][183] * vector[18] +matrix[19][183] * vector[19] +matrix[20][183] * vector[20] +matrix[21][183] * vector[21] +matrix[22][183] * vector[22] +matrix[23][183] * vector[23] +matrix[24][183] * vector[24] +matrix[25][183] * vector[25] +matrix[26][183] * vector[26] +matrix[27][183] * vector[27] +matrix[28][183] * vector[28] +matrix[29][183] * vector[29] +matrix[30][183] * vector[30] +matrix[31][183] * vector[31] +matrix[32][183] * vector[32] +matrix[33][183] * vector[33] +matrix[34][183] * vector[34] +matrix[35][183] * vector[35] +matrix[36][183] * vector[36] +matrix[37][183] * vector[37] +matrix[38][183] * vector[38] +matrix[39][183] * vector[39] +matrix[40][183] * vector[40] +matrix[41][183] * vector[41] +matrix[42][183] * vector[42] +matrix[43][183] * vector[43] +matrix[44][183] * vector[44] +matrix[45][183] * vector[45] +matrix[46][183] * vector[46] +matrix[47][183] * vector[47] +matrix[48][183] * vector[48] +matrix[49][183] * vector[49] +matrix[50][183] * vector[50] +matrix[51][183] * vector[51] +matrix[52][183] * vector[52] +matrix[53][183] * vector[53] +matrix[54][183] * vector[54] +matrix[55][183] * vector[55] +matrix[56][183] * vector[56] +matrix[57][183] * vector[57] +matrix[58][183] * vector[58] +matrix[59][183] * vector[59] +matrix[60][183] * vector[60] +matrix[61][183] * vector[61] +matrix[62][183] * vector[62] +matrix[63][183] * vector[63] +matrix[64][183] * vector[64] +matrix[65][183] * vector[65] +matrix[66][183] * vector[66] +matrix[67][183] * vector[67] +matrix[68][183] * vector[68] +matrix[69][183] * vector[69] +matrix[70][183] * vector[70] +matrix[71][183] * vector[71] +matrix[72][183] * vector[72] +matrix[73][183] * vector[73] +matrix[74][183] * vector[74] +matrix[75][183] * vector[75] +matrix[76][183] * vector[76] +matrix[77][183] * vector[77] +matrix[78][183] * vector[78] +matrix[79][183] * vector[79] +matrix[80][183] * vector[80] +matrix[81][183] * vector[81] +matrix[82][183] * vector[82] +matrix[83][183] * vector[83] +matrix[84][183] * vector[84] +matrix[85][183] * vector[85] +matrix[86][183] * vector[86] +matrix[87][183] * vector[87] +matrix[88][183] * vector[88] +matrix[89][183] * vector[89] +matrix[90][183] * vector[90] +matrix[91][183] * vector[91] +matrix[92][183] * vector[92] +matrix[93][183] * vector[93] +matrix[94][183] * vector[94] +matrix[95][183] * vector[95] +matrix[96][183] * vector[96] +matrix[97][183] * vector[97] +matrix[98][183] * vector[98] +matrix[99][183] * vector[99] +b[183];
assign result[184] = matrix[0][184] * vector[0] +matrix[1][184] * vector[1] +matrix[2][184] * vector[2] +matrix[3][184] * vector[3] +matrix[4][184] * vector[4] +matrix[5][184] * vector[5] +matrix[6][184] * vector[6] +matrix[7][184] * vector[7] +matrix[8][184] * vector[8] +matrix[9][184] * vector[9] +matrix[10][184] * vector[10] +matrix[11][184] * vector[11] +matrix[12][184] * vector[12] +matrix[13][184] * vector[13] +matrix[14][184] * vector[14] +matrix[15][184] * vector[15] +matrix[16][184] * vector[16] +matrix[17][184] * vector[17] +matrix[18][184] * vector[18] +matrix[19][184] * vector[19] +matrix[20][184] * vector[20] +matrix[21][184] * vector[21] +matrix[22][184] * vector[22] +matrix[23][184] * vector[23] +matrix[24][184] * vector[24] +matrix[25][184] * vector[25] +matrix[26][184] * vector[26] +matrix[27][184] * vector[27] +matrix[28][184] * vector[28] +matrix[29][184] * vector[29] +matrix[30][184] * vector[30] +matrix[31][184] * vector[31] +matrix[32][184] * vector[32] +matrix[33][184] * vector[33] +matrix[34][184] * vector[34] +matrix[35][184] * vector[35] +matrix[36][184] * vector[36] +matrix[37][184] * vector[37] +matrix[38][184] * vector[38] +matrix[39][184] * vector[39] +matrix[40][184] * vector[40] +matrix[41][184] * vector[41] +matrix[42][184] * vector[42] +matrix[43][184] * vector[43] +matrix[44][184] * vector[44] +matrix[45][184] * vector[45] +matrix[46][184] * vector[46] +matrix[47][184] * vector[47] +matrix[48][184] * vector[48] +matrix[49][184] * vector[49] +matrix[50][184] * vector[50] +matrix[51][184] * vector[51] +matrix[52][184] * vector[52] +matrix[53][184] * vector[53] +matrix[54][184] * vector[54] +matrix[55][184] * vector[55] +matrix[56][184] * vector[56] +matrix[57][184] * vector[57] +matrix[58][184] * vector[58] +matrix[59][184] * vector[59] +matrix[60][184] * vector[60] +matrix[61][184] * vector[61] +matrix[62][184] * vector[62] +matrix[63][184] * vector[63] +matrix[64][184] * vector[64] +matrix[65][184] * vector[65] +matrix[66][184] * vector[66] +matrix[67][184] * vector[67] +matrix[68][184] * vector[68] +matrix[69][184] * vector[69] +matrix[70][184] * vector[70] +matrix[71][184] * vector[71] +matrix[72][184] * vector[72] +matrix[73][184] * vector[73] +matrix[74][184] * vector[74] +matrix[75][184] * vector[75] +matrix[76][184] * vector[76] +matrix[77][184] * vector[77] +matrix[78][184] * vector[78] +matrix[79][184] * vector[79] +matrix[80][184] * vector[80] +matrix[81][184] * vector[81] +matrix[82][184] * vector[82] +matrix[83][184] * vector[83] +matrix[84][184] * vector[84] +matrix[85][184] * vector[85] +matrix[86][184] * vector[86] +matrix[87][184] * vector[87] +matrix[88][184] * vector[88] +matrix[89][184] * vector[89] +matrix[90][184] * vector[90] +matrix[91][184] * vector[91] +matrix[92][184] * vector[92] +matrix[93][184] * vector[93] +matrix[94][184] * vector[94] +matrix[95][184] * vector[95] +matrix[96][184] * vector[96] +matrix[97][184] * vector[97] +matrix[98][184] * vector[98] +matrix[99][184] * vector[99] +b[184];
assign result[185] = matrix[0][185] * vector[0] +matrix[1][185] * vector[1] +matrix[2][185] * vector[2] +matrix[3][185] * vector[3] +matrix[4][185] * vector[4] +matrix[5][185] * vector[5] +matrix[6][185] * vector[6] +matrix[7][185] * vector[7] +matrix[8][185] * vector[8] +matrix[9][185] * vector[9] +matrix[10][185] * vector[10] +matrix[11][185] * vector[11] +matrix[12][185] * vector[12] +matrix[13][185] * vector[13] +matrix[14][185] * vector[14] +matrix[15][185] * vector[15] +matrix[16][185] * vector[16] +matrix[17][185] * vector[17] +matrix[18][185] * vector[18] +matrix[19][185] * vector[19] +matrix[20][185] * vector[20] +matrix[21][185] * vector[21] +matrix[22][185] * vector[22] +matrix[23][185] * vector[23] +matrix[24][185] * vector[24] +matrix[25][185] * vector[25] +matrix[26][185] * vector[26] +matrix[27][185] * vector[27] +matrix[28][185] * vector[28] +matrix[29][185] * vector[29] +matrix[30][185] * vector[30] +matrix[31][185] * vector[31] +matrix[32][185] * vector[32] +matrix[33][185] * vector[33] +matrix[34][185] * vector[34] +matrix[35][185] * vector[35] +matrix[36][185] * vector[36] +matrix[37][185] * vector[37] +matrix[38][185] * vector[38] +matrix[39][185] * vector[39] +matrix[40][185] * vector[40] +matrix[41][185] * vector[41] +matrix[42][185] * vector[42] +matrix[43][185] * vector[43] +matrix[44][185] * vector[44] +matrix[45][185] * vector[45] +matrix[46][185] * vector[46] +matrix[47][185] * vector[47] +matrix[48][185] * vector[48] +matrix[49][185] * vector[49] +matrix[50][185] * vector[50] +matrix[51][185] * vector[51] +matrix[52][185] * vector[52] +matrix[53][185] * vector[53] +matrix[54][185] * vector[54] +matrix[55][185] * vector[55] +matrix[56][185] * vector[56] +matrix[57][185] * vector[57] +matrix[58][185] * vector[58] +matrix[59][185] * vector[59] +matrix[60][185] * vector[60] +matrix[61][185] * vector[61] +matrix[62][185] * vector[62] +matrix[63][185] * vector[63] +matrix[64][185] * vector[64] +matrix[65][185] * vector[65] +matrix[66][185] * vector[66] +matrix[67][185] * vector[67] +matrix[68][185] * vector[68] +matrix[69][185] * vector[69] +matrix[70][185] * vector[70] +matrix[71][185] * vector[71] +matrix[72][185] * vector[72] +matrix[73][185] * vector[73] +matrix[74][185] * vector[74] +matrix[75][185] * vector[75] +matrix[76][185] * vector[76] +matrix[77][185] * vector[77] +matrix[78][185] * vector[78] +matrix[79][185] * vector[79] +matrix[80][185] * vector[80] +matrix[81][185] * vector[81] +matrix[82][185] * vector[82] +matrix[83][185] * vector[83] +matrix[84][185] * vector[84] +matrix[85][185] * vector[85] +matrix[86][185] * vector[86] +matrix[87][185] * vector[87] +matrix[88][185] * vector[88] +matrix[89][185] * vector[89] +matrix[90][185] * vector[90] +matrix[91][185] * vector[91] +matrix[92][185] * vector[92] +matrix[93][185] * vector[93] +matrix[94][185] * vector[94] +matrix[95][185] * vector[95] +matrix[96][185] * vector[96] +matrix[97][185] * vector[97] +matrix[98][185] * vector[98] +matrix[99][185] * vector[99] +b[185];
assign result[186] = matrix[0][186] * vector[0] +matrix[1][186] * vector[1] +matrix[2][186] * vector[2] +matrix[3][186] * vector[3] +matrix[4][186] * vector[4] +matrix[5][186] * vector[5] +matrix[6][186] * vector[6] +matrix[7][186] * vector[7] +matrix[8][186] * vector[8] +matrix[9][186] * vector[9] +matrix[10][186] * vector[10] +matrix[11][186] * vector[11] +matrix[12][186] * vector[12] +matrix[13][186] * vector[13] +matrix[14][186] * vector[14] +matrix[15][186] * vector[15] +matrix[16][186] * vector[16] +matrix[17][186] * vector[17] +matrix[18][186] * vector[18] +matrix[19][186] * vector[19] +matrix[20][186] * vector[20] +matrix[21][186] * vector[21] +matrix[22][186] * vector[22] +matrix[23][186] * vector[23] +matrix[24][186] * vector[24] +matrix[25][186] * vector[25] +matrix[26][186] * vector[26] +matrix[27][186] * vector[27] +matrix[28][186] * vector[28] +matrix[29][186] * vector[29] +matrix[30][186] * vector[30] +matrix[31][186] * vector[31] +matrix[32][186] * vector[32] +matrix[33][186] * vector[33] +matrix[34][186] * vector[34] +matrix[35][186] * vector[35] +matrix[36][186] * vector[36] +matrix[37][186] * vector[37] +matrix[38][186] * vector[38] +matrix[39][186] * vector[39] +matrix[40][186] * vector[40] +matrix[41][186] * vector[41] +matrix[42][186] * vector[42] +matrix[43][186] * vector[43] +matrix[44][186] * vector[44] +matrix[45][186] * vector[45] +matrix[46][186] * vector[46] +matrix[47][186] * vector[47] +matrix[48][186] * vector[48] +matrix[49][186] * vector[49] +matrix[50][186] * vector[50] +matrix[51][186] * vector[51] +matrix[52][186] * vector[52] +matrix[53][186] * vector[53] +matrix[54][186] * vector[54] +matrix[55][186] * vector[55] +matrix[56][186] * vector[56] +matrix[57][186] * vector[57] +matrix[58][186] * vector[58] +matrix[59][186] * vector[59] +matrix[60][186] * vector[60] +matrix[61][186] * vector[61] +matrix[62][186] * vector[62] +matrix[63][186] * vector[63] +matrix[64][186] * vector[64] +matrix[65][186] * vector[65] +matrix[66][186] * vector[66] +matrix[67][186] * vector[67] +matrix[68][186] * vector[68] +matrix[69][186] * vector[69] +matrix[70][186] * vector[70] +matrix[71][186] * vector[71] +matrix[72][186] * vector[72] +matrix[73][186] * vector[73] +matrix[74][186] * vector[74] +matrix[75][186] * vector[75] +matrix[76][186] * vector[76] +matrix[77][186] * vector[77] +matrix[78][186] * vector[78] +matrix[79][186] * vector[79] +matrix[80][186] * vector[80] +matrix[81][186] * vector[81] +matrix[82][186] * vector[82] +matrix[83][186] * vector[83] +matrix[84][186] * vector[84] +matrix[85][186] * vector[85] +matrix[86][186] * vector[86] +matrix[87][186] * vector[87] +matrix[88][186] * vector[88] +matrix[89][186] * vector[89] +matrix[90][186] * vector[90] +matrix[91][186] * vector[91] +matrix[92][186] * vector[92] +matrix[93][186] * vector[93] +matrix[94][186] * vector[94] +matrix[95][186] * vector[95] +matrix[96][186] * vector[96] +matrix[97][186] * vector[97] +matrix[98][186] * vector[98] +matrix[99][186] * vector[99] +b[186];
assign result[187] = matrix[0][187] * vector[0] +matrix[1][187] * vector[1] +matrix[2][187] * vector[2] +matrix[3][187] * vector[3] +matrix[4][187] * vector[4] +matrix[5][187] * vector[5] +matrix[6][187] * vector[6] +matrix[7][187] * vector[7] +matrix[8][187] * vector[8] +matrix[9][187] * vector[9] +matrix[10][187] * vector[10] +matrix[11][187] * vector[11] +matrix[12][187] * vector[12] +matrix[13][187] * vector[13] +matrix[14][187] * vector[14] +matrix[15][187] * vector[15] +matrix[16][187] * vector[16] +matrix[17][187] * vector[17] +matrix[18][187] * vector[18] +matrix[19][187] * vector[19] +matrix[20][187] * vector[20] +matrix[21][187] * vector[21] +matrix[22][187] * vector[22] +matrix[23][187] * vector[23] +matrix[24][187] * vector[24] +matrix[25][187] * vector[25] +matrix[26][187] * vector[26] +matrix[27][187] * vector[27] +matrix[28][187] * vector[28] +matrix[29][187] * vector[29] +matrix[30][187] * vector[30] +matrix[31][187] * vector[31] +matrix[32][187] * vector[32] +matrix[33][187] * vector[33] +matrix[34][187] * vector[34] +matrix[35][187] * vector[35] +matrix[36][187] * vector[36] +matrix[37][187] * vector[37] +matrix[38][187] * vector[38] +matrix[39][187] * vector[39] +matrix[40][187] * vector[40] +matrix[41][187] * vector[41] +matrix[42][187] * vector[42] +matrix[43][187] * vector[43] +matrix[44][187] * vector[44] +matrix[45][187] * vector[45] +matrix[46][187] * vector[46] +matrix[47][187] * vector[47] +matrix[48][187] * vector[48] +matrix[49][187] * vector[49] +matrix[50][187] * vector[50] +matrix[51][187] * vector[51] +matrix[52][187] * vector[52] +matrix[53][187] * vector[53] +matrix[54][187] * vector[54] +matrix[55][187] * vector[55] +matrix[56][187] * vector[56] +matrix[57][187] * vector[57] +matrix[58][187] * vector[58] +matrix[59][187] * vector[59] +matrix[60][187] * vector[60] +matrix[61][187] * vector[61] +matrix[62][187] * vector[62] +matrix[63][187] * vector[63] +matrix[64][187] * vector[64] +matrix[65][187] * vector[65] +matrix[66][187] * vector[66] +matrix[67][187] * vector[67] +matrix[68][187] * vector[68] +matrix[69][187] * vector[69] +matrix[70][187] * vector[70] +matrix[71][187] * vector[71] +matrix[72][187] * vector[72] +matrix[73][187] * vector[73] +matrix[74][187] * vector[74] +matrix[75][187] * vector[75] +matrix[76][187] * vector[76] +matrix[77][187] * vector[77] +matrix[78][187] * vector[78] +matrix[79][187] * vector[79] +matrix[80][187] * vector[80] +matrix[81][187] * vector[81] +matrix[82][187] * vector[82] +matrix[83][187] * vector[83] +matrix[84][187] * vector[84] +matrix[85][187] * vector[85] +matrix[86][187] * vector[86] +matrix[87][187] * vector[87] +matrix[88][187] * vector[88] +matrix[89][187] * vector[89] +matrix[90][187] * vector[90] +matrix[91][187] * vector[91] +matrix[92][187] * vector[92] +matrix[93][187] * vector[93] +matrix[94][187] * vector[94] +matrix[95][187] * vector[95] +matrix[96][187] * vector[96] +matrix[97][187] * vector[97] +matrix[98][187] * vector[98] +matrix[99][187] * vector[99] +b[187];
assign result[188] = matrix[0][188] * vector[0] +matrix[1][188] * vector[1] +matrix[2][188] * vector[2] +matrix[3][188] * vector[3] +matrix[4][188] * vector[4] +matrix[5][188] * vector[5] +matrix[6][188] * vector[6] +matrix[7][188] * vector[7] +matrix[8][188] * vector[8] +matrix[9][188] * vector[9] +matrix[10][188] * vector[10] +matrix[11][188] * vector[11] +matrix[12][188] * vector[12] +matrix[13][188] * vector[13] +matrix[14][188] * vector[14] +matrix[15][188] * vector[15] +matrix[16][188] * vector[16] +matrix[17][188] * vector[17] +matrix[18][188] * vector[18] +matrix[19][188] * vector[19] +matrix[20][188] * vector[20] +matrix[21][188] * vector[21] +matrix[22][188] * vector[22] +matrix[23][188] * vector[23] +matrix[24][188] * vector[24] +matrix[25][188] * vector[25] +matrix[26][188] * vector[26] +matrix[27][188] * vector[27] +matrix[28][188] * vector[28] +matrix[29][188] * vector[29] +matrix[30][188] * vector[30] +matrix[31][188] * vector[31] +matrix[32][188] * vector[32] +matrix[33][188] * vector[33] +matrix[34][188] * vector[34] +matrix[35][188] * vector[35] +matrix[36][188] * vector[36] +matrix[37][188] * vector[37] +matrix[38][188] * vector[38] +matrix[39][188] * vector[39] +matrix[40][188] * vector[40] +matrix[41][188] * vector[41] +matrix[42][188] * vector[42] +matrix[43][188] * vector[43] +matrix[44][188] * vector[44] +matrix[45][188] * vector[45] +matrix[46][188] * vector[46] +matrix[47][188] * vector[47] +matrix[48][188] * vector[48] +matrix[49][188] * vector[49] +matrix[50][188] * vector[50] +matrix[51][188] * vector[51] +matrix[52][188] * vector[52] +matrix[53][188] * vector[53] +matrix[54][188] * vector[54] +matrix[55][188] * vector[55] +matrix[56][188] * vector[56] +matrix[57][188] * vector[57] +matrix[58][188] * vector[58] +matrix[59][188] * vector[59] +matrix[60][188] * vector[60] +matrix[61][188] * vector[61] +matrix[62][188] * vector[62] +matrix[63][188] * vector[63] +matrix[64][188] * vector[64] +matrix[65][188] * vector[65] +matrix[66][188] * vector[66] +matrix[67][188] * vector[67] +matrix[68][188] * vector[68] +matrix[69][188] * vector[69] +matrix[70][188] * vector[70] +matrix[71][188] * vector[71] +matrix[72][188] * vector[72] +matrix[73][188] * vector[73] +matrix[74][188] * vector[74] +matrix[75][188] * vector[75] +matrix[76][188] * vector[76] +matrix[77][188] * vector[77] +matrix[78][188] * vector[78] +matrix[79][188] * vector[79] +matrix[80][188] * vector[80] +matrix[81][188] * vector[81] +matrix[82][188] * vector[82] +matrix[83][188] * vector[83] +matrix[84][188] * vector[84] +matrix[85][188] * vector[85] +matrix[86][188] * vector[86] +matrix[87][188] * vector[87] +matrix[88][188] * vector[88] +matrix[89][188] * vector[89] +matrix[90][188] * vector[90] +matrix[91][188] * vector[91] +matrix[92][188] * vector[92] +matrix[93][188] * vector[93] +matrix[94][188] * vector[94] +matrix[95][188] * vector[95] +matrix[96][188] * vector[96] +matrix[97][188] * vector[97] +matrix[98][188] * vector[98] +matrix[99][188] * vector[99] +b[188];
assign result[189] = matrix[0][189] * vector[0] +matrix[1][189] * vector[1] +matrix[2][189] * vector[2] +matrix[3][189] * vector[3] +matrix[4][189] * vector[4] +matrix[5][189] * vector[5] +matrix[6][189] * vector[6] +matrix[7][189] * vector[7] +matrix[8][189] * vector[8] +matrix[9][189] * vector[9] +matrix[10][189] * vector[10] +matrix[11][189] * vector[11] +matrix[12][189] * vector[12] +matrix[13][189] * vector[13] +matrix[14][189] * vector[14] +matrix[15][189] * vector[15] +matrix[16][189] * vector[16] +matrix[17][189] * vector[17] +matrix[18][189] * vector[18] +matrix[19][189] * vector[19] +matrix[20][189] * vector[20] +matrix[21][189] * vector[21] +matrix[22][189] * vector[22] +matrix[23][189] * vector[23] +matrix[24][189] * vector[24] +matrix[25][189] * vector[25] +matrix[26][189] * vector[26] +matrix[27][189] * vector[27] +matrix[28][189] * vector[28] +matrix[29][189] * vector[29] +matrix[30][189] * vector[30] +matrix[31][189] * vector[31] +matrix[32][189] * vector[32] +matrix[33][189] * vector[33] +matrix[34][189] * vector[34] +matrix[35][189] * vector[35] +matrix[36][189] * vector[36] +matrix[37][189] * vector[37] +matrix[38][189] * vector[38] +matrix[39][189] * vector[39] +matrix[40][189] * vector[40] +matrix[41][189] * vector[41] +matrix[42][189] * vector[42] +matrix[43][189] * vector[43] +matrix[44][189] * vector[44] +matrix[45][189] * vector[45] +matrix[46][189] * vector[46] +matrix[47][189] * vector[47] +matrix[48][189] * vector[48] +matrix[49][189] * vector[49] +matrix[50][189] * vector[50] +matrix[51][189] * vector[51] +matrix[52][189] * vector[52] +matrix[53][189] * vector[53] +matrix[54][189] * vector[54] +matrix[55][189] * vector[55] +matrix[56][189] * vector[56] +matrix[57][189] * vector[57] +matrix[58][189] * vector[58] +matrix[59][189] * vector[59] +matrix[60][189] * vector[60] +matrix[61][189] * vector[61] +matrix[62][189] * vector[62] +matrix[63][189] * vector[63] +matrix[64][189] * vector[64] +matrix[65][189] * vector[65] +matrix[66][189] * vector[66] +matrix[67][189] * vector[67] +matrix[68][189] * vector[68] +matrix[69][189] * vector[69] +matrix[70][189] * vector[70] +matrix[71][189] * vector[71] +matrix[72][189] * vector[72] +matrix[73][189] * vector[73] +matrix[74][189] * vector[74] +matrix[75][189] * vector[75] +matrix[76][189] * vector[76] +matrix[77][189] * vector[77] +matrix[78][189] * vector[78] +matrix[79][189] * vector[79] +matrix[80][189] * vector[80] +matrix[81][189] * vector[81] +matrix[82][189] * vector[82] +matrix[83][189] * vector[83] +matrix[84][189] * vector[84] +matrix[85][189] * vector[85] +matrix[86][189] * vector[86] +matrix[87][189] * vector[87] +matrix[88][189] * vector[88] +matrix[89][189] * vector[89] +matrix[90][189] * vector[90] +matrix[91][189] * vector[91] +matrix[92][189] * vector[92] +matrix[93][189] * vector[93] +matrix[94][189] * vector[94] +matrix[95][189] * vector[95] +matrix[96][189] * vector[96] +matrix[97][189] * vector[97] +matrix[98][189] * vector[98] +matrix[99][189] * vector[99] +b[189];
assign result[190] = matrix[0][190] * vector[0] +matrix[1][190] * vector[1] +matrix[2][190] * vector[2] +matrix[3][190] * vector[3] +matrix[4][190] * vector[4] +matrix[5][190] * vector[5] +matrix[6][190] * vector[6] +matrix[7][190] * vector[7] +matrix[8][190] * vector[8] +matrix[9][190] * vector[9] +matrix[10][190] * vector[10] +matrix[11][190] * vector[11] +matrix[12][190] * vector[12] +matrix[13][190] * vector[13] +matrix[14][190] * vector[14] +matrix[15][190] * vector[15] +matrix[16][190] * vector[16] +matrix[17][190] * vector[17] +matrix[18][190] * vector[18] +matrix[19][190] * vector[19] +matrix[20][190] * vector[20] +matrix[21][190] * vector[21] +matrix[22][190] * vector[22] +matrix[23][190] * vector[23] +matrix[24][190] * vector[24] +matrix[25][190] * vector[25] +matrix[26][190] * vector[26] +matrix[27][190] * vector[27] +matrix[28][190] * vector[28] +matrix[29][190] * vector[29] +matrix[30][190] * vector[30] +matrix[31][190] * vector[31] +matrix[32][190] * vector[32] +matrix[33][190] * vector[33] +matrix[34][190] * vector[34] +matrix[35][190] * vector[35] +matrix[36][190] * vector[36] +matrix[37][190] * vector[37] +matrix[38][190] * vector[38] +matrix[39][190] * vector[39] +matrix[40][190] * vector[40] +matrix[41][190] * vector[41] +matrix[42][190] * vector[42] +matrix[43][190] * vector[43] +matrix[44][190] * vector[44] +matrix[45][190] * vector[45] +matrix[46][190] * vector[46] +matrix[47][190] * vector[47] +matrix[48][190] * vector[48] +matrix[49][190] * vector[49] +matrix[50][190] * vector[50] +matrix[51][190] * vector[51] +matrix[52][190] * vector[52] +matrix[53][190] * vector[53] +matrix[54][190] * vector[54] +matrix[55][190] * vector[55] +matrix[56][190] * vector[56] +matrix[57][190] * vector[57] +matrix[58][190] * vector[58] +matrix[59][190] * vector[59] +matrix[60][190] * vector[60] +matrix[61][190] * vector[61] +matrix[62][190] * vector[62] +matrix[63][190] * vector[63] +matrix[64][190] * vector[64] +matrix[65][190] * vector[65] +matrix[66][190] * vector[66] +matrix[67][190] * vector[67] +matrix[68][190] * vector[68] +matrix[69][190] * vector[69] +matrix[70][190] * vector[70] +matrix[71][190] * vector[71] +matrix[72][190] * vector[72] +matrix[73][190] * vector[73] +matrix[74][190] * vector[74] +matrix[75][190] * vector[75] +matrix[76][190] * vector[76] +matrix[77][190] * vector[77] +matrix[78][190] * vector[78] +matrix[79][190] * vector[79] +matrix[80][190] * vector[80] +matrix[81][190] * vector[81] +matrix[82][190] * vector[82] +matrix[83][190] * vector[83] +matrix[84][190] * vector[84] +matrix[85][190] * vector[85] +matrix[86][190] * vector[86] +matrix[87][190] * vector[87] +matrix[88][190] * vector[88] +matrix[89][190] * vector[89] +matrix[90][190] * vector[90] +matrix[91][190] * vector[91] +matrix[92][190] * vector[92] +matrix[93][190] * vector[93] +matrix[94][190] * vector[94] +matrix[95][190] * vector[95] +matrix[96][190] * vector[96] +matrix[97][190] * vector[97] +matrix[98][190] * vector[98] +matrix[99][190] * vector[99] +b[190];
assign result[191] = matrix[0][191] * vector[0] +matrix[1][191] * vector[1] +matrix[2][191] * vector[2] +matrix[3][191] * vector[3] +matrix[4][191] * vector[4] +matrix[5][191] * vector[5] +matrix[6][191] * vector[6] +matrix[7][191] * vector[7] +matrix[8][191] * vector[8] +matrix[9][191] * vector[9] +matrix[10][191] * vector[10] +matrix[11][191] * vector[11] +matrix[12][191] * vector[12] +matrix[13][191] * vector[13] +matrix[14][191] * vector[14] +matrix[15][191] * vector[15] +matrix[16][191] * vector[16] +matrix[17][191] * vector[17] +matrix[18][191] * vector[18] +matrix[19][191] * vector[19] +matrix[20][191] * vector[20] +matrix[21][191] * vector[21] +matrix[22][191] * vector[22] +matrix[23][191] * vector[23] +matrix[24][191] * vector[24] +matrix[25][191] * vector[25] +matrix[26][191] * vector[26] +matrix[27][191] * vector[27] +matrix[28][191] * vector[28] +matrix[29][191] * vector[29] +matrix[30][191] * vector[30] +matrix[31][191] * vector[31] +matrix[32][191] * vector[32] +matrix[33][191] * vector[33] +matrix[34][191] * vector[34] +matrix[35][191] * vector[35] +matrix[36][191] * vector[36] +matrix[37][191] * vector[37] +matrix[38][191] * vector[38] +matrix[39][191] * vector[39] +matrix[40][191] * vector[40] +matrix[41][191] * vector[41] +matrix[42][191] * vector[42] +matrix[43][191] * vector[43] +matrix[44][191] * vector[44] +matrix[45][191] * vector[45] +matrix[46][191] * vector[46] +matrix[47][191] * vector[47] +matrix[48][191] * vector[48] +matrix[49][191] * vector[49] +matrix[50][191] * vector[50] +matrix[51][191] * vector[51] +matrix[52][191] * vector[52] +matrix[53][191] * vector[53] +matrix[54][191] * vector[54] +matrix[55][191] * vector[55] +matrix[56][191] * vector[56] +matrix[57][191] * vector[57] +matrix[58][191] * vector[58] +matrix[59][191] * vector[59] +matrix[60][191] * vector[60] +matrix[61][191] * vector[61] +matrix[62][191] * vector[62] +matrix[63][191] * vector[63] +matrix[64][191] * vector[64] +matrix[65][191] * vector[65] +matrix[66][191] * vector[66] +matrix[67][191] * vector[67] +matrix[68][191] * vector[68] +matrix[69][191] * vector[69] +matrix[70][191] * vector[70] +matrix[71][191] * vector[71] +matrix[72][191] * vector[72] +matrix[73][191] * vector[73] +matrix[74][191] * vector[74] +matrix[75][191] * vector[75] +matrix[76][191] * vector[76] +matrix[77][191] * vector[77] +matrix[78][191] * vector[78] +matrix[79][191] * vector[79] +matrix[80][191] * vector[80] +matrix[81][191] * vector[81] +matrix[82][191] * vector[82] +matrix[83][191] * vector[83] +matrix[84][191] * vector[84] +matrix[85][191] * vector[85] +matrix[86][191] * vector[86] +matrix[87][191] * vector[87] +matrix[88][191] * vector[88] +matrix[89][191] * vector[89] +matrix[90][191] * vector[90] +matrix[91][191] * vector[91] +matrix[92][191] * vector[92] +matrix[93][191] * vector[93] +matrix[94][191] * vector[94] +matrix[95][191] * vector[95] +matrix[96][191] * vector[96] +matrix[97][191] * vector[97] +matrix[98][191] * vector[98] +matrix[99][191] * vector[99] +b[191];
assign result[192] = matrix[0][192] * vector[0] +matrix[1][192] * vector[1] +matrix[2][192] * vector[2] +matrix[3][192] * vector[3] +matrix[4][192] * vector[4] +matrix[5][192] * vector[5] +matrix[6][192] * vector[6] +matrix[7][192] * vector[7] +matrix[8][192] * vector[8] +matrix[9][192] * vector[9] +matrix[10][192] * vector[10] +matrix[11][192] * vector[11] +matrix[12][192] * vector[12] +matrix[13][192] * vector[13] +matrix[14][192] * vector[14] +matrix[15][192] * vector[15] +matrix[16][192] * vector[16] +matrix[17][192] * vector[17] +matrix[18][192] * vector[18] +matrix[19][192] * vector[19] +matrix[20][192] * vector[20] +matrix[21][192] * vector[21] +matrix[22][192] * vector[22] +matrix[23][192] * vector[23] +matrix[24][192] * vector[24] +matrix[25][192] * vector[25] +matrix[26][192] * vector[26] +matrix[27][192] * vector[27] +matrix[28][192] * vector[28] +matrix[29][192] * vector[29] +matrix[30][192] * vector[30] +matrix[31][192] * vector[31] +matrix[32][192] * vector[32] +matrix[33][192] * vector[33] +matrix[34][192] * vector[34] +matrix[35][192] * vector[35] +matrix[36][192] * vector[36] +matrix[37][192] * vector[37] +matrix[38][192] * vector[38] +matrix[39][192] * vector[39] +matrix[40][192] * vector[40] +matrix[41][192] * vector[41] +matrix[42][192] * vector[42] +matrix[43][192] * vector[43] +matrix[44][192] * vector[44] +matrix[45][192] * vector[45] +matrix[46][192] * vector[46] +matrix[47][192] * vector[47] +matrix[48][192] * vector[48] +matrix[49][192] * vector[49] +matrix[50][192] * vector[50] +matrix[51][192] * vector[51] +matrix[52][192] * vector[52] +matrix[53][192] * vector[53] +matrix[54][192] * vector[54] +matrix[55][192] * vector[55] +matrix[56][192] * vector[56] +matrix[57][192] * vector[57] +matrix[58][192] * vector[58] +matrix[59][192] * vector[59] +matrix[60][192] * vector[60] +matrix[61][192] * vector[61] +matrix[62][192] * vector[62] +matrix[63][192] * vector[63] +matrix[64][192] * vector[64] +matrix[65][192] * vector[65] +matrix[66][192] * vector[66] +matrix[67][192] * vector[67] +matrix[68][192] * vector[68] +matrix[69][192] * vector[69] +matrix[70][192] * vector[70] +matrix[71][192] * vector[71] +matrix[72][192] * vector[72] +matrix[73][192] * vector[73] +matrix[74][192] * vector[74] +matrix[75][192] * vector[75] +matrix[76][192] * vector[76] +matrix[77][192] * vector[77] +matrix[78][192] * vector[78] +matrix[79][192] * vector[79] +matrix[80][192] * vector[80] +matrix[81][192] * vector[81] +matrix[82][192] * vector[82] +matrix[83][192] * vector[83] +matrix[84][192] * vector[84] +matrix[85][192] * vector[85] +matrix[86][192] * vector[86] +matrix[87][192] * vector[87] +matrix[88][192] * vector[88] +matrix[89][192] * vector[89] +matrix[90][192] * vector[90] +matrix[91][192] * vector[91] +matrix[92][192] * vector[92] +matrix[93][192] * vector[93] +matrix[94][192] * vector[94] +matrix[95][192] * vector[95] +matrix[96][192] * vector[96] +matrix[97][192] * vector[97] +matrix[98][192] * vector[98] +matrix[99][192] * vector[99] +b[192];
assign result[193] = matrix[0][193] * vector[0] +matrix[1][193] * vector[1] +matrix[2][193] * vector[2] +matrix[3][193] * vector[3] +matrix[4][193] * vector[4] +matrix[5][193] * vector[5] +matrix[6][193] * vector[6] +matrix[7][193] * vector[7] +matrix[8][193] * vector[8] +matrix[9][193] * vector[9] +matrix[10][193] * vector[10] +matrix[11][193] * vector[11] +matrix[12][193] * vector[12] +matrix[13][193] * vector[13] +matrix[14][193] * vector[14] +matrix[15][193] * vector[15] +matrix[16][193] * vector[16] +matrix[17][193] * vector[17] +matrix[18][193] * vector[18] +matrix[19][193] * vector[19] +matrix[20][193] * vector[20] +matrix[21][193] * vector[21] +matrix[22][193] * vector[22] +matrix[23][193] * vector[23] +matrix[24][193] * vector[24] +matrix[25][193] * vector[25] +matrix[26][193] * vector[26] +matrix[27][193] * vector[27] +matrix[28][193] * vector[28] +matrix[29][193] * vector[29] +matrix[30][193] * vector[30] +matrix[31][193] * vector[31] +matrix[32][193] * vector[32] +matrix[33][193] * vector[33] +matrix[34][193] * vector[34] +matrix[35][193] * vector[35] +matrix[36][193] * vector[36] +matrix[37][193] * vector[37] +matrix[38][193] * vector[38] +matrix[39][193] * vector[39] +matrix[40][193] * vector[40] +matrix[41][193] * vector[41] +matrix[42][193] * vector[42] +matrix[43][193] * vector[43] +matrix[44][193] * vector[44] +matrix[45][193] * vector[45] +matrix[46][193] * vector[46] +matrix[47][193] * vector[47] +matrix[48][193] * vector[48] +matrix[49][193] * vector[49] +matrix[50][193] * vector[50] +matrix[51][193] * vector[51] +matrix[52][193] * vector[52] +matrix[53][193] * vector[53] +matrix[54][193] * vector[54] +matrix[55][193] * vector[55] +matrix[56][193] * vector[56] +matrix[57][193] * vector[57] +matrix[58][193] * vector[58] +matrix[59][193] * vector[59] +matrix[60][193] * vector[60] +matrix[61][193] * vector[61] +matrix[62][193] * vector[62] +matrix[63][193] * vector[63] +matrix[64][193] * vector[64] +matrix[65][193] * vector[65] +matrix[66][193] * vector[66] +matrix[67][193] * vector[67] +matrix[68][193] * vector[68] +matrix[69][193] * vector[69] +matrix[70][193] * vector[70] +matrix[71][193] * vector[71] +matrix[72][193] * vector[72] +matrix[73][193] * vector[73] +matrix[74][193] * vector[74] +matrix[75][193] * vector[75] +matrix[76][193] * vector[76] +matrix[77][193] * vector[77] +matrix[78][193] * vector[78] +matrix[79][193] * vector[79] +matrix[80][193] * vector[80] +matrix[81][193] * vector[81] +matrix[82][193] * vector[82] +matrix[83][193] * vector[83] +matrix[84][193] * vector[84] +matrix[85][193] * vector[85] +matrix[86][193] * vector[86] +matrix[87][193] * vector[87] +matrix[88][193] * vector[88] +matrix[89][193] * vector[89] +matrix[90][193] * vector[90] +matrix[91][193] * vector[91] +matrix[92][193] * vector[92] +matrix[93][193] * vector[93] +matrix[94][193] * vector[94] +matrix[95][193] * vector[95] +matrix[96][193] * vector[96] +matrix[97][193] * vector[97] +matrix[98][193] * vector[98] +matrix[99][193] * vector[99] +b[193];
assign result[194] = matrix[0][194] * vector[0] +matrix[1][194] * vector[1] +matrix[2][194] * vector[2] +matrix[3][194] * vector[3] +matrix[4][194] * vector[4] +matrix[5][194] * vector[5] +matrix[6][194] * vector[6] +matrix[7][194] * vector[7] +matrix[8][194] * vector[8] +matrix[9][194] * vector[9] +matrix[10][194] * vector[10] +matrix[11][194] * vector[11] +matrix[12][194] * vector[12] +matrix[13][194] * vector[13] +matrix[14][194] * vector[14] +matrix[15][194] * vector[15] +matrix[16][194] * vector[16] +matrix[17][194] * vector[17] +matrix[18][194] * vector[18] +matrix[19][194] * vector[19] +matrix[20][194] * vector[20] +matrix[21][194] * vector[21] +matrix[22][194] * vector[22] +matrix[23][194] * vector[23] +matrix[24][194] * vector[24] +matrix[25][194] * vector[25] +matrix[26][194] * vector[26] +matrix[27][194] * vector[27] +matrix[28][194] * vector[28] +matrix[29][194] * vector[29] +matrix[30][194] * vector[30] +matrix[31][194] * vector[31] +matrix[32][194] * vector[32] +matrix[33][194] * vector[33] +matrix[34][194] * vector[34] +matrix[35][194] * vector[35] +matrix[36][194] * vector[36] +matrix[37][194] * vector[37] +matrix[38][194] * vector[38] +matrix[39][194] * vector[39] +matrix[40][194] * vector[40] +matrix[41][194] * vector[41] +matrix[42][194] * vector[42] +matrix[43][194] * vector[43] +matrix[44][194] * vector[44] +matrix[45][194] * vector[45] +matrix[46][194] * vector[46] +matrix[47][194] * vector[47] +matrix[48][194] * vector[48] +matrix[49][194] * vector[49] +matrix[50][194] * vector[50] +matrix[51][194] * vector[51] +matrix[52][194] * vector[52] +matrix[53][194] * vector[53] +matrix[54][194] * vector[54] +matrix[55][194] * vector[55] +matrix[56][194] * vector[56] +matrix[57][194] * vector[57] +matrix[58][194] * vector[58] +matrix[59][194] * vector[59] +matrix[60][194] * vector[60] +matrix[61][194] * vector[61] +matrix[62][194] * vector[62] +matrix[63][194] * vector[63] +matrix[64][194] * vector[64] +matrix[65][194] * vector[65] +matrix[66][194] * vector[66] +matrix[67][194] * vector[67] +matrix[68][194] * vector[68] +matrix[69][194] * vector[69] +matrix[70][194] * vector[70] +matrix[71][194] * vector[71] +matrix[72][194] * vector[72] +matrix[73][194] * vector[73] +matrix[74][194] * vector[74] +matrix[75][194] * vector[75] +matrix[76][194] * vector[76] +matrix[77][194] * vector[77] +matrix[78][194] * vector[78] +matrix[79][194] * vector[79] +matrix[80][194] * vector[80] +matrix[81][194] * vector[81] +matrix[82][194] * vector[82] +matrix[83][194] * vector[83] +matrix[84][194] * vector[84] +matrix[85][194] * vector[85] +matrix[86][194] * vector[86] +matrix[87][194] * vector[87] +matrix[88][194] * vector[88] +matrix[89][194] * vector[89] +matrix[90][194] * vector[90] +matrix[91][194] * vector[91] +matrix[92][194] * vector[92] +matrix[93][194] * vector[93] +matrix[94][194] * vector[94] +matrix[95][194] * vector[95] +matrix[96][194] * vector[96] +matrix[97][194] * vector[97] +matrix[98][194] * vector[98] +matrix[99][194] * vector[99] +b[194];
assign result[195] = matrix[0][195] * vector[0] +matrix[1][195] * vector[1] +matrix[2][195] * vector[2] +matrix[3][195] * vector[3] +matrix[4][195] * vector[4] +matrix[5][195] * vector[5] +matrix[6][195] * vector[6] +matrix[7][195] * vector[7] +matrix[8][195] * vector[8] +matrix[9][195] * vector[9] +matrix[10][195] * vector[10] +matrix[11][195] * vector[11] +matrix[12][195] * vector[12] +matrix[13][195] * vector[13] +matrix[14][195] * vector[14] +matrix[15][195] * vector[15] +matrix[16][195] * vector[16] +matrix[17][195] * vector[17] +matrix[18][195] * vector[18] +matrix[19][195] * vector[19] +matrix[20][195] * vector[20] +matrix[21][195] * vector[21] +matrix[22][195] * vector[22] +matrix[23][195] * vector[23] +matrix[24][195] * vector[24] +matrix[25][195] * vector[25] +matrix[26][195] * vector[26] +matrix[27][195] * vector[27] +matrix[28][195] * vector[28] +matrix[29][195] * vector[29] +matrix[30][195] * vector[30] +matrix[31][195] * vector[31] +matrix[32][195] * vector[32] +matrix[33][195] * vector[33] +matrix[34][195] * vector[34] +matrix[35][195] * vector[35] +matrix[36][195] * vector[36] +matrix[37][195] * vector[37] +matrix[38][195] * vector[38] +matrix[39][195] * vector[39] +matrix[40][195] * vector[40] +matrix[41][195] * vector[41] +matrix[42][195] * vector[42] +matrix[43][195] * vector[43] +matrix[44][195] * vector[44] +matrix[45][195] * vector[45] +matrix[46][195] * vector[46] +matrix[47][195] * vector[47] +matrix[48][195] * vector[48] +matrix[49][195] * vector[49] +matrix[50][195] * vector[50] +matrix[51][195] * vector[51] +matrix[52][195] * vector[52] +matrix[53][195] * vector[53] +matrix[54][195] * vector[54] +matrix[55][195] * vector[55] +matrix[56][195] * vector[56] +matrix[57][195] * vector[57] +matrix[58][195] * vector[58] +matrix[59][195] * vector[59] +matrix[60][195] * vector[60] +matrix[61][195] * vector[61] +matrix[62][195] * vector[62] +matrix[63][195] * vector[63] +matrix[64][195] * vector[64] +matrix[65][195] * vector[65] +matrix[66][195] * vector[66] +matrix[67][195] * vector[67] +matrix[68][195] * vector[68] +matrix[69][195] * vector[69] +matrix[70][195] * vector[70] +matrix[71][195] * vector[71] +matrix[72][195] * vector[72] +matrix[73][195] * vector[73] +matrix[74][195] * vector[74] +matrix[75][195] * vector[75] +matrix[76][195] * vector[76] +matrix[77][195] * vector[77] +matrix[78][195] * vector[78] +matrix[79][195] * vector[79] +matrix[80][195] * vector[80] +matrix[81][195] * vector[81] +matrix[82][195] * vector[82] +matrix[83][195] * vector[83] +matrix[84][195] * vector[84] +matrix[85][195] * vector[85] +matrix[86][195] * vector[86] +matrix[87][195] * vector[87] +matrix[88][195] * vector[88] +matrix[89][195] * vector[89] +matrix[90][195] * vector[90] +matrix[91][195] * vector[91] +matrix[92][195] * vector[92] +matrix[93][195] * vector[93] +matrix[94][195] * vector[94] +matrix[95][195] * vector[95] +matrix[96][195] * vector[96] +matrix[97][195] * vector[97] +matrix[98][195] * vector[98] +matrix[99][195] * vector[99] +b[195];
assign result[196] = matrix[0][196] * vector[0] +matrix[1][196] * vector[1] +matrix[2][196] * vector[2] +matrix[3][196] * vector[3] +matrix[4][196] * vector[4] +matrix[5][196] * vector[5] +matrix[6][196] * vector[6] +matrix[7][196] * vector[7] +matrix[8][196] * vector[8] +matrix[9][196] * vector[9] +matrix[10][196] * vector[10] +matrix[11][196] * vector[11] +matrix[12][196] * vector[12] +matrix[13][196] * vector[13] +matrix[14][196] * vector[14] +matrix[15][196] * vector[15] +matrix[16][196] * vector[16] +matrix[17][196] * vector[17] +matrix[18][196] * vector[18] +matrix[19][196] * vector[19] +matrix[20][196] * vector[20] +matrix[21][196] * vector[21] +matrix[22][196] * vector[22] +matrix[23][196] * vector[23] +matrix[24][196] * vector[24] +matrix[25][196] * vector[25] +matrix[26][196] * vector[26] +matrix[27][196] * vector[27] +matrix[28][196] * vector[28] +matrix[29][196] * vector[29] +matrix[30][196] * vector[30] +matrix[31][196] * vector[31] +matrix[32][196] * vector[32] +matrix[33][196] * vector[33] +matrix[34][196] * vector[34] +matrix[35][196] * vector[35] +matrix[36][196] * vector[36] +matrix[37][196] * vector[37] +matrix[38][196] * vector[38] +matrix[39][196] * vector[39] +matrix[40][196] * vector[40] +matrix[41][196] * vector[41] +matrix[42][196] * vector[42] +matrix[43][196] * vector[43] +matrix[44][196] * vector[44] +matrix[45][196] * vector[45] +matrix[46][196] * vector[46] +matrix[47][196] * vector[47] +matrix[48][196] * vector[48] +matrix[49][196] * vector[49] +matrix[50][196] * vector[50] +matrix[51][196] * vector[51] +matrix[52][196] * vector[52] +matrix[53][196] * vector[53] +matrix[54][196] * vector[54] +matrix[55][196] * vector[55] +matrix[56][196] * vector[56] +matrix[57][196] * vector[57] +matrix[58][196] * vector[58] +matrix[59][196] * vector[59] +matrix[60][196] * vector[60] +matrix[61][196] * vector[61] +matrix[62][196] * vector[62] +matrix[63][196] * vector[63] +matrix[64][196] * vector[64] +matrix[65][196] * vector[65] +matrix[66][196] * vector[66] +matrix[67][196] * vector[67] +matrix[68][196] * vector[68] +matrix[69][196] * vector[69] +matrix[70][196] * vector[70] +matrix[71][196] * vector[71] +matrix[72][196] * vector[72] +matrix[73][196] * vector[73] +matrix[74][196] * vector[74] +matrix[75][196] * vector[75] +matrix[76][196] * vector[76] +matrix[77][196] * vector[77] +matrix[78][196] * vector[78] +matrix[79][196] * vector[79] +matrix[80][196] * vector[80] +matrix[81][196] * vector[81] +matrix[82][196] * vector[82] +matrix[83][196] * vector[83] +matrix[84][196] * vector[84] +matrix[85][196] * vector[85] +matrix[86][196] * vector[86] +matrix[87][196] * vector[87] +matrix[88][196] * vector[88] +matrix[89][196] * vector[89] +matrix[90][196] * vector[90] +matrix[91][196] * vector[91] +matrix[92][196] * vector[92] +matrix[93][196] * vector[93] +matrix[94][196] * vector[94] +matrix[95][196] * vector[95] +matrix[96][196] * vector[96] +matrix[97][196] * vector[97] +matrix[98][196] * vector[98] +matrix[99][196] * vector[99] +b[196];
assign result[197] = matrix[0][197] * vector[0] +matrix[1][197] * vector[1] +matrix[2][197] * vector[2] +matrix[3][197] * vector[3] +matrix[4][197] * vector[4] +matrix[5][197] * vector[5] +matrix[6][197] * vector[6] +matrix[7][197] * vector[7] +matrix[8][197] * vector[8] +matrix[9][197] * vector[9] +matrix[10][197] * vector[10] +matrix[11][197] * vector[11] +matrix[12][197] * vector[12] +matrix[13][197] * vector[13] +matrix[14][197] * vector[14] +matrix[15][197] * vector[15] +matrix[16][197] * vector[16] +matrix[17][197] * vector[17] +matrix[18][197] * vector[18] +matrix[19][197] * vector[19] +matrix[20][197] * vector[20] +matrix[21][197] * vector[21] +matrix[22][197] * vector[22] +matrix[23][197] * vector[23] +matrix[24][197] * vector[24] +matrix[25][197] * vector[25] +matrix[26][197] * vector[26] +matrix[27][197] * vector[27] +matrix[28][197] * vector[28] +matrix[29][197] * vector[29] +matrix[30][197] * vector[30] +matrix[31][197] * vector[31] +matrix[32][197] * vector[32] +matrix[33][197] * vector[33] +matrix[34][197] * vector[34] +matrix[35][197] * vector[35] +matrix[36][197] * vector[36] +matrix[37][197] * vector[37] +matrix[38][197] * vector[38] +matrix[39][197] * vector[39] +matrix[40][197] * vector[40] +matrix[41][197] * vector[41] +matrix[42][197] * vector[42] +matrix[43][197] * vector[43] +matrix[44][197] * vector[44] +matrix[45][197] * vector[45] +matrix[46][197] * vector[46] +matrix[47][197] * vector[47] +matrix[48][197] * vector[48] +matrix[49][197] * vector[49] +matrix[50][197] * vector[50] +matrix[51][197] * vector[51] +matrix[52][197] * vector[52] +matrix[53][197] * vector[53] +matrix[54][197] * vector[54] +matrix[55][197] * vector[55] +matrix[56][197] * vector[56] +matrix[57][197] * vector[57] +matrix[58][197] * vector[58] +matrix[59][197] * vector[59] +matrix[60][197] * vector[60] +matrix[61][197] * vector[61] +matrix[62][197] * vector[62] +matrix[63][197] * vector[63] +matrix[64][197] * vector[64] +matrix[65][197] * vector[65] +matrix[66][197] * vector[66] +matrix[67][197] * vector[67] +matrix[68][197] * vector[68] +matrix[69][197] * vector[69] +matrix[70][197] * vector[70] +matrix[71][197] * vector[71] +matrix[72][197] * vector[72] +matrix[73][197] * vector[73] +matrix[74][197] * vector[74] +matrix[75][197] * vector[75] +matrix[76][197] * vector[76] +matrix[77][197] * vector[77] +matrix[78][197] * vector[78] +matrix[79][197] * vector[79] +matrix[80][197] * vector[80] +matrix[81][197] * vector[81] +matrix[82][197] * vector[82] +matrix[83][197] * vector[83] +matrix[84][197] * vector[84] +matrix[85][197] * vector[85] +matrix[86][197] * vector[86] +matrix[87][197] * vector[87] +matrix[88][197] * vector[88] +matrix[89][197] * vector[89] +matrix[90][197] * vector[90] +matrix[91][197] * vector[91] +matrix[92][197] * vector[92] +matrix[93][197] * vector[93] +matrix[94][197] * vector[94] +matrix[95][197] * vector[95] +matrix[96][197] * vector[96] +matrix[97][197] * vector[97] +matrix[98][197] * vector[98] +matrix[99][197] * vector[99] +b[197];
assign result[198] = matrix[0][198] * vector[0] +matrix[1][198] * vector[1] +matrix[2][198] * vector[2] +matrix[3][198] * vector[3] +matrix[4][198] * vector[4] +matrix[5][198] * vector[5] +matrix[6][198] * vector[6] +matrix[7][198] * vector[7] +matrix[8][198] * vector[8] +matrix[9][198] * vector[9] +matrix[10][198] * vector[10] +matrix[11][198] * vector[11] +matrix[12][198] * vector[12] +matrix[13][198] * vector[13] +matrix[14][198] * vector[14] +matrix[15][198] * vector[15] +matrix[16][198] * vector[16] +matrix[17][198] * vector[17] +matrix[18][198] * vector[18] +matrix[19][198] * vector[19] +matrix[20][198] * vector[20] +matrix[21][198] * vector[21] +matrix[22][198] * vector[22] +matrix[23][198] * vector[23] +matrix[24][198] * vector[24] +matrix[25][198] * vector[25] +matrix[26][198] * vector[26] +matrix[27][198] * vector[27] +matrix[28][198] * vector[28] +matrix[29][198] * vector[29] +matrix[30][198] * vector[30] +matrix[31][198] * vector[31] +matrix[32][198] * vector[32] +matrix[33][198] * vector[33] +matrix[34][198] * vector[34] +matrix[35][198] * vector[35] +matrix[36][198] * vector[36] +matrix[37][198] * vector[37] +matrix[38][198] * vector[38] +matrix[39][198] * vector[39] +matrix[40][198] * vector[40] +matrix[41][198] * vector[41] +matrix[42][198] * vector[42] +matrix[43][198] * vector[43] +matrix[44][198] * vector[44] +matrix[45][198] * vector[45] +matrix[46][198] * vector[46] +matrix[47][198] * vector[47] +matrix[48][198] * vector[48] +matrix[49][198] * vector[49] +matrix[50][198] * vector[50] +matrix[51][198] * vector[51] +matrix[52][198] * vector[52] +matrix[53][198] * vector[53] +matrix[54][198] * vector[54] +matrix[55][198] * vector[55] +matrix[56][198] * vector[56] +matrix[57][198] * vector[57] +matrix[58][198] * vector[58] +matrix[59][198] * vector[59] +matrix[60][198] * vector[60] +matrix[61][198] * vector[61] +matrix[62][198] * vector[62] +matrix[63][198] * vector[63] +matrix[64][198] * vector[64] +matrix[65][198] * vector[65] +matrix[66][198] * vector[66] +matrix[67][198] * vector[67] +matrix[68][198] * vector[68] +matrix[69][198] * vector[69] +matrix[70][198] * vector[70] +matrix[71][198] * vector[71] +matrix[72][198] * vector[72] +matrix[73][198] * vector[73] +matrix[74][198] * vector[74] +matrix[75][198] * vector[75] +matrix[76][198] * vector[76] +matrix[77][198] * vector[77] +matrix[78][198] * vector[78] +matrix[79][198] * vector[79] +matrix[80][198] * vector[80] +matrix[81][198] * vector[81] +matrix[82][198] * vector[82] +matrix[83][198] * vector[83] +matrix[84][198] * vector[84] +matrix[85][198] * vector[85] +matrix[86][198] * vector[86] +matrix[87][198] * vector[87] +matrix[88][198] * vector[88] +matrix[89][198] * vector[89] +matrix[90][198] * vector[90] +matrix[91][198] * vector[91] +matrix[92][198] * vector[92] +matrix[93][198] * vector[93] +matrix[94][198] * vector[94] +matrix[95][198] * vector[95] +matrix[96][198] * vector[96] +matrix[97][198] * vector[97] +matrix[98][198] * vector[98] +matrix[99][198] * vector[99] +b[198];
assign result[199] = matrix[0][199] * vector[0] +matrix[1][199] * vector[1] +matrix[2][199] * vector[2] +matrix[3][199] * vector[3] +matrix[4][199] * vector[4] +matrix[5][199] * vector[5] +matrix[6][199] * vector[6] +matrix[7][199] * vector[7] +matrix[8][199] * vector[8] +matrix[9][199] * vector[9] +matrix[10][199] * vector[10] +matrix[11][199] * vector[11] +matrix[12][199] * vector[12] +matrix[13][199] * vector[13] +matrix[14][199] * vector[14] +matrix[15][199] * vector[15] +matrix[16][199] * vector[16] +matrix[17][199] * vector[17] +matrix[18][199] * vector[18] +matrix[19][199] * vector[19] +matrix[20][199] * vector[20] +matrix[21][199] * vector[21] +matrix[22][199] * vector[22] +matrix[23][199] * vector[23] +matrix[24][199] * vector[24] +matrix[25][199] * vector[25] +matrix[26][199] * vector[26] +matrix[27][199] * vector[27] +matrix[28][199] * vector[28] +matrix[29][199] * vector[29] +matrix[30][199] * vector[30] +matrix[31][199] * vector[31] +matrix[32][199] * vector[32] +matrix[33][199] * vector[33] +matrix[34][199] * vector[34] +matrix[35][199] * vector[35] +matrix[36][199] * vector[36] +matrix[37][199] * vector[37] +matrix[38][199] * vector[38] +matrix[39][199] * vector[39] +matrix[40][199] * vector[40] +matrix[41][199] * vector[41] +matrix[42][199] * vector[42] +matrix[43][199] * vector[43] +matrix[44][199] * vector[44] +matrix[45][199] * vector[45] +matrix[46][199] * vector[46] +matrix[47][199] * vector[47] +matrix[48][199] * vector[48] +matrix[49][199] * vector[49] +matrix[50][199] * vector[50] +matrix[51][199] * vector[51] +matrix[52][199] * vector[52] +matrix[53][199] * vector[53] +matrix[54][199] * vector[54] +matrix[55][199] * vector[55] +matrix[56][199] * vector[56] +matrix[57][199] * vector[57] +matrix[58][199] * vector[58] +matrix[59][199] * vector[59] +matrix[60][199] * vector[60] +matrix[61][199] * vector[61] +matrix[62][199] * vector[62] +matrix[63][199] * vector[63] +matrix[64][199] * vector[64] +matrix[65][199] * vector[65] +matrix[66][199] * vector[66] +matrix[67][199] * vector[67] +matrix[68][199] * vector[68] +matrix[69][199] * vector[69] +matrix[70][199] * vector[70] +matrix[71][199] * vector[71] +matrix[72][199] * vector[72] +matrix[73][199] * vector[73] +matrix[74][199] * vector[74] +matrix[75][199] * vector[75] +matrix[76][199] * vector[76] +matrix[77][199] * vector[77] +matrix[78][199] * vector[78] +matrix[79][199] * vector[79] +matrix[80][199] * vector[80] +matrix[81][199] * vector[81] +matrix[82][199] * vector[82] +matrix[83][199] * vector[83] +matrix[84][199] * vector[84] +matrix[85][199] * vector[85] +matrix[86][199] * vector[86] +matrix[87][199] * vector[87] +matrix[88][199] * vector[88] +matrix[89][199] * vector[89] +matrix[90][199] * vector[90] +matrix[91][199] * vector[91] +matrix[92][199] * vector[92] +matrix[93][199] * vector[93] +matrix[94][199] * vector[94] +matrix[95][199] * vector[95] +matrix[96][199] * vector[96] +matrix[97][199] * vector[97] +matrix[98][199] * vector[98] +matrix[99][199] * vector[99] +b[199];
assign result[200] = matrix[0][200] * vector[0] +matrix[1][200] * vector[1] +matrix[2][200] * vector[2] +matrix[3][200] * vector[3] +matrix[4][200] * vector[4] +matrix[5][200] * vector[5] +matrix[6][200] * vector[6] +matrix[7][200] * vector[7] +matrix[8][200] * vector[8] +matrix[9][200] * vector[9] +matrix[10][200] * vector[10] +matrix[11][200] * vector[11] +matrix[12][200] * vector[12] +matrix[13][200] * vector[13] +matrix[14][200] * vector[14] +matrix[15][200] * vector[15] +matrix[16][200] * vector[16] +matrix[17][200] * vector[17] +matrix[18][200] * vector[18] +matrix[19][200] * vector[19] +matrix[20][200] * vector[20] +matrix[21][200] * vector[21] +matrix[22][200] * vector[22] +matrix[23][200] * vector[23] +matrix[24][200] * vector[24] +matrix[25][200] * vector[25] +matrix[26][200] * vector[26] +matrix[27][200] * vector[27] +matrix[28][200] * vector[28] +matrix[29][200] * vector[29] +matrix[30][200] * vector[30] +matrix[31][200] * vector[31] +matrix[32][200] * vector[32] +matrix[33][200] * vector[33] +matrix[34][200] * vector[34] +matrix[35][200] * vector[35] +matrix[36][200] * vector[36] +matrix[37][200] * vector[37] +matrix[38][200] * vector[38] +matrix[39][200] * vector[39] +matrix[40][200] * vector[40] +matrix[41][200] * vector[41] +matrix[42][200] * vector[42] +matrix[43][200] * vector[43] +matrix[44][200] * vector[44] +matrix[45][200] * vector[45] +matrix[46][200] * vector[46] +matrix[47][200] * vector[47] +matrix[48][200] * vector[48] +matrix[49][200] * vector[49] +matrix[50][200] * vector[50] +matrix[51][200] * vector[51] +matrix[52][200] * vector[52] +matrix[53][200] * vector[53] +matrix[54][200] * vector[54] +matrix[55][200] * vector[55] +matrix[56][200] * vector[56] +matrix[57][200] * vector[57] +matrix[58][200] * vector[58] +matrix[59][200] * vector[59] +matrix[60][200] * vector[60] +matrix[61][200] * vector[61] +matrix[62][200] * vector[62] +matrix[63][200] * vector[63] +matrix[64][200] * vector[64] +matrix[65][200] * vector[65] +matrix[66][200] * vector[66] +matrix[67][200] * vector[67] +matrix[68][200] * vector[68] +matrix[69][200] * vector[69] +matrix[70][200] * vector[70] +matrix[71][200] * vector[71] +matrix[72][200] * vector[72] +matrix[73][200] * vector[73] +matrix[74][200] * vector[74] +matrix[75][200] * vector[75] +matrix[76][200] * vector[76] +matrix[77][200] * vector[77] +matrix[78][200] * vector[78] +matrix[79][200] * vector[79] +matrix[80][200] * vector[80] +matrix[81][200] * vector[81] +matrix[82][200] * vector[82] +matrix[83][200] * vector[83] +matrix[84][200] * vector[84] +matrix[85][200] * vector[85] +matrix[86][200] * vector[86] +matrix[87][200] * vector[87] +matrix[88][200] * vector[88] +matrix[89][200] * vector[89] +matrix[90][200] * vector[90] +matrix[91][200] * vector[91] +matrix[92][200] * vector[92] +matrix[93][200] * vector[93] +matrix[94][200] * vector[94] +matrix[95][200] * vector[95] +matrix[96][200] * vector[96] +matrix[97][200] * vector[97] +matrix[98][200] * vector[98] +matrix[99][200] * vector[99] +b[200];
assign result[201] = matrix[0][201] * vector[0] +matrix[1][201] * vector[1] +matrix[2][201] * vector[2] +matrix[3][201] * vector[3] +matrix[4][201] * vector[4] +matrix[5][201] * vector[5] +matrix[6][201] * vector[6] +matrix[7][201] * vector[7] +matrix[8][201] * vector[8] +matrix[9][201] * vector[9] +matrix[10][201] * vector[10] +matrix[11][201] * vector[11] +matrix[12][201] * vector[12] +matrix[13][201] * vector[13] +matrix[14][201] * vector[14] +matrix[15][201] * vector[15] +matrix[16][201] * vector[16] +matrix[17][201] * vector[17] +matrix[18][201] * vector[18] +matrix[19][201] * vector[19] +matrix[20][201] * vector[20] +matrix[21][201] * vector[21] +matrix[22][201] * vector[22] +matrix[23][201] * vector[23] +matrix[24][201] * vector[24] +matrix[25][201] * vector[25] +matrix[26][201] * vector[26] +matrix[27][201] * vector[27] +matrix[28][201] * vector[28] +matrix[29][201] * vector[29] +matrix[30][201] * vector[30] +matrix[31][201] * vector[31] +matrix[32][201] * vector[32] +matrix[33][201] * vector[33] +matrix[34][201] * vector[34] +matrix[35][201] * vector[35] +matrix[36][201] * vector[36] +matrix[37][201] * vector[37] +matrix[38][201] * vector[38] +matrix[39][201] * vector[39] +matrix[40][201] * vector[40] +matrix[41][201] * vector[41] +matrix[42][201] * vector[42] +matrix[43][201] * vector[43] +matrix[44][201] * vector[44] +matrix[45][201] * vector[45] +matrix[46][201] * vector[46] +matrix[47][201] * vector[47] +matrix[48][201] * vector[48] +matrix[49][201] * vector[49] +matrix[50][201] * vector[50] +matrix[51][201] * vector[51] +matrix[52][201] * vector[52] +matrix[53][201] * vector[53] +matrix[54][201] * vector[54] +matrix[55][201] * vector[55] +matrix[56][201] * vector[56] +matrix[57][201] * vector[57] +matrix[58][201] * vector[58] +matrix[59][201] * vector[59] +matrix[60][201] * vector[60] +matrix[61][201] * vector[61] +matrix[62][201] * vector[62] +matrix[63][201] * vector[63] +matrix[64][201] * vector[64] +matrix[65][201] * vector[65] +matrix[66][201] * vector[66] +matrix[67][201] * vector[67] +matrix[68][201] * vector[68] +matrix[69][201] * vector[69] +matrix[70][201] * vector[70] +matrix[71][201] * vector[71] +matrix[72][201] * vector[72] +matrix[73][201] * vector[73] +matrix[74][201] * vector[74] +matrix[75][201] * vector[75] +matrix[76][201] * vector[76] +matrix[77][201] * vector[77] +matrix[78][201] * vector[78] +matrix[79][201] * vector[79] +matrix[80][201] * vector[80] +matrix[81][201] * vector[81] +matrix[82][201] * vector[82] +matrix[83][201] * vector[83] +matrix[84][201] * vector[84] +matrix[85][201] * vector[85] +matrix[86][201] * vector[86] +matrix[87][201] * vector[87] +matrix[88][201] * vector[88] +matrix[89][201] * vector[89] +matrix[90][201] * vector[90] +matrix[91][201] * vector[91] +matrix[92][201] * vector[92] +matrix[93][201] * vector[93] +matrix[94][201] * vector[94] +matrix[95][201] * vector[95] +matrix[96][201] * vector[96] +matrix[97][201] * vector[97] +matrix[98][201] * vector[98] +matrix[99][201] * vector[99] +b[201];
assign result[202] = matrix[0][202] * vector[0] +matrix[1][202] * vector[1] +matrix[2][202] * vector[2] +matrix[3][202] * vector[3] +matrix[4][202] * vector[4] +matrix[5][202] * vector[5] +matrix[6][202] * vector[6] +matrix[7][202] * vector[7] +matrix[8][202] * vector[8] +matrix[9][202] * vector[9] +matrix[10][202] * vector[10] +matrix[11][202] * vector[11] +matrix[12][202] * vector[12] +matrix[13][202] * vector[13] +matrix[14][202] * vector[14] +matrix[15][202] * vector[15] +matrix[16][202] * vector[16] +matrix[17][202] * vector[17] +matrix[18][202] * vector[18] +matrix[19][202] * vector[19] +matrix[20][202] * vector[20] +matrix[21][202] * vector[21] +matrix[22][202] * vector[22] +matrix[23][202] * vector[23] +matrix[24][202] * vector[24] +matrix[25][202] * vector[25] +matrix[26][202] * vector[26] +matrix[27][202] * vector[27] +matrix[28][202] * vector[28] +matrix[29][202] * vector[29] +matrix[30][202] * vector[30] +matrix[31][202] * vector[31] +matrix[32][202] * vector[32] +matrix[33][202] * vector[33] +matrix[34][202] * vector[34] +matrix[35][202] * vector[35] +matrix[36][202] * vector[36] +matrix[37][202] * vector[37] +matrix[38][202] * vector[38] +matrix[39][202] * vector[39] +matrix[40][202] * vector[40] +matrix[41][202] * vector[41] +matrix[42][202] * vector[42] +matrix[43][202] * vector[43] +matrix[44][202] * vector[44] +matrix[45][202] * vector[45] +matrix[46][202] * vector[46] +matrix[47][202] * vector[47] +matrix[48][202] * vector[48] +matrix[49][202] * vector[49] +matrix[50][202] * vector[50] +matrix[51][202] * vector[51] +matrix[52][202] * vector[52] +matrix[53][202] * vector[53] +matrix[54][202] * vector[54] +matrix[55][202] * vector[55] +matrix[56][202] * vector[56] +matrix[57][202] * vector[57] +matrix[58][202] * vector[58] +matrix[59][202] * vector[59] +matrix[60][202] * vector[60] +matrix[61][202] * vector[61] +matrix[62][202] * vector[62] +matrix[63][202] * vector[63] +matrix[64][202] * vector[64] +matrix[65][202] * vector[65] +matrix[66][202] * vector[66] +matrix[67][202] * vector[67] +matrix[68][202] * vector[68] +matrix[69][202] * vector[69] +matrix[70][202] * vector[70] +matrix[71][202] * vector[71] +matrix[72][202] * vector[72] +matrix[73][202] * vector[73] +matrix[74][202] * vector[74] +matrix[75][202] * vector[75] +matrix[76][202] * vector[76] +matrix[77][202] * vector[77] +matrix[78][202] * vector[78] +matrix[79][202] * vector[79] +matrix[80][202] * vector[80] +matrix[81][202] * vector[81] +matrix[82][202] * vector[82] +matrix[83][202] * vector[83] +matrix[84][202] * vector[84] +matrix[85][202] * vector[85] +matrix[86][202] * vector[86] +matrix[87][202] * vector[87] +matrix[88][202] * vector[88] +matrix[89][202] * vector[89] +matrix[90][202] * vector[90] +matrix[91][202] * vector[91] +matrix[92][202] * vector[92] +matrix[93][202] * vector[93] +matrix[94][202] * vector[94] +matrix[95][202] * vector[95] +matrix[96][202] * vector[96] +matrix[97][202] * vector[97] +matrix[98][202] * vector[98] +matrix[99][202] * vector[99] +b[202];
assign result[203] = matrix[0][203] * vector[0] +matrix[1][203] * vector[1] +matrix[2][203] * vector[2] +matrix[3][203] * vector[3] +matrix[4][203] * vector[4] +matrix[5][203] * vector[5] +matrix[6][203] * vector[6] +matrix[7][203] * vector[7] +matrix[8][203] * vector[8] +matrix[9][203] * vector[9] +matrix[10][203] * vector[10] +matrix[11][203] * vector[11] +matrix[12][203] * vector[12] +matrix[13][203] * vector[13] +matrix[14][203] * vector[14] +matrix[15][203] * vector[15] +matrix[16][203] * vector[16] +matrix[17][203] * vector[17] +matrix[18][203] * vector[18] +matrix[19][203] * vector[19] +matrix[20][203] * vector[20] +matrix[21][203] * vector[21] +matrix[22][203] * vector[22] +matrix[23][203] * vector[23] +matrix[24][203] * vector[24] +matrix[25][203] * vector[25] +matrix[26][203] * vector[26] +matrix[27][203] * vector[27] +matrix[28][203] * vector[28] +matrix[29][203] * vector[29] +matrix[30][203] * vector[30] +matrix[31][203] * vector[31] +matrix[32][203] * vector[32] +matrix[33][203] * vector[33] +matrix[34][203] * vector[34] +matrix[35][203] * vector[35] +matrix[36][203] * vector[36] +matrix[37][203] * vector[37] +matrix[38][203] * vector[38] +matrix[39][203] * vector[39] +matrix[40][203] * vector[40] +matrix[41][203] * vector[41] +matrix[42][203] * vector[42] +matrix[43][203] * vector[43] +matrix[44][203] * vector[44] +matrix[45][203] * vector[45] +matrix[46][203] * vector[46] +matrix[47][203] * vector[47] +matrix[48][203] * vector[48] +matrix[49][203] * vector[49] +matrix[50][203] * vector[50] +matrix[51][203] * vector[51] +matrix[52][203] * vector[52] +matrix[53][203] * vector[53] +matrix[54][203] * vector[54] +matrix[55][203] * vector[55] +matrix[56][203] * vector[56] +matrix[57][203] * vector[57] +matrix[58][203] * vector[58] +matrix[59][203] * vector[59] +matrix[60][203] * vector[60] +matrix[61][203] * vector[61] +matrix[62][203] * vector[62] +matrix[63][203] * vector[63] +matrix[64][203] * vector[64] +matrix[65][203] * vector[65] +matrix[66][203] * vector[66] +matrix[67][203] * vector[67] +matrix[68][203] * vector[68] +matrix[69][203] * vector[69] +matrix[70][203] * vector[70] +matrix[71][203] * vector[71] +matrix[72][203] * vector[72] +matrix[73][203] * vector[73] +matrix[74][203] * vector[74] +matrix[75][203] * vector[75] +matrix[76][203] * vector[76] +matrix[77][203] * vector[77] +matrix[78][203] * vector[78] +matrix[79][203] * vector[79] +matrix[80][203] * vector[80] +matrix[81][203] * vector[81] +matrix[82][203] * vector[82] +matrix[83][203] * vector[83] +matrix[84][203] * vector[84] +matrix[85][203] * vector[85] +matrix[86][203] * vector[86] +matrix[87][203] * vector[87] +matrix[88][203] * vector[88] +matrix[89][203] * vector[89] +matrix[90][203] * vector[90] +matrix[91][203] * vector[91] +matrix[92][203] * vector[92] +matrix[93][203] * vector[93] +matrix[94][203] * vector[94] +matrix[95][203] * vector[95] +matrix[96][203] * vector[96] +matrix[97][203] * vector[97] +matrix[98][203] * vector[98] +matrix[99][203] * vector[99] +b[203];
assign result[204] = matrix[0][204] * vector[0] +matrix[1][204] * vector[1] +matrix[2][204] * vector[2] +matrix[3][204] * vector[3] +matrix[4][204] * vector[4] +matrix[5][204] * vector[5] +matrix[6][204] * vector[6] +matrix[7][204] * vector[7] +matrix[8][204] * vector[8] +matrix[9][204] * vector[9] +matrix[10][204] * vector[10] +matrix[11][204] * vector[11] +matrix[12][204] * vector[12] +matrix[13][204] * vector[13] +matrix[14][204] * vector[14] +matrix[15][204] * vector[15] +matrix[16][204] * vector[16] +matrix[17][204] * vector[17] +matrix[18][204] * vector[18] +matrix[19][204] * vector[19] +matrix[20][204] * vector[20] +matrix[21][204] * vector[21] +matrix[22][204] * vector[22] +matrix[23][204] * vector[23] +matrix[24][204] * vector[24] +matrix[25][204] * vector[25] +matrix[26][204] * vector[26] +matrix[27][204] * vector[27] +matrix[28][204] * vector[28] +matrix[29][204] * vector[29] +matrix[30][204] * vector[30] +matrix[31][204] * vector[31] +matrix[32][204] * vector[32] +matrix[33][204] * vector[33] +matrix[34][204] * vector[34] +matrix[35][204] * vector[35] +matrix[36][204] * vector[36] +matrix[37][204] * vector[37] +matrix[38][204] * vector[38] +matrix[39][204] * vector[39] +matrix[40][204] * vector[40] +matrix[41][204] * vector[41] +matrix[42][204] * vector[42] +matrix[43][204] * vector[43] +matrix[44][204] * vector[44] +matrix[45][204] * vector[45] +matrix[46][204] * vector[46] +matrix[47][204] * vector[47] +matrix[48][204] * vector[48] +matrix[49][204] * vector[49] +matrix[50][204] * vector[50] +matrix[51][204] * vector[51] +matrix[52][204] * vector[52] +matrix[53][204] * vector[53] +matrix[54][204] * vector[54] +matrix[55][204] * vector[55] +matrix[56][204] * vector[56] +matrix[57][204] * vector[57] +matrix[58][204] * vector[58] +matrix[59][204] * vector[59] +matrix[60][204] * vector[60] +matrix[61][204] * vector[61] +matrix[62][204] * vector[62] +matrix[63][204] * vector[63] +matrix[64][204] * vector[64] +matrix[65][204] * vector[65] +matrix[66][204] * vector[66] +matrix[67][204] * vector[67] +matrix[68][204] * vector[68] +matrix[69][204] * vector[69] +matrix[70][204] * vector[70] +matrix[71][204] * vector[71] +matrix[72][204] * vector[72] +matrix[73][204] * vector[73] +matrix[74][204] * vector[74] +matrix[75][204] * vector[75] +matrix[76][204] * vector[76] +matrix[77][204] * vector[77] +matrix[78][204] * vector[78] +matrix[79][204] * vector[79] +matrix[80][204] * vector[80] +matrix[81][204] * vector[81] +matrix[82][204] * vector[82] +matrix[83][204] * vector[83] +matrix[84][204] * vector[84] +matrix[85][204] * vector[85] +matrix[86][204] * vector[86] +matrix[87][204] * vector[87] +matrix[88][204] * vector[88] +matrix[89][204] * vector[89] +matrix[90][204] * vector[90] +matrix[91][204] * vector[91] +matrix[92][204] * vector[92] +matrix[93][204] * vector[93] +matrix[94][204] * vector[94] +matrix[95][204] * vector[95] +matrix[96][204] * vector[96] +matrix[97][204] * vector[97] +matrix[98][204] * vector[98] +matrix[99][204] * vector[99] +b[204];
assign result[205] = matrix[0][205] * vector[0] +matrix[1][205] * vector[1] +matrix[2][205] * vector[2] +matrix[3][205] * vector[3] +matrix[4][205] * vector[4] +matrix[5][205] * vector[5] +matrix[6][205] * vector[6] +matrix[7][205] * vector[7] +matrix[8][205] * vector[8] +matrix[9][205] * vector[9] +matrix[10][205] * vector[10] +matrix[11][205] * vector[11] +matrix[12][205] * vector[12] +matrix[13][205] * vector[13] +matrix[14][205] * vector[14] +matrix[15][205] * vector[15] +matrix[16][205] * vector[16] +matrix[17][205] * vector[17] +matrix[18][205] * vector[18] +matrix[19][205] * vector[19] +matrix[20][205] * vector[20] +matrix[21][205] * vector[21] +matrix[22][205] * vector[22] +matrix[23][205] * vector[23] +matrix[24][205] * vector[24] +matrix[25][205] * vector[25] +matrix[26][205] * vector[26] +matrix[27][205] * vector[27] +matrix[28][205] * vector[28] +matrix[29][205] * vector[29] +matrix[30][205] * vector[30] +matrix[31][205] * vector[31] +matrix[32][205] * vector[32] +matrix[33][205] * vector[33] +matrix[34][205] * vector[34] +matrix[35][205] * vector[35] +matrix[36][205] * vector[36] +matrix[37][205] * vector[37] +matrix[38][205] * vector[38] +matrix[39][205] * vector[39] +matrix[40][205] * vector[40] +matrix[41][205] * vector[41] +matrix[42][205] * vector[42] +matrix[43][205] * vector[43] +matrix[44][205] * vector[44] +matrix[45][205] * vector[45] +matrix[46][205] * vector[46] +matrix[47][205] * vector[47] +matrix[48][205] * vector[48] +matrix[49][205] * vector[49] +matrix[50][205] * vector[50] +matrix[51][205] * vector[51] +matrix[52][205] * vector[52] +matrix[53][205] * vector[53] +matrix[54][205] * vector[54] +matrix[55][205] * vector[55] +matrix[56][205] * vector[56] +matrix[57][205] * vector[57] +matrix[58][205] * vector[58] +matrix[59][205] * vector[59] +matrix[60][205] * vector[60] +matrix[61][205] * vector[61] +matrix[62][205] * vector[62] +matrix[63][205] * vector[63] +matrix[64][205] * vector[64] +matrix[65][205] * vector[65] +matrix[66][205] * vector[66] +matrix[67][205] * vector[67] +matrix[68][205] * vector[68] +matrix[69][205] * vector[69] +matrix[70][205] * vector[70] +matrix[71][205] * vector[71] +matrix[72][205] * vector[72] +matrix[73][205] * vector[73] +matrix[74][205] * vector[74] +matrix[75][205] * vector[75] +matrix[76][205] * vector[76] +matrix[77][205] * vector[77] +matrix[78][205] * vector[78] +matrix[79][205] * vector[79] +matrix[80][205] * vector[80] +matrix[81][205] * vector[81] +matrix[82][205] * vector[82] +matrix[83][205] * vector[83] +matrix[84][205] * vector[84] +matrix[85][205] * vector[85] +matrix[86][205] * vector[86] +matrix[87][205] * vector[87] +matrix[88][205] * vector[88] +matrix[89][205] * vector[89] +matrix[90][205] * vector[90] +matrix[91][205] * vector[91] +matrix[92][205] * vector[92] +matrix[93][205] * vector[93] +matrix[94][205] * vector[94] +matrix[95][205] * vector[95] +matrix[96][205] * vector[96] +matrix[97][205] * vector[97] +matrix[98][205] * vector[98] +matrix[99][205] * vector[99] +b[205];
assign result[206] = matrix[0][206] * vector[0] +matrix[1][206] * vector[1] +matrix[2][206] * vector[2] +matrix[3][206] * vector[3] +matrix[4][206] * vector[4] +matrix[5][206] * vector[5] +matrix[6][206] * vector[6] +matrix[7][206] * vector[7] +matrix[8][206] * vector[8] +matrix[9][206] * vector[9] +matrix[10][206] * vector[10] +matrix[11][206] * vector[11] +matrix[12][206] * vector[12] +matrix[13][206] * vector[13] +matrix[14][206] * vector[14] +matrix[15][206] * vector[15] +matrix[16][206] * vector[16] +matrix[17][206] * vector[17] +matrix[18][206] * vector[18] +matrix[19][206] * vector[19] +matrix[20][206] * vector[20] +matrix[21][206] * vector[21] +matrix[22][206] * vector[22] +matrix[23][206] * vector[23] +matrix[24][206] * vector[24] +matrix[25][206] * vector[25] +matrix[26][206] * vector[26] +matrix[27][206] * vector[27] +matrix[28][206] * vector[28] +matrix[29][206] * vector[29] +matrix[30][206] * vector[30] +matrix[31][206] * vector[31] +matrix[32][206] * vector[32] +matrix[33][206] * vector[33] +matrix[34][206] * vector[34] +matrix[35][206] * vector[35] +matrix[36][206] * vector[36] +matrix[37][206] * vector[37] +matrix[38][206] * vector[38] +matrix[39][206] * vector[39] +matrix[40][206] * vector[40] +matrix[41][206] * vector[41] +matrix[42][206] * vector[42] +matrix[43][206] * vector[43] +matrix[44][206] * vector[44] +matrix[45][206] * vector[45] +matrix[46][206] * vector[46] +matrix[47][206] * vector[47] +matrix[48][206] * vector[48] +matrix[49][206] * vector[49] +matrix[50][206] * vector[50] +matrix[51][206] * vector[51] +matrix[52][206] * vector[52] +matrix[53][206] * vector[53] +matrix[54][206] * vector[54] +matrix[55][206] * vector[55] +matrix[56][206] * vector[56] +matrix[57][206] * vector[57] +matrix[58][206] * vector[58] +matrix[59][206] * vector[59] +matrix[60][206] * vector[60] +matrix[61][206] * vector[61] +matrix[62][206] * vector[62] +matrix[63][206] * vector[63] +matrix[64][206] * vector[64] +matrix[65][206] * vector[65] +matrix[66][206] * vector[66] +matrix[67][206] * vector[67] +matrix[68][206] * vector[68] +matrix[69][206] * vector[69] +matrix[70][206] * vector[70] +matrix[71][206] * vector[71] +matrix[72][206] * vector[72] +matrix[73][206] * vector[73] +matrix[74][206] * vector[74] +matrix[75][206] * vector[75] +matrix[76][206] * vector[76] +matrix[77][206] * vector[77] +matrix[78][206] * vector[78] +matrix[79][206] * vector[79] +matrix[80][206] * vector[80] +matrix[81][206] * vector[81] +matrix[82][206] * vector[82] +matrix[83][206] * vector[83] +matrix[84][206] * vector[84] +matrix[85][206] * vector[85] +matrix[86][206] * vector[86] +matrix[87][206] * vector[87] +matrix[88][206] * vector[88] +matrix[89][206] * vector[89] +matrix[90][206] * vector[90] +matrix[91][206] * vector[91] +matrix[92][206] * vector[92] +matrix[93][206] * vector[93] +matrix[94][206] * vector[94] +matrix[95][206] * vector[95] +matrix[96][206] * vector[96] +matrix[97][206] * vector[97] +matrix[98][206] * vector[98] +matrix[99][206] * vector[99] +b[206];
assign result[207] = matrix[0][207] * vector[0] +matrix[1][207] * vector[1] +matrix[2][207] * vector[2] +matrix[3][207] * vector[3] +matrix[4][207] * vector[4] +matrix[5][207] * vector[5] +matrix[6][207] * vector[6] +matrix[7][207] * vector[7] +matrix[8][207] * vector[8] +matrix[9][207] * vector[9] +matrix[10][207] * vector[10] +matrix[11][207] * vector[11] +matrix[12][207] * vector[12] +matrix[13][207] * vector[13] +matrix[14][207] * vector[14] +matrix[15][207] * vector[15] +matrix[16][207] * vector[16] +matrix[17][207] * vector[17] +matrix[18][207] * vector[18] +matrix[19][207] * vector[19] +matrix[20][207] * vector[20] +matrix[21][207] * vector[21] +matrix[22][207] * vector[22] +matrix[23][207] * vector[23] +matrix[24][207] * vector[24] +matrix[25][207] * vector[25] +matrix[26][207] * vector[26] +matrix[27][207] * vector[27] +matrix[28][207] * vector[28] +matrix[29][207] * vector[29] +matrix[30][207] * vector[30] +matrix[31][207] * vector[31] +matrix[32][207] * vector[32] +matrix[33][207] * vector[33] +matrix[34][207] * vector[34] +matrix[35][207] * vector[35] +matrix[36][207] * vector[36] +matrix[37][207] * vector[37] +matrix[38][207] * vector[38] +matrix[39][207] * vector[39] +matrix[40][207] * vector[40] +matrix[41][207] * vector[41] +matrix[42][207] * vector[42] +matrix[43][207] * vector[43] +matrix[44][207] * vector[44] +matrix[45][207] * vector[45] +matrix[46][207] * vector[46] +matrix[47][207] * vector[47] +matrix[48][207] * vector[48] +matrix[49][207] * vector[49] +matrix[50][207] * vector[50] +matrix[51][207] * vector[51] +matrix[52][207] * vector[52] +matrix[53][207] * vector[53] +matrix[54][207] * vector[54] +matrix[55][207] * vector[55] +matrix[56][207] * vector[56] +matrix[57][207] * vector[57] +matrix[58][207] * vector[58] +matrix[59][207] * vector[59] +matrix[60][207] * vector[60] +matrix[61][207] * vector[61] +matrix[62][207] * vector[62] +matrix[63][207] * vector[63] +matrix[64][207] * vector[64] +matrix[65][207] * vector[65] +matrix[66][207] * vector[66] +matrix[67][207] * vector[67] +matrix[68][207] * vector[68] +matrix[69][207] * vector[69] +matrix[70][207] * vector[70] +matrix[71][207] * vector[71] +matrix[72][207] * vector[72] +matrix[73][207] * vector[73] +matrix[74][207] * vector[74] +matrix[75][207] * vector[75] +matrix[76][207] * vector[76] +matrix[77][207] * vector[77] +matrix[78][207] * vector[78] +matrix[79][207] * vector[79] +matrix[80][207] * vector[80] +matrix[81][207] * vector[81] +matrix[82][207] * vector[82] +matrix[83][207] * vector[83] +matrix[84][207] * vector[84] +matrix[85][207] * vector[85] +matrix[86][207] * vector[86] +matrix[87][207] * vector[87] +matrix[88][207] * vector[88] +matrix[89][207] * vector[89] +matrix[90][207] * vector[90] +matrix[91][207] * vector[91] +matrix[92][207] * vector[92] +matrix[93][207] * vector[93] +matrix[94][207] * vector[94] +matrix[95][207] * vector[95] +matrix[96][207] * vector[96] +matrix[97][207] * vector[97] +matrix[98][207] * vector[98] +matrix[99][207] * vector[99] +b[207];
assign result[208] = matrix[0][208] * vector[0] +matrix[1][208] * vector[1] +matrix[2][208] * vector[2] +matrix[3][208] * vector[3] +matrix[4][208] * vector[4] +matrix[5][208] * vector[5] +matrix[6][208] * vector[6] +matrix[7][208] * vector[7] +matrix[8][208] * vector[8] +matrix[9][208] * vector[9] +matrix[10][208] * vector[10] +matrix[11][208] * vector[11] +matrix[12][208] * vector[12] +matrix[13][208] * vector[13] +matrix[14][208] * vector[14] +matrix[15][208] * vector[15] +matrix[16][208] * vector[16] +matrix[17][208] * vector[17] +matrix[18][208] * vector[18] +matrix[19][208] * vector[19] +matrix[20][208] * vector[20] +matrix[21][208] * vector[21] +matrix[22][208] * vector[22] +matrix[23][208] * vector[23] +matrix[24][208] * vector[24] +matrix[25][208] * vector[25] +matrix[26][208] * vector[26] +matrix[27][208] * vector[27] +matrix[28][208] * vector[28] +matrix[29][208] * vector[29] +matrix[30][208] * vector[30] +matrix[31][208] * vector[31] +matrix[32][208] * vector[32] +matrix[33][208] * vector[33] +matrix[34][208] * vector[34] +matrix[35][208] * vector[35] +matrix[36][208] * vector[36] +matrix[37][208] * vector[37] +matrix[38][208] * vector[38] +matrix[39][208] * vector[39] +matrix[40][208] * vector[40] +matrix[41][208] * vector[41] +matrix[42][208] * vector[42] +matrix[43][208] * vector[43] +matrix[44][208] * vector[44] +matrix[45][208] * vector[45] +matrix[46][208] * vector[46] +matrix[47][208] * vector[47] +matrix[48][208] * vector[48] +matrix[49][208] * vector[49] +matrix[50][208] * vector[50] +matrix[51][208] * vector[51] +matrix[52][208] * vector[52] +matrix[53][208] * vector[53] +matrix[54][208] * vector[54] +matrix[55][208] * vector[55] +matrix[56][208] * vector[56] +matrix[57][208] * vector[57] +matrix[58][208] * vector[58] +matrix[59][208] * vector[59] +matrix[60][208] * vector[60] +matrix[61][208] * vector[61] +matrix[62][208] * vector[62] +matrix[63][208] * vector[63] +matrix[64][208] * vector[64] +matrix[65][208] * vector[65] +matrix[66][208] * vector[66] +matrix[67][208] * vector[67] +matrix[68][208] * vector[68] +matrix[69][208] * vector[69] +matrix[70][208] * vector[70] +matrix[71][208] * vector[71] +matrix[72][208] * vector[72] +matrix[73][208] * vector[73] +matrix[74][208] * vector[74] +matrix[75][208] * vector[75] +matrix[76][208] * vector[76] +matrix[77][208] * vector[77] +matrix[78][208] * vector[78] +matrix[79][208] * vector[79] +matrix[80][208] * vector[80] +matrix[81][208] * vector[81] +matrix[82][208] * vector[82] +matrix[83][208] * vector[83] +matrix[84][208] * vector[84] +matrix[85][208] * vector[85] +matrix[86][208] * vector[86] +matrix[87][208] * vector[87] +matrix[88][208] * vector[88] +matrix[89][208] * vector[89] +matrix[90][208] * vector[90] +matrix[91][208] * vector[91] +matrix[92][208] * vector[92] +matrix[93][208] * vector[93] +matrix[94][208] * vector[94] +matrix[95][208] * vector[95] +matrix[96][208] * vector[96] +matrix[97][208] * vector[97] +matrix[98][208] * vector[98] +matrix[99][208] * vector[99] +b[208];
assign result[209] = matrix[0][209] * vector[0] +matrix[1][209] * vector[1] +matrix[2][209] * vector[2] +matrix[3][209] * vector[3] +matrix[4][209] * vector[4] +matrix[5][209] * vector[5] +matrix[6][209] * vector[6] +matrix[7][209] * vector[7] +matrix[8][209] * vector[8] +matrix[9][209] * vector[9] +matrix[10][209] * vector[10] +matrix[11][209] * vector[11] +matrix[12][209] * vector[12] +matrix[13][209] * vector[13] +matrix[14][209] * vector[14] +matrix[15][209] * vector[15] +matrix[16][209] * vector[16] +matrix[17][209] * vector[17] +matrix[18][209] * vector[18] +matrix[19][209] * vector[19] +matrix[20][209] * vector[20] +matrix[21][209] * vector[21] +matrix[22][209] * vector[22] +matrix[23][209] * vector[23] +matrix[24][209] * vector[24] +matrix[25][209] * vector[25] +matrix[26][209] * vector[26] +matrix[27][209] * vector[27] +matrix[28][209] * vector[28] +matrix[29][209] * vector[29] +matrix[30][209] * vector[30] +matrix[31][209] * vector[31] +matrix[32][209] * vector[32] +matrix[33][209] * vector[33] +matrix[34][209] * vector[34] +matrix[35][209] * vector[35] +matrix[36][209] * vector[36] +matrix[37][209] * vector[37] +matrix[38][209] * vector[38] +matrix[39][209] * vector[39] +matrix[40][209] * vector[40] +matrix[41][209] * vector[41] +matrix[42][209] * vector[42] +matrix[43][209] * vector[43] +matrix[44][209] * vector[44] +matrix[45][209] * vector[45] +matrix[46][209] * vector[46] +matrix[47][209] * vector[47] +matrix[48][209] * vector[48] +matrix[49][209] * vector[49] +matrix[50][209] * vector[50] +matrix[51][209] * vector[51] +matrix[52][209] * vector[52] +matrix[53][209] * vector[53] +matrix[54][209] * vector[54] +matrix[55][209] * vector[55] +matrix[56][209] * vector[56] +matrix[57][209] * vector[57] +matrix[58][209] * vector[58] +matrix[59][209] * vector[59] +matrix[60][209] * vector[60] +matrix[61][209] * vector[61] +matrix[62][209] * vector[62] +matrix[63][209] * vector[63] +matrix[64][209] * vector[64] +matrix[65][209] * vector[65] +matrix[66][209] * vector[66] +matrix[67][209] * vector[67] +matrix[68][209] * vector[68] +matrix[69][209] * vector[69] +matrix[70][209] * vector[70] +matrix[71][209] * vector[71] +matrix[72][209] * vector[72] +matrix[73][209] * vector[73] +matrix[74][209] * vector[74] +matrix[75][209] * vector[75] +matrix[76][209] * vector[76] +matrix[77][209] * vector[77] +matrix[78][209] * vector[78] +matrix[79][209] * vector[79] +matrix[80][209] * vector[80] +matrix[81][209] * vector[81] +matrix[82][209] * vector[82] +matrix[83][209] * vector[83] +matrix[84][209] * vector[84] +matrix[85][209] * vector[85] +matrix[86][209] * vector[86] +matrix[87][209] * vector[87] +matrix[88][209] * vector[88] +matrix[89][209] * vector[89] +matrix[90][209] * vector[90] +matrix[91][209] * vector[91] +matrix[92][209] * vector[92] +matrix[93][209] * vector[93] +matrix[94][209] * vector[94] +matrix[95][209] * vector[95] +matrix[96][209] * vector[96] +matrix[97][209] * vector[97] +matrix[98][209] * vector[98] +matrix[99][209] * vector[99] +b[209];
assign result[210] = matrix[0][210] * vector[0] +matrix[1][210] * vector[1] +matrix[2][210] * vector[2] +matrix[3][210] * vector[3] +matrix[4][210] * vector[4] +matrix[5][210] * vector[5] +matrix[6][210] * vector[6] +matrix[7][210] * vector[7] +matrix[8][210] * vector[8] +matrix[9][210] * vector[9] +matrix[10][210] * vector[10] +matrix[11][210] * vector[11] +matrix[12][210] * vector[12] +matrix[13][210] * vector[13] +matrix[14][210] * vector[14] +matrix[15][210] * vector[15] +matrix[16][210] * vector[16] +matrix[17][210] * vector[17] +matrix[18][210] * vector[18] +matrix[19][210] * vector[19] +matrix[20][210] * vector[20] +matrix[21][210] * vector[21] +matrix[22][210] * vector[22] +matrix[23][210] * vector[23] +matrix[24][210] * vector[24] +matrix[25][210] * vector[25] +matrix[26][210] * vector[26] +matrix[27][210] * vector[27] +matrix[28][210] * vector[28] +matrix[29][210] * vector[29] +matrix[30][210] * vector[30] +matrix[31][210] * vector[31] +matrix[32][210] * vector[32] +matrix[33][210] * vector[33] +matrix[34][210] * vector[34] +matrix[35][210] * vector[35] +matrix[36][210] * vector[36] +matrix[37][210] * vector[37] +matrix[38][210] * vector[38] +matrix[39][210] * vector[39] +matrix[40][210] * vector[40] +matrix[41][210] * vector[41] +matrix[42][210] * vector[42] +matrix[43][210] * vector[43] +matrix[44][210] * vector[44] +matrix[45][210] * vector[45] +matrix[46][210] * vector[46] +matrix[47][210] * vector[47] +matrix[48][210] * vector[48] +matrix[49][210] * vector[49] +matrix[50][210] * vector[50] +matrix[51][210] * vector[51] +matrix[52][210] * vector[52] +matrix[53][210] * vector[53] +matrix[54][210] * vector[54] +matrix[55][210] * vector[55] +matrix[56][210] * vector[56] +matrix[57][210] * vector[57] +matrix[58][210] * vector[58] +matrix[59][210] * vector[59] +matrix[60][210] * vector[60] +matrix[61][210] * vector[61] +matrix[62][210] * vector[62] +matrix[63][210] * vector[63] +matrix[64][210] * vector[64] +matrix[65][210] * vector[65] +matrix[66][210] * vector[66] +matrix[67][210] * vector[67] +matrix[68][210] * vector[68] +matrix[69][210] * vector[69] +matrix[70][210] * vector[70] +matrix[71][210] * vector[71] +matrix[72][210] * vector[72] +matrix[73][210] * vector[73] +matrix[74][210] * vector[74] +matrix[75][210] * vector[75] +matrix[76][210] * vector[76] +matrix[77][210] * vector[77] +matrix[78][210] * vector[78] +matrix[79][210] * vector[79] +matrix[80][210] * vector[80] +matrix[81][210] * vector[81] +matrix[82][210] * vector[82] +matrix[83][210] * vector[83] +matrix[84][210] * vector[84] +matrix[85][210] * vector[85] +matrix[86][210] * vector[86] +matrix[87][210] * vector[87] +matrix[88][210] * vector[88] +matrix[89][210] * vector[89] +matrix[90][210] * vector[90] +matrix[91][210] * vector[91] +matrix[92][210] * vector[92] +matrix[93][210] * vector[93] +matrix[94][210] * vector[94] +matrix[95][210] * vector[95] +matrix[96][210] * vector[96] +matrix[97][210] * vector[97] +matrix[98][210] * vector[98] +matrix[99][210] * vector[99] +b[210];
assign result[211] = matrix[0][211] * vector[0] +matrix[1][211] * vector[1] +matrix[2][211] * vector[2] +matrix[3][211] * vector[3] +matrix[4][211] * vector[4] +matrix[5][211] * vector[5] +matrix[6][211] * vector[6] +matrix[7][211] * vector[7] +matrix[8][211] * vector[8] +matrix[9][211] * vector[9] +matrix[10][211] * vector[10] +matrix[11][211] * vector[11] +matrix[12][211] * vector[12] +matrix[13][211] * vector[13] +matrix[14][211] * vector[14] +matrix[15][211] * vector[15] +matrix[16][211] * vector[16] +matrix[17][211] * vector[17] +matrix[18][211] * vector[18] +matrix[19][211] * vector[19] +matrix[20][211] * vector[20] +matrix[21][211] * vector[21] +matrix[22][211] * vector[22] +matrix[23][211] * vector[23] +matrix[24][211] * vector[24] +matrix[25][211] * vector[25] +matrix[26][211] * vector[26] +matrix[27][211] * vector[27] +matrix[28][211] * vector[28] +matrix[29][211] * vector[29] +matrix[30][211] * vector[30] +matrix[31][211] * vector[31] +matrix[32][211] * vector[32] +matrix[33][211] * vector[33] +matrix[34][211] * vector[34] +matrix[35][211] * vector[35] +matrix[36][211] * vector[36] +matrix[37][211] * vector[37] +matrix[38][211] * vector[38] +matrix[39][211] * vector[39] +matrix[40][211] * vector[40] +matrix[41][211] * vector[41] +matrix[42][211] * vector[42] +matrix[43][211] * vector[43] +matrix[44][211] * vector[44] +matrix[45][211] * vector[45] +matrix[46][211] * vector[46] +matrix[47][211] * vector[47] +matrix[48][211] * vector[48] +matrix[49][211] * vector[49] +matrix[50][211] * vector[50] +matrix[51][211] * vector[51] +matrix[52][211] * vector[52] +matrix[53][211] * vector[53] +matrix[54][211] * vector[54] +matrix[55][211] * vector[55] +matrix[56][211] * vector[56] +matrix[57][211] * vector[57] +matrix[58][211] * vector[58] +matrix[59][211] * vector[59] +matrix[60][211] * vector[60] +matrix[61][211] * vector[61] +matrix[62][211] * vector[62] +matrix[63][211] * vector[63] +matrix[64][211] * vector[64] +matrix[65][211] * vector[65] +matrix[66][211] * vector[66] +matrix[67][211] * vector[67] +matrix[68][211] * vector[68] +matrix[69][211] * vector[69] +matrix[70][211] * vector[70] +matrix[71][211] * vector[71] +matrix[72][211] * vector[72] +matrix[73][211] * vector[73] +matrix[74][211] * vector[74] +matrix[75][211] * vector[75] +matrix[76][211] * vector[76] +matrix[77][211] * vector[77] +matrix[78][211] * vector[78] +matrix[79][211] * vector[79] +matrix[80][211] * vector[80] +matrix[81][211] * vector[81] +matrix[82][211] * vector[82] +matrix[83][211] * vector[83] +matrix[84][211] * vector[84] +matrix[85][211] * vector[85] +matrix[86][211] * vector[86] +matrix[87][211] * vector[87] +matrix[88][211] * vector[88] +matrix[89][211] * vector[89] +matrix[90][211] * vector[90] +matrix[91][211] * vector[91] +matrix[92][211] * vector[92] +matrix[93][211] * vector[93] +matrix[94][211] * vector[94] +matrix[95][211] * vector[95] +matrix[96][211] * vector[96] +matrix[97][211] * vector[97] +matrix[98][211] * vector[98] +matrix[99][211] * vector[99] +b[211];
assign result[212] = matrix[0][212] * vector[0] +matrix[1][212] * vector[1] +matrix[2][212] * vector[2] +matrix[3][212] * vector[3] +matrix[4][212] * vector[4] +matrix[5][212] * vector[5] +matrix[6][212] * vector[6] +matrix[7][212] * vector[7] +matrix[8][212] * vector[8] +matrix[9][212] * vector[9] +matrix[10][212] * vector[10] +matrix[11][212] * vector[11] +matrix[12][212] * vector[12] +matrix[13][212] * vector[13] +matrix[14][212] * vector[14] +matrix[15][212] * vector[15] +matrix[16][212] * vector[16] +matrix[17][212] * vector[17] +matrix[18][212] * vector[18] +matrix[19][212] * vector[19] +matrix[20][212] * vector[20] +matrix[21][212] * vector[21] +matrix[22][212] * vector[22] +matrix[23][212] * vector[23] +matrix[24][212] * vector[24] +matrix[25][212] * vector[25] +matrix[26][212] * vector[26] +matrix[27][212] * vector[27] +matrix[28][212] * vector[28] +matrix[29][212] * vector[29] +matrix[30][212] * vector[30] +matrix[31][212] * vector[31] +matrix[32][212] * vector[32] +matrix[33][212] * vector[33] +matrix[34][212] * vector[34] +matrix[35][212] * vector[35] +matrix[36][212] * vector[36] +matrix[37][212] * vector[37] +matrix[38][212] * vector[38] +matrix[39][212] * vector[39] +matrix[40][212] * vector[40] +matrix[41][212] * vector[41] +matrix[42][212] * vector[42] +matrix[43][212] * vector[43] +matrix[44][212] * vector[44] +matrix[45][212] * vector[45] +matrix[46][212] * vector[46] +matrix[47][212] * vector[47] +matrix[48][212] * vector[48] +matrix[49][212] * vector[49] +matrix[50][212] * vector[50] +matrix[51][212] * vector[51] +matrix[52][212] * vector[52] +matrix[53][212] * vector[53] +matrix[54][212] * vector[54] +matrix[55][212] * vector[55] +matrix[56][212] * vector[56] +matrix[57][212] * vector[57] +matrix[58][212] * vector[58] +matrix[59][212] * vector[59] +matrix[60][212] * vector[60] +matrix[61][212] * vector[61] +matrix[62][212] * vector[62] +matrix[63][212] * vector[63] +matrix[64][212] * vector[64] +matrix[65][212] * vector[65] +matrix[66][212] * vector[66] +matrix[67][212] * vector[67] +matrix[68][212] * vector[68] +matrix[69][212] * vector[69] +matrix[70][212] * vector[70] +matrix[71][212] * vector[71] +matrix[72][212] * vector[72] +matrix[73][212] * vector[73] +matrix[74][212] * vector[74] +matrix[75][212] * vector[75] +matrix[76][212] * vector[76] +matrix[77][212] * vector[77] +matrix[78][212] * vector[78] +matrix[79][212] * vector[79] +matrix[80][212] * vector[80] +matrix[81][212] * vector[81] +matrix[82][212] * vector[82] +matrix[83][212] * vector[83] +matrix[84][212] * vector[84] +matrix[85][212] * vector[85] +matrix[86][212] * vector[86] +matrix[87][212] * vector[87] +matrix[88][212] * vector[88] +matrix[89][212] * vector[89] +matrix[90][212] * vector[90] +matrix[91][212] * vector[91] +matrix[92][212] * vector[92] +matrix[93][212] * vector[93] +matrix[94][212] * vector[94] +matrix[95][212] * vector[95] +matrix[96][212] * vector[96] +matrix[97][212] * vector[97] +matrix[98][212] * vector[98] +matrix[99][212] * vector[99] +b[212];
assign result[213] = matrix[0][213] * vector[0] +matrix[1][213] * vector[1] +matrix[2][213] * vector[2] +matrix[3][213] * vector[3] +matrix[4][213] * vector[4] +matrix[5][213] * vector[5] +matrix[6][213] * vector[6] +matrix[7][213] * vector[7] +matrix[8][213] * vector[8] +matrix[9][213] * vector[9] +matrix[10][213] * vector[10] +matrix[11][213] * vector[11] +matrix[12][213] * vector[12] +matrix[13][213] * vector[13] +matrix[14][213] * vector[14] +matrix[15][213] * vector[15] +matrix[16][213] * vector[16] +matrix[17][213] * vector[17] +matrix[18][213] * vector[18] +matrix[19][213] * vector[19] +matrix[20][213] * vector[20] +matrix[21][213] * vector[21] +matrix[22][213] * vector[22] +matrix[23][213] * vector[23] +matrix[24][213] * vector[24] +matrix[25][213] * vector[25] +matrix[26][213] * vector[26] +matrix[27][213] * vector[27] +matrix[28][213] * vector[28] +matrix[29][213] * vector[29] +matrix[30][213] * vector[30] +matrix[31][213] * vector[31] +matrix[32][213] * vector[32] +matrix[33][213] * vector[33] +matrix[34][213] * vector[34] +matrix[35][213] * vector[35] +matrix[36][213] * vector[36] +matrix[37][213] * vector[37] +matrix[38][213] * vector[38] +matrix[39][213] * vector[39] +matrix[40][213] * vector[40] +matrix[41][213] * vector[41] +matrix[42][213] * vector[42] +matrix[43][213] * vector[43] +matrix[44][213] * vector[44] +matrix[45][213] * vector[45] +matrix[46][213] * vector[46] +matrix[47][213] * vector[47] +matrix[48][213] * vector[48] +matrix[49][213] * vector[49] +matrix[50][213] * vector[50] +matrix[51][213] * vector[51] +matrix[52][213] * vector[52] +matrix[53][213] * vector[53] +matrix[54][213] * vector[54] +matrix[55][213] * vector[55] +matrix[56][213] * vector[56] +matrix[57][213] * vector[57] +matrix[58][213] * vector[58] +matrix[59][213] * vector[59] +matrix[60][213] * vector[60] +matrix[61][213] * vector[61] +matrix[62][213] * vector[62] +matrix[63][213] * vector[63] +matrix[64][213] * vector[64] +matrix[65][213] * vector[65] +matrix[66][213] * vector[66] +matrix[67][213] * vector[67] +matrix[68][213] * vector[68] +matrix[69][213] * vector[69] +matrix[70][213] * vector[70] +matrix[71][213] * vector[71] +matrix[72][213] * vector[72] +matrix[73][213] * vector[73] +matrix[74][213] * vector[74] +matrix[75][213] * vector[75] +matrix[76][213] * vector[76] +matrix[77][213] * vector[77] +matrix[78][213] * vector[78] +matrix[79][213] * vector[79] +matrix[80][213] * vector[80] +matrix[81][213] * vector[81] +matrix[82][213] * vector[82] +matrix[83][213] * vector[83] +matrix[84][213] * vector[84] +matrix[85][213] * vector[85] +matrix[86][213] * vector[86] +matrix[87][213] * vector[87] +matrix[88][213] * vector[88] +matrix[89][213] * vector[89] +matrix[90][213] * vector[90] +matrix[91][213] * vector[91] +matrix[92][213] * vector[92] +matrix[93][213] * vector[93] +matrix[94][213] * vector[94] +matrix[95][213] * vector[95] +matrix[96][213] * vector[96] +matrix[97][213] * vector[97] +matrix[98][213] * vector[98] +matrix[99][213] * vector[99] +b[213];
assign result[214] = matrix[0][214] * vector[0] +matrix[1][214] * vector[1] +matrix[2][214] * vector[2] +matrix[3][214] * vector[3] +matrix[4][214] * vector[4] +matrix[5][214] * vector[5] +matrix[6][214] * vector[6] +matrix[7][214] * vector[7] +matrix[8][214] * vector[8] +matrix[9][214] * vector[9] +matrix[10][214] * vector[10] +matrix[11][214] * vector[11] +matrix[12][214] * vector[12] +matrix[13][214] * vector[13] +matrix[14][214] * vector[14] +matrix[15][214] * vector[15] +matrix[16][214] * vector[16] +matrix[17][214] * vector[17] +matrix[18][214] * vector[18] +matrix[19][214] * vector[19] +matrix[20][214] * vector[20] +matrix[21][214] * vector[21] +matrix[22][214] * vector[22] +matrix[23][214] * vector[23] +matrix[24][214] * vector[24] +matrix[25][214] * vector[25] +matrix[26][214] * vector[26] +matrix[27][214] * vector[27] +matrix[28][214] * vector[28] +matrix[29][214] * vector[29] +matrix[30][214] * vector[30] +matrix[31][214] * vector[31] +matrix[32][214] * vector[32] +matrix[33][214] * vector[33] +matrix[34][214] * vector[34] +matrix[35][214] * vector[35] +matrix[36][214] * vector[36] +matrix[37][214] * vector[37] +matrix[38][214] * vector[38] +matrix[39][214] * vector[39] +matrix[40][214] * vector[40] +matrix[41][214] * vector[41] +matrix[42][214] * vector[42] +matrix[43][214] * vector[43] +matrix[44][214] * vector[44] +matrix[45][214] * vector[45] +matrix[46][214] * vector[46] +matrix[47][214] * vector[47] +matrix[48][214] * vector[48] +matrix[49][214] * vector[49] +matrix[50][214] * vector[50] +matrix[51][214] * vector[51] +matrix[52][214] * vector[52] +matrix[53][214] * vector[53] +matrix[54][214] * vector[54] +matrix[55][214] * vector[55] +matrix[56][214] * vector[56] +matrix[57][214] * vector[57] +matrix[58][214] * vector[58] +matrix[59][214] * vector[59] +matrix[60][214] * vector[60] +matrix[61][214] * vector[61] +matrix[62][214] * vector[62] +matrix[63][214] * vector[63] +matrix[64][214] * vector[64] +matrix[65][214] * vector[65] +matrix[66][214] * vector[66] +matrix[67][214] * vector[67] +matrix[68][214] * vector[68] +matrix[69][214] * vector[69] +matrix[70][214] * vector[70] +matrix[71][214] * vector[71] +matrix[72][214] * vector[72] +matrix[73][214] * vector[73] +matrix[74][214] * vector[74] +matrix[75][214] * vector[75] +matrix[76][214] * vector[76] +matrix[77][214] * vector[77] +matrix[78][214] * vector[78] +matrix[79][214] * vector[79] +matrix[80][214] * vector[80] +matrix[81][214] * vector[81] +matrix[82][214] * vector[82] +matrix[83][214] * vector[83] +matrix[84][214] * vector[84] +matrix[85][214] * vector[85] +matrix[86][214] * vector[86] +matrix[87][214] * vector[87] +matrix[88][214] * vector[88] +matrix[89][214] * vector[89] +matrix[90][214] * vector[90] +matrix[91][214] * vector[91] +matrix[92][214] * vector[92] +matrix[93][214] * vector[93] +matrix[94][214] * vector[94] +matrix[95][214] * vector[95] +matrix[96][214] * vector[96] +matrix[97][214] * vector[97] +matrix[98][214] * vector[98] +matrix[99][214] * vector[99] +b[214];
assign result[215] = matrix[0][215] * vector[0] +matrix[1][215] * vector[1] +matrix[2][215] * vector[2] +matrix[3][215] * vector[3] +matrix[4][215] * vector[4] +matrix[5][215] * vector[5] +matrix[6][215] * vector[6] +matrix[7][215] * vector[7] +matrix[8][215] * vector[8] +matrix[9][215] * vector[9] +matrix[10][215] * vector[10] +matrix[11][215] * vector[11] +matrix[12][215] * vector[12] +matrix[13][215] * vector[13] +matrix[14][215] * vector[14] +matrix[15][215] * vector[15] +matrix[16][215] * vector[16] +matrix[17][215] * vector[17] +matrix[18][215] * vector[18] +matrix[19][215] * vector[19] +matrix[20][215] * vector[20] +matrix[21][215] * vector[21] +matrix[22][215] * vector[22] +matrix[23][215] * vector[23] +matrix[24][215] * vector[24] +matrix[25][215] * vector[25] +matrix[26][215] * vector[26] +matrix[27][215] * vector[27] +matrix[28][215] * vector[28] +matrix[29][215] * vector[29] +matrix[30][215] * vector[30] +matrix[31][215] * vector[31] +matrix[32][215] * vector[32] +matrix[33][215] * vector[33] +matrix[34][215] * vector[34] +matrix[35][215] * vector[35] +matrix[36][215] * vector[36] +matrix[37][215] * vector[37] +matrix[38][215] * vector[38] +matrix[39][215] * vector[39] +matrix[40][215] * vector[40] +matrix[41][215] * vector[41] +matrix[42][215] * vector[42] +matrix[43][215] * vector[43] +matrix[44][215] * vector[44] +matrix[45][215] * vector[45] +matrix[46][215] * vector[46] +matrix[47][215] * vector[47] +matrix[48][215] * vector[48] +matrix[49][215] * vector[49] +matrix[50][215] * vector[50] +matrix[51][215] * vector[51] +matrix[52][215] * vector[52] +matrix[53][215] * vector[53] +matrix[54][215] * vector[54] +matrix[55][215] * vector[55] +matrix[56][215] * vector[56] +matrix[57][215] * vector[57] +matrix[58][215] * vector[58] +matrix[59][215] * vector[59] +matrix[60][215] * vector[60] +matrix[61][215] * vector[61] +matrix[62][215] * vector[62] +matrix[63][215] * vector[63] +matrix[64][215] * vector[64] +matrix[65][215] * vector[65] +matrix[66][215] * vector[66] +matrix[67][215] * vector[67] +matrix[68][215] * vector[68] +matrix[69][215] * vector[69] +matrix[70][215] * vector[70] +matrix[71][215] * vector[71] +matrix[72][215] * vector[72] +matrix[73][215] * vector[73] +matrix[74][215] * vector[74] +matrix[75][215] * vector[75] +matrix[76][215] * vector[76] +matrix[77][215] * vector[77] +matrix[78][215] * vector[78] +matrix[79][215] * vector[79] +matrix[80][215] * vector[80] +matrix[81][215] * vector[81] +matrix[82][215] * vector[82] +matrix[83][215] * vector[83] +matrix[84][215] * vector[84] +matrix[85][215] * vector[85] +matrix[86][215] * vector[86] +matrix[87][215] * vector[87] +matrix[88][215] * vector[88] +matrix[89][215] * vector[89] +matrix[90][215] * vector[90] +matrix[91][215] * vector[91] +matrix[92][215] * vector[92] +matrix[93][215] * vector[93] +matrix[94][215] * vector[94] +matrix[95][215] * vector[95] +matrix[96][215] * vector[96] +matrix[97][215] * vector[97] +matrix[98][215] * vector[98] +matrix[99][215] * vector[99] +b[215];
assign result[216] = matrix[0][216] * vector[0] +matrix[1][216] * vector[1] +matrix[2][216] * vector[2] +matrix[3][216] * vector[3] +matrix[4][216] * vector[4] +matrix[5][216] * vector[5] +matrix[6][216] * vector[6] +matrix[7][216] * vector[7] +matrix[8][216] * vector[8] +matrix[9][216] * vector[9] +matrix[10][216] * vector[10] +matrix[11][216] * vector[11] +matrix[12][216] * vector[12] +matrix[13][216] * vector[13] +matrix[14][216] * vector[14] +matrix[15][216] * vector[15] +matrix[16][216] * vector[16] +matrix[17][216] * vector[17] +matrix[18][216] * vector[18] +matrix[19][216] * vector[19] +matrix[20][216] * vector[20] +matrix[21][216] * vector[21] +matrix[22][216] * vector[22] +matrix[23][216] * vector[23] +matrix[24][216] * vector[24] +matrix[25][216] * vector[25] +matrix[26][216] * vector[26] +matrix[27][216] * vector[27] +matrix[28][216] * vector[28] +matrix[29][216] * vector[29] +matrix[30][216] * vector[30] +matrix[31][216] * vector[31] +matrix[32][216] * vector[32] +matrix[33][216] * vector[33] +matrix[34][216] * vector[34] +matrix[35][216] * vector[35] +matrix[36][216] * vector[36] +matrix[37][216] * vector[37] +matrix[38][216] * vector[38] +matrix[39][216] * vector[39] +matrix[40][216] * vector[40] +matrix[41][216] * vector[41] +matrix[42][216] * vector[42] +matrix[43][216] * vector[43] +matrix[44][216] * vector[44] +matrix[45][216] * vector[45] +matrix[46][216] * vector[46] +matrix[47][216] * vector[47] +matrix[48][216] * vector[48] +matrix[49][216] * vector[49] +matrix[50][216] * vector[50] +matrix[51][216] * vector[51] +matrix[52][216] * vector[52] +matrix[53][216] * vector[53] +matrix[54][216] * vector[54] +matrix[55][216] * vector[55] +matrix[56][216] * vector[56] +matrix[57][216] * vector[57] +matrix[58][216] * vector[58] +matrix[59][216] * vector[59] +matrix[60][216] * vector[60] +matrix[61][216] * vector[61] +matrix[62][216] * vector[62] +matrix[63][216] * vector[63] +matrix[64][216] * vector[64] +matrix[65][216] * vector[65] +matrix[66][216] * vector[66] +matrix[67][216] * vector[67] +matrix[68][216] * vector[68] +matrix[69][216] * vector[69] +matrix[70][216] * vector[70] +matrix[71][216] * vector[71] +matrix[72][216] * vector[72] +matrix[73][216] * vector[73] +matrix[74][216] * vector[74] +matrix[75][216] * vector[75] +matrix[76][216] * vector[76] +matrix[77][216] * vector[77] +matrix[78][216] * vector[78] +matrix[79][216] * vector[79] +matrix[80][216] * vector[80] +matrix[81][216] * vector[81] +matrix[82][216] * vector[82] +matrix[83][216] * vector[83] +matrix[84][216] * vector[84] +matrix[85][216] * vector[85] +matrix[86][216] * vector[86] +matrix[87][216] * vector[87] +matrix[88][216] * vector[88] +matrix[89][216] * vector[89] +matrix[90][216] * vector[90] +matrix[91][216] * vector[91] +matrix[92][216] * vector[92] +matrix[93][216] * vector[93] +matrix[94][216] * vector[94] +matrix[95][216] * vector[95] +matrix[96][216] * vector[96] +matrix[97][216] * vector[97] +matrix[98][216] * vector[98] +matrix[99][216] * vector[99] +b[216];
assign result[217] = matrix[0][217] * vector[0] +matrix[1][217] * vector[1] +matrix[2][217] * vector[2] +matrix[3][217] * vector[3] +matrix[4][217] * vector[4] +matrix[5][217] * vector[5] +matrix[6][217] * vector[6] +matrix[7][217] * vector[7] +matrix[8][217] * vector[8] +matrix[9][217] * vector[9] +matrix[10][217] * vector[10] +matrix[11][217] * vector[11] +matrix[12][217] * vector[12] +matrix[13][217] * vector[13] +matrix[14][217] * vector[14] +matrix[15][217] * vector[15] +matrix[16][217] * vector[16] +matrix[17][217] * vector[17] +matrix[18][217] * vector[18] +matrix[19][217] * vector[19] +matrix[20][217] * vector[20] +matrix[21][217] * vector[21] +matrix[22][217] * vector[22] +matrix[23][217] * vector[23] +matrix[24][217] * vector[24] +matrix[25][217] * vector[25] +matrix[26][217] * vector[26] +matrix[27][217] * vector[27] +matrix[28][217] * vector[28] +matrix[29][217] * vector[29] +matrix[30][217] * vector[30] +matrix[31][217] * vector[31] +matrix[32][217] * vector[32] +matrix[33][217] * vector[33] +matrix[34][217] * vector[34] +matrix[35][217] * vector[35] +matrix[36][217] * vector[36] +matrix[37][217] * vector[37] +matrix[38][217] * vector[38] +matrix[39][217] * vector[39] +matrix[40][217] * vector[40] +matrix[41][217] * vector[41] +matrix[42][217] * vector[42] +matrix[43][217] * vector[43] +matrix[44][217] * vector[44] +matrix[45][217] * vector[45] +matrix[46][217] * vector[46] +matrix[47][217] * vector[47] +matrix[48][217] * vector[48] +matrix[49][217] * vector[49] +matrix[50][217] * vector[50] +matrix[51][217] * vector[51] +matrix[52][217] * vector[52] +matrix[53][217] * vector[53] +matrix[54][217] * vector[54] +matrix[55][217] * vector[55] +matrix[56][217] * vector[56] +matrix[57][217] * vector[57] +matrix[58][217] * vector[58] +matrix[59][217] * vector[59] +matrix[60][217] * vector[60] +matrix[61][217] * vector[61] +matrix[62][217] * vector[62] +matrix[63][217] * vector[63] +matrix[64][217] * vector[64] +matrix[65][217] * vector[65] +matrix[66][217] * vector[66] +matrix[67][217] * vector[67] +matrix[68][217] * vector[68] +matrix[69][217] * vector[69] +matrix[70][217] * vector[70] +matrix[71][217] * vector[71] +matrix[72][217] * vector[72] +matrix[73][217] * vector[73] +matrix[74][217] * vector[74] +matrix[75][217] * vector[75] +matrix[76][217] * vector[76] +matrix[77][217] * vector[77] +matrix[78][217] * vector[78] +matrix[79][217] * vector[79] +matrix[80][217] * vector[80] +matrix[81][217] * vector[81] +matrix[82][217] * vector[82] +matrix[83][217] * vector[83] +matrix[84][217] * vector[84] +matrix[85][217] * vector[85] +matrix[86][217] * vector[86] +matrix[87][217] * vector[87] +matrix[88][217] * vector[88] +matrix[89][217] * vector[89] +matrix[90][217] * vector[90] +matrix[91][217] * vector[91] +matrix[92][217] * vector[92] +matrix[93][217] * vector[93] +matrix[94][217] * vector[94] +matrix[95][217] * vector[95] +matrix[96][217] * vector[96] +matrix[97][217] * vector[97] +matrix[98][217] * vector[98] +matrix[99][217] * vector[99] +b[217];
assign result[218] = matrix[0][218] * vector[0] +matrix[1][218] * vector[1] +matrix[2][218] * vector[2] +matrix[3][218] * vector[3] +matrix[4][218] * vector[4] +matrix[5][218] * vector[5] +matrix[6][218] * vector[6] +matrix[7][218] * vector[7] +matrix[8][218] * vector[8] +matrix[9][218] * vector[9] +matrix[10][218] * vector[10] +matrix[11][218] * vector[11] +matrix[12][218] * vector[12] +matrix[13][218] * vector[13] +matrix[14][218] * vector[14] +matrix[15][218] * vector[15] +matrix[16][218] * vector[16] +matrix[17][218] * vector[17] +matrix[18][218] * vector[18] +matrix[19][218] * vector[19] +matrix[20][218] * vector[20] +matrix[21][218] * vector[21] +matrix[22][218] * vector[22] +matrix[23][218] * vector[23] +matrix[24][218] * vector[24] +matrix[25][218] * vector[25] +matrix[26][218] * vector[26] +matrix[27][218] * vector[27] +matrix[28][218] * vector[28] +matrix[29][218] * vector[29] +matrix[30][218] * vector[30] +matrix[31][218] * vector[31] +matrix[32][218] * vector[32] +matrix[33][218] * vector[33] +matrix[34][218] * vector[34] +matrix[35][218] * vector[35] +matrix[36][218] * vector[36] +matrix[37][218] * vector[37] +matrix[38][218] * vector[38] +matrix[39][218] * vector[39] +matrix[40][218] * vector[40] +matrix[41][218] * vector[41] +matrix[42][218] * vector[42] +matrix[43][218] * vector[43] +matrix[44][218] * vector[44] +matrix[45][218] * vector[45] +matrix[46][218] * vector[46] +matrix[47][218] * vector[47] +matrix[48][218] * vector[48] +matrix[49][218] * vector[49] +matrix[50][218] * vector[50] +matrix[51][218] * vector[51] +matrix[52][218] * vector[52] +matrix[53][218] * vector[53] +matrix[54][218] * vector[54] +matrix[55][218] * vector[55] +matrix[56][218] * vector[56] +matrix[57][218] * vector[57] +matrix[58][218] * vector[58] +matrix[59][218] * vector[59] +matrix[60][218] * vector[60] +matrix[61][218] * vector[61] +matrix[62][218] * vector[62] +matrix[63][218] * vector[63] +matrix[64][218] * vector[64] +matrix[65][218] * vector[65] +matrix[66][218] * vector[66] +matrix[67][218] * vector[67] +matrix[68][218] * vector[68] +matrix[69][218] * vector[69] +matrix[70][218] * vector[70] +matrix[71][218] * vector[71] +matrix[72][218] * vector[72] +matrix[73][218] * vector[73] +matrix[74][218] * vector[74] +matrix[75][218] * vector[75] +matrix[76][218] * vector[76] +matrix[77][218] * vector[77] +matrix[78][218] * vector[78] +matrix[79][218] * vector[79] +matrix[80][218] * vector[80] +matrix[81][218] * vector[81] +matrix[82][218] * vector[82] +matrix[83][218] * vector[83] +matrix[84][218] * vector[84] +matrix[85][218] * vector[85] +matrix[86][218] * vector[86] +matrix[87][218] * vector[87] +matrix[88][218] * vector[88] +matrix[89][218] * vector[89] +matrix[90][218] * vector[90] +matrix[91][218] * vector[91] +matrix[92][218] * vector[92] +matrix[93][218] * vector[93] +matrix[94][218] * vector[94] +matrix[95][218] * vector[95] +matrix[96][218] * vector[96] +matrix[97][218] * vector[97] +matrix[98][218] * vector[98] +matrix[99][218] * vector[99] +b[218];
assign result[219] = matrix[0][219] * vector[0] +matrix[1][219] * vector[1] +matrix[2][219] * vector[2] +matrix[3][219] * vector[3] +matrix[4][219] * vector[4] +matrix[5][219] * vector[5] +matrix[6][219] * vector[6] +matrix[7][219] * vector[7] +matrix[8][219] * vector[8] +matrix[9][219] * vector[9] +matrix[10][219] * vector[10] +matrix[11][219] * vector[11] +matrix[12][219] * vector[12] +matrix[13][219] * vector[13] +matrix[14][219] * vector[14] +matrix[15][219] * vector[15] +matrix[16][219] * vector[16] +matrix[17][219] * vector[17] +matrix[18][219] * vector[18] +matrix[19][219] * vector[19] +matrix[20][219] * vector[20] +matrix[21][219] * vector[21] +matrix[22][219] * vector[22] +matrix[23][219] * vector[23] +matrix[24][219] * vector[24] +matrix[25][219] * vector[25] +matrix[26][219] * vector[26] +matrix[27][219] * vector[27] +matrix[28][219] * vector[28] +matrix[29][219] * vector[29] +matrix[30][219] * vector[30] +matrix[31][219] * vector[31] +matrix[32][219] * vector[32] +matrix[33][219] * vector[33] +matrix[34][219] * vector[34] +matrix[35][219] * vector[35] +matrix[36][219] * vector[36] +matrix[37][219] * vector[37] +matrix[38][219] * vector[38] +matrix[39][219] * vector[39] +matrix[40][219] * vector[40] +matrix[41][219] * vector[41] +matrix[42][219] * vector[42] +matrix[43][219] * vector[43] +matrix[44][219] * vector[44] +matrix[45][219] * vector[45] +matrix[46][219] * vector[46] +matrix[47][219] * vector[47] +matrix[48][219] * vector[48] +matrix[49][219] * vector[49] +matrix[50][219] * vector[50] +matrix[51][219] * vector[51] +matrix[52][219] * vector[52] +matrix[53][219] * vector[53] +matrix[54][219] * vector[54] +matrix[55][219] * vector[55] +matrix[56][219] * vector[56] +matrix[57][219] * vector[57] +matrix[58][219] * vector[58] +matrix[59][219] * vector[59] +matrix[60][219] * vector[60] +matrix[61][219] * vector[61] +matrix[62][219] * vector[62] +matrix[63][219] * vector[63] +matrix[64][219] * vector[64] +matrix[65][219] * vector[65] +matrix[66][219] * vector[66] +matrix[67][219] * vector[67] +matrix[68][219] * vector[68] +matrix[69][219] * vector[69] +matrix[70][219] * vector[70] +matrix[71][219] * vector[71] +matrix[72][219] * vector[72] +matrix[73][219] * vector[73] +matrix[74][219] * vector[74] +matrix[75][219] * vector[75] +matrix[76][219] * vector[76] +matrix[77][219] * vector[77] +matrix[78][219] * vector[78] +matrix[79][219] * vector[79] +matrix[80][219] * vector[80] +matrix[81][219] * vector[81] +matrix[82][219] * vector[82] +matrix[83][219] * vector[83] +matrix[84][219] * vector[84] +matrix[85][219] * vector[85] +matrix[86][219] * vector[86] +matrix[87][219] * vector[87] +matrix[88][219] * vector[88] +matrix[89][219] * vector[89] +matrix[90][219] * vector[90] +matrix[91][219] * vector[91] +matrix[92][219] * vector[92] +matrix[93][219] * vector[93] +matrix[94][219] * vector[94] +matrix[95][219] * vector[95] +matrix[96][219] * vector[96] +matrix[97][219] * vector[97] +matrix[98][219] * vector[98] +matrix[99][219] * vector[99] +b[219];
assign result[220] = matrix[0][220] * vector[0] +matrix[1][220] * vector[1] +matrix[2][220] * vector[2] +matrix[3][220] * vector[3] +matrix[4][220] * vector[4] +matrix[5][220] * vector[5] +matrix[6][220] * vector[6] +matrix[7][220] * vector[7] +matrix[8][220] * vector[8] +matrix[9][220] * vector[9] +matrix[10][220] * vector[10] +matrix[11][220] * vector[11] +matrix[12][220] * vector[12] +matrix[13][220] * vector[13] +matrix[14][220] * vector[14] +matrix[15][220] * vector[15] +matrix[16][220] * vector[16] +matrix[17][220] * vector[17] +matrix[18][220] * vector[18] +matrix[19][220] * vector[19] +matrix[20][220] * vector[20] +matrix[21][220] * vector[21] +matrix[22][220] * vector[22] +matrix[23][220] * vector[23] +matrix[24][220] * vector[24] +matrix[25][220] * vector[25] +matrix[26][220] * vector[26] +matrix[27][220] * vector[27] +matrix[28][220] * vector[28] +matrix[29][220] * vector[29] +matrix[30][220] * vector[30] +matrix[31][220] * vector[31] +matrix[32][220] * vector[32] +matrix[33][220] * vector[33] +matrix[34][220] * vector[34] +matrix[35][220] * vector[35] +matrix[36][220] * vector[36] +matrix[37][220] * vector[37] +matrix[38][220] * vector[38] +matrix[39][220] * vector[39] +matrix[40][220] * vector[40] +matrix[41][220] * vector[41] +matrix[42][220] * vector[42] +matrix[43][220] * vector[43] +matrix[44][220] * vector[44] +matrix[45][220] * vector[45] +matrix[46][220] * vector[46] +matrix[47][220] * vector[47] +matrix[48][220] * vector[48] +matrix[49][220] * vector[49] +matrix[50][220] * vector[50] +matrix[51][220] * vector[51] +matrix[52][220] * vector[52] +matrix[53][220] * vector[53] +matrix[54][220] * vector[54] +matrix[55][220] * vector[55] +matrix[56][220] * vector[56] +matrix[57][220] * vector[57] +matrix[58][220] * vector[58] +matrix[59][220] * vector[59] +matrix[60][220] * vector[60] +matrix[61][220] * vector[61] +matrix[62][220] * vector[62] +matrix[63][220] * vector[63] +matrix[64][220] * vector[64] +matrix[65][220] * vector[65] +matrix[66][220] * vector[66] +matrix[67][220] * vector[67] +matrix[68][220] * vector[68] +matrix[69][220] * vector[69] +matrix[70][220] * vector[70] +matrix[71][220] * vector[71] +matrix[72][220] * vector[72] +matrix[73][220] * vector[73] +matrix[74][220] * vector[74] +matrix[75][220] * vector[75] +matrix[76][220] * vector[76] +matrix[77][220] * vector[77] +matrix[78][220] * vector[78] +matrix[79][220] * vector[79] +matrix[80][220] * vector[80] +matrix[81][220] * vector[81] +matrix[82][220] * vector[82] +matrix[83][220] * vector[83] +matrix[84][220] * vector[84] +matrix[85][220] * vector[85] +matrix[86][220] * vector[86] +matrix[87][220] * vector[87] +matrix[88][220] * vector[88] +matrix[89][220] * vector[89] +matrix[90][220] * vector[90] +matrix[91][220] * vector[91] +matrix[92][220] * vector[92] +matrix[93][220] * vector[93] +matrix[94][220] * vector[94] +matrix[95][220] * vector[95] +matrix[96][220] * vector[96] +matrix[97][220] * vector[97] +matrix[98][220] * vector[98] +matrix[99][220] * vector[99] +b[220];
assign result[221] = matrix[0][221] * vector[0] +matrix[1][221] * vector[1] +matrix[2][221] * vector[2] +matrix[3][221] * vector[3] +matrix[4][221] * vector[4] +matrix[5][221] * vector[5] +matrix[6][221] * vector[6] +matrix[7][221] * vector[7] +matrix[8][221] * vector[8] +matrix[9][221] * vector[9] +matrix[10][221] * vector[10] +matrix[11][221] * vector[11] +matrix[12][221] * vector[12] +matrix[13][221] * vector[13] +matrix[14][221] * vector[14] +matrix[15][221] * vector[15] +matrix[16][221] * vector[16] +matrix[17][221] * vector[17] +matrix[18][221] * vector[18] +matrix[19][221] * vector[19] +matrix[20][221] * vector[20] +matrix[21][221] * vector[21] +matrix[22][221] * vector[22] +matrix[23][221] * vector[23] +matrix[24][221] * vector[24] +matrix[25][221] * vector[25] +matrix[26][221] * vector[26] +matrix[27][221] * vector[27] +matrix[28][221] * vector[28] +matrix[29][221] * vector[29] +matrix[30][221] * vector[30] +matrix[31][221] * vector[31] +matrix[32][221] * vector[32] +matrix[33][221] * vector[33] +matrix[34][221] * vector[34] +matrix[35][221] * vector[35] +matrix[36][221] * vector[36] +matrix[37][221] * vector[37] +matrix[38][221] * vector[38] +matrix[39][221] * vector[39] +matrix[40][221] * vector[40] +matrix[41][221] * vector[41] +matrix[42][221] * vector[42] +matrix[43][221] * vector[43] +matrix[44][221] * vector[44] +matrix[45][221] * vector[45] +matrix[46][221] * vector[46] +matrix[47][221] * vector[47] +matrix[48][221] * vector[48] +matrix[49][221] * vector[49] +matrix[50][221] * vector[50] +matrix[51][221] * vector[51] +matrix[52][221] * vector[52] +matrix[53][221] * vector[53] +matrix[54][221] * vector[54] +matrix[55][221] * vector[55] +matrix[56][221] * vector[56] +matrix[57][221] * vector[57] +matrix[58][221] * vector[58] +matrix[59][221] * vector[59] +matrix[60][221] * vector[60] +matrix[61][221] * vector[61] +matrix[62][221] * vector[62] +matrix[63][221] * vector[63] +matrix[64][221] * vector[64] +matrix[65][221] * vector[65] +matrix[66][221] * vector[66] +matrix[67][221] * vector[67] +matrix[68][221] * vector[68] +matrix[69][221] * vector[69] +matrix[70][221] * vector[70] +matrix[71][221] * vector[71] +matrix[72][221] * vector[72] +matrix[73][221] * vector[73] +matrix[74][221] * vector[74] +matrix[75][221] * vector[75] +matrix[76][221] * vector[76] +matrix[77][221] * vector[77] +matrix[78][221] * vector[78] +matrix[79][221] * vector[79] +matrix[80][221] * vector[80] +matrix[81][221] * vector[81] +matrix[82][221] * vector[82] +matrix[83][221] * vector[83] +matrix[84][221] * vector[84] +matrix[85][221] * vector[85] +matrix[86][221] * vector[86] +matrix[87][221] * vector[87] +matrix[88][221] * vector[88] +matrix[89][221] * vector[89] +matrix[90][221] * vector[90] +matrix[91][221] * vector[91] +matrix[92][221] * vector[92] +matrix[93][221] * vector[93] +matrix[94][221] * vector[94] +matrix[95][221] * vector[95] +matrix[96][221] * vector[96] +matrix[97][221] * vector[97] +matrix[98][221] * vector[98] +matrix[99][221] * vector[99] +b[221];
assign result[222] = matrix[0][222] * vector[0] +matrix[1][222] * vector[1] +matrix[2][222] * vector[2] +matrix[3][222] * vector[3] +matrix[4][222] * vector[4] +matrix[5][222] * vector[5] +matrix[6][222] * vector[6] +matrix[7][222] * vector[7] +matrix[8][222] * vector[8] +matrix[9][222] * vector[9] +matrix[10][222] * vector[10] +matrix[11][222] * vector[11] +matrix[12][222] * vector[12] +matrix[13][222] * vector[13] +matrix[14][222] * vector[14] +matrix[15][222] * vector[15] +matrix[16][222] * vector[16] +matrix[17][222] * vector[17] +matrix[18][222] * vector[18] +matrix[19][222] * vector[19] +matrix[20][222] * vector[20] +matrix[21][222] * vector[21] +matrix[22][222] * vector[22] +matrix[23][222] * vector[23] +matrix[24][222] * vector[24] +matrix[25][222] * vector[25] +matrix[26][222] * vector[26] +matrix[27][222] * vector[27] +matrix[28][222] * vector[28] +matrix[29][222] * vector[29] +matrix[30][222] * vector[30] +matrix[31][222] * vector[31] +matrix[32][222] * vector[32] +matrix[33][222] * vector[33] +matrix[34][222] * vector[34] +matrix[35][222] * vector[35] +matrix[36][222] * vector[36] +matrix[37][222] * vector[37] +matrix[38][222] * vector[38] +matrix[39][222] * vector[39] +matrix[40][222] * vector[40] +matrix[41][222] * vector[41] +matrix[42][222] * vector[42] +matrix[43][222] * vector[43] +matrix[44][222] * vector[44] +matrix[45][222] * vector[45] +matrix[46][222] * vector[46] +matrix[47][222] * vector[47] +matrix[48][222] * vector[48] +matrix[49][222] * vector[49] +matrix[50][222] * vector[50] +matrix[51][222] * vector[51] +matrix[52][222] * vector[52] +matrix[53][222] * vector[53] +matrix[54][222] * vector[54] +matrix[55][222] * vector[55] +matrix[56][222] * vector[56] +matrix[57][222] * vector[57] +matrix[58][222] * vector[58] +matrix[59][222] * vector[59] +matrix[60][222] * vector[60] +matrix[61][222] * vector[61] +matrix[62][222] * vector[62] +matrix[63][222] * vector[63] +matrix[64][222] * vector[64] +matrix[65][222] * vector[65] +matrix[66][222] * vector[66] +matrix[67][222] * vector[67] +matrix[68][222] * vector[68] +matrix[69][222] * vector[69] +matrix[70][222] * vector[70] +matrix[71][222] * vector[71] +matrix[72][222] * vector[72] +matrix[73][222] * vector[73] +matrix[74][222] * vector[74] +matrix[75][222] * vector[75] +matrix[76][222] * vector[76] +matrix[77][222] * vector[77] +matrix[78][222] * vector[78] +matrix[79][222] * vector[79] +matrix[80][222] * vector[80] +matrix[81][222] * vector[81] +matrix[82][222] * vector[82] +matrix[83][222] * vector[83] +matrix[84][222] * vector[84] +matrix[85][222] * vector[85] +matrix[86][222] * vector[86] +matrix[87][222] * vector[87] +matrix[88][222] * vector[88] +matrix[89][222] * vector[89] +matrix[90][222] * vector[90] +matrix[91][222] * vector[91] +matrix[92][222] * vector[92] +matrix[93][222] * vector[93] +matrix[94][222] * vector[94] +matrix[95][222] * vector[95] +matrix[96][222] * vector[96] +matrix[97][222] * vector[97] +matrix[98][222] * vector[98] +matrix[99][222] * vector[99] +b[222];
assign result[223] = matrix[0][223] * vector[0] +matrix[1][223] * vector[1] +matrix[2][223] * vector[2] +matrix[3][223] * vector[3] +matrix[4][223] * vector[4] +matrix[5][223] * vector[5] +matrix[6][223] * vector[6] +matrix[7][223] * vector[7] +matrix[8][223] * vector[8] +matrix[9][223] * vector[9] +matrix[10][223] * vector[10] +matrix[11][223] * vector[11] +matrix[12][223] * vector[12] +matrix[13][223] * vector[13] +matrix[14][223] * vector[14] +matrix[15][223] * vector[15] +matrix[16][223] * vector[16] +matrix[17][223] * vector[17] +matrix[18][223] * vector[18] +matrix[19][223] * vector[19] +matrix[20][223] * vector[20] +matrix[21][223] * vector[21] +matrix[22][223] * vector[22] +matrix[23][223] * vector[23] +matrix[24][223] * vector[24] +matrix[25][223] * vector[25] +matrix[26][223] * vector[26] +matrix[27][223] * vector[27] +matrix[28][223] * vector[28] +matrix[29][223] * vector[29] +matrix[30][223] * vector[30] +matrix[31][223] * vector[31] +matrix[32][223] * vector[32] +matrix[33][223] * vector[33] +matrix[34][223] * vector[34] +matrix[35][223] * vector[35] +matrix[36][223] * vector[36] +matrix[37][223] * vector[37] +matrix[38][223] * vector[38] +matrix[39][223] * vector[39] +matrix[40][223] * vector[40] +matrix[41][223] * vector[41] +matrix[42][223] * vector[42] +matrix[43][223] * vector[43] +matrix[44][223] * vector[44] +matrix[45][223] * vector[45] +matrix[46][223] * vector[46] +matrix[47][223] * vector[47] +matrix[48][223] * vector[48] +matrix[49][223] * vector[49] +matrix[50][223] * vector[50] +matrix[51][223] * vector[51] +matrix[52][223] * vector[52] +matrix[53][223] * vector[53] +matrix[54][223] * vector[54] +matrix[55][223] * vector[55] +matrix[56][223] * vector[56] +matrix[57][223] * vector[57] +matrix[58][223] * vector[58] +matrix[59][223] * vector[59] +matrix[60][223] * vector[60] +matrix[61][223] * vector[61] +matrix[62][223] * vector[62] +matrix[63][223] * vector[63] +matrix[64][223] * vector[64] +matrix[65][223] * vector[65] +matrix[66][223] * vector[66] +matrix[67][223] * vector[67] +matrix[68][223] * vector[68] +matrix[69][223] * vector[69] +matrix[70][223] * vector[70] +matrix[71][223] * vector[71] +matrix[72][223] * vector[72] +matrix[73][223] * vector[73] +matrix[74][223] * vector[74] +matrix[75][223] * vector[75] +matrix[76][223] * vector[76] +matrix[77][223] * vector[77] +matrix[78][223] * vector[78] +matrix[79][223] * vector[79] +matrix[80][223] * vector[80] +matrix[81][223] * vector[81] +matrix[82][223] * vector[82] +matrix[83][223] * vector[83] +matrix[84][223] * vector[84] +matrix[85][223] * vector[85] +matrix[86][223] * vector[86] +matrix[87][223] * vector[87] +matrix[88][223] * vector[88] +matrix[89][223] * vector[89] +matrix[90][223] * vector[90] +matrix[91][223] * vector[91] +matrix[92][223] * vector[92] +matrix[93][223] * vector[93] +matrix[94][223] * vector[94] +matrix[95][223] * vector[95] +matrix[96][223] * vector[96] +matrix[97][223] * vector[97] +matrix[98][223] * vector[98] +matrix[99][223] * vector[99] +b[223];
assign result[224] = matrix[0][224] * vector[0] +matrix[1][224] * vector[1] +matrix[2][224] * vector[2] +matrix[3][224] * vector[3] +matrix[4][224] * vector[4] +matrix[5][224] * vector[5] +matrix[6][224] * vector[6] +matrix[7][224] * vector[7] +matrix[8][224] * vector[8] +matrix[9][224] * vector[9] +matrix[10][224] * vector[10] +matrix[11][224] * vector[11] +matrix[12][224] * vector[12] +matrix[13][224] * vector[13] +matrix[14][224] * vector[14] +matrix[15][224] * vector[15] +matrix[16][224] * vector[16] +matrix[17][224] * vector[17] +matrix[18][224] * vector[18] +matrix[19][224] * vector[19] +matrix[20][224] * vector[20] +matrix[21][224] * vector[21] +matrix[22][224] * vector[22] +matrix[23][224] * vector[23] +matrix[24][224] * vector[24] +matrix[25][224] * vector[25] +matrix[26][224] * vector[26] +matrix[27][224] * vector[27] +matrix[28][224] * vector[28] +matrix[29][224] * vector[29] +matrix[30][224] * vector[30] +matrix[31][224] * vector[31] +matrix[32][224] * vector[32] +matrix[33][224] * vector[33] +matrix[34][224] * vector[34] +matrix[35][224] * vector[35] +matrix[36][224] * vector[36] +matrix[37][224] * vector[37] +matrix[38][224] * vector[38] +matrix[39][224] * vector[39] +matrix[40][224] * vector[40] +matrix[41][224] * vector[41] +matrix[42][224] * vector[42] +matrix[43][224] * vector[43] +matrix[44][224] * vector[44] +matrix[45][224] * vector[45] +matrix[46][224] * vector[46] +matrix[47][224] * vector[47] +matrix[48][224] * vector[48] +matrix[49][224] * vector[49] +matrix[50][224] * vector[50] +matrix[51][224] * vector[51] +matrix[52][224] * vector[52] +matrix[53][224] * vector[53] +matrix[54][224] * vector[54] +matrix[55][224] * vector[55] +matrix[56][224] * vector[56] +matrix[57][224] * vector[57] +matrix[58][224] * vector[58] +matrix[59][224] * vector[59] +matrix[60][224] * vector[60] +matrix[61][224] * vector[61] +matrix[62][224] * vector[62] +matrix[63][224] * vector[63] +matrix[64][224] * vector[64] +matrix[65][224] * vector[65] +matrix[66][224] * vector[66] +matrix[67][224] * vector[67] +matrix[68][224] * vector[68] +matrix[69][224] * vector[69] +matrix[70][224] * vector[70] +matrix[71][224] * vector[71] +matrix[72][224] * vector[72] +matrix[73][224] * vector[73] +matrix[74][224] * vector[74] +matrix[75][224] * vector[75] +matrix[76][224] * vector[76] +matrix[77][224] * vector[77] +matrix[78][224] * vector[78] +matrix[79][224] * vector[79] +matrix[80][224] * vector[80] +matrix[81][224] * vector[81] +matrix[82][224] * vector[82] +matrix[83][224] * vector[83] +matrix[84][224] * vector[84] +matrix[85][224] * vector[85] +matrix[86][224] * vector[86] +matrix[87][224] * vector[87] +matrix[88][224] * vector[88] +matrix[89][224] * vector[89] +matrix[90][224] * vector[90] +matrix[91][224] * vector[91] +matrix[92][224] * vector[92] +matrix[93][224] * vector[93] +matrix[94][224] * vector[94] +matrix[95][224] * vector[95] +matrix[96][224] * vector[96] +matrix[97][224] * vector[97] +matrix[98][224] * vector[98] +matrix[99][224] * vector[99] +b[224];
assign result[225] = matrix[0][225] * vector[0] +matrix[1][225] * vector[1] +matrix[2][225] * vector[2] +matrix[3][225] * vector[3] +matrix[4][225] * vector[4] +matrix[5][225] * vector[5] +matrix[6][225] * vector[6] +matrix[7][225] * vector[7] +matrix[8][225] * vector[8] +matrix[9][225] * vector[9] +matrix[10][225] * vector[10] +matrix[11][225] * vector[11] +matrix[12][225] * vector[12] +matrix[13][225] * vector[13] +matrix[14][225] * vector[14] +matrix[15][225] * vector[15] +matrix[16][225] * vector[16] +matrix[17][225] * vector[17] +matrix[18][225] * vector[18] +matrix[19][225] * vector[19] +matrix[20][225] * vector[20] +matrix[21][225] * vector[21] +matrix[22][225] * vector[22] +matrix[23][225] * vector[23] +matrix[24][225] * vector[24] +matrix[25][225] * vector[25] +matrix[26][225] * vector[26] +matrix[27][225] * vector[27] +matrix[28][225] * vector[28] +matrix[29][225] * vector[29] +matrix[30][225] * vector[30] +matrix[31][225] * vector[31] +matrix[32][225] * vector[32] +matrix[33][225] * vector[33] +matrix[34][225] * vector[34] +matrix[35][225] * vector[35] +matrix[36][225] * vector[36] +matrix[37][225] * vector[37] +matrix[38][225] * vector[38] +matrix[39][225] * vector[39] +matrix[40][225] * vector[40] +matrix[41][225] * vector[41] +matrix[42][225] * vector[42] +matrix[43][225] * vector[43] +matrix[44][225] * vector[44] +matrix[45][225] * vector[45] +matrix[46][225] * vector[46] +matrix[47][225] * vector[47] +matrix[48][225] * vector[48] +matrix[49][225] * vector[49] +matrix[50][225] * vector[50] +matrix[51][225] * vector[51] +matrix[52][225] * vector[52] +matrix[53][225] * vector[53] +matrix[54][225] * vector[54] +matrix[55][225] * vector[55] +matrix[56][225] * vector[56] +matrix[57][225] * vector[57] +matrix[58][225] * vector[58] +matrix[59][225] * vector[59] +matrix[60][225] * vector[60] +matrix[61][225] * vector[61] +matrix[62][225] * vector[62] +matrix[63][225] * vector[63] +matrix[64][225] * vector[64] +matrix[65][225] * vector[65] +matrix[66][225] * vector[66] +matrix[67][225] * vector[67] +matrix[68][225] * vector[68] +matrix[69][225] * vector[69] +matrix[70][225] * vector[70] +matrix[71][225] * vector[71] +matrix[72][225] * vector[72] +matrix[73][225] * vector[73] +matrix[74][225] * vector[74] +matrix[75][225] * vector[75] +matrix[76][225] * vector[76] +matrix[77][225] * vector[77] +matrix[78][225] * vector[78] +matrix[79][225] * vector[79] +matrix[80][225] * vector[80] +matrix[81][225] * vector[81] +matrix[82][225] * vector[82] +matrix[83][225] * vector[83] +matrix[84][225] * vector[84] +matrix[85][225] * vector[85] +matrix[86][225] * vector[86] +matrix[87][225] * vector[87] +matrix[88][225] * vector[88] +matrix[89][225] * vector[89] +matrix[90][225] * vector[90] +matrix[91][225] * vector[91] +matrix[92][225] * vector[92] +matrix[93][225] * vector[93] +matrix[94][225] * vector[94] +matrix[95][225] * vector[95] +matrix[96][225] * vector[96] +matrix[97][225] * vector[97] +matrix[98][225] * vector[98] +matrix[99][225] * vector[99] +b[225];
assign result[226] = matrix[0][226] * vector[0] +matrix[1][226] * vector[1] +matrix[2][226] * vector[2] +matrix[3][226] * vector[3] +matrix[4][226] * vector[4] +matrix[5][226] * vector[5] +matrix[6][226] * vector[6] +matrix[7][226] * vector[7] +matrix[8][226] * vector[8] +matrix[9][226] * vector[9] +matrix[10][226] * vector[10] +matrix[11][226] * vector[11] +matrix[12][226] * vector[12] +matrix[13][226] * vector[13] +matrix[14][226] * vector[14] +matrix[15][226] * vector[15] +matrix[16][226] * vector[16] +matrix[17][226] * vector[17] +matrix[18][226] * vector[18] +matrix[19][226] * vector[19] +matrix[20][226] * vector[20] +matrix[21][226] * vector[21] +matrix[22][226] * vector[22] +matrix[23][226] * vector[23] +matrix[24][226] * vector[24] +matrix[25][226] * vector[25] +matrix[26][226] * vector[26] +matrix[27][226] * vector[27] +matrix[28][226] * vector[28] +matrix[29][226] * vector[29] +matrix[30][226] * vector[30] +matrix[31][226] * vector[31] +matrix[32][226] * vector[32] +matrix[33][226] * vector[33] +matrix[34][226] * vector[34] +matrix[35][226] * vector[35] +matrix[36][226] * vector[36] +matrix[37][226] * vector[37] +matrix[38][226] * vector[38] +matrix[39][226] * vector[39] +matrix[40][226] * vector[40] +matrix[41][226] * vector[41] +matrix[42][226] * vector[42] +matrix[43][226] * vector[43] +matrix[44][226] * vector[44] +matrix[45][226] * vector[45] +matrix[46][226] * vector[46] +matrix[47][226] * vector[47] +matrix[48][226] * vector[48] +matrix[49][226] * vector[49] +matrix[50][226] * vector[50] +matrix[51][226] * vector[51] +matrix[52][226] * vector[52] +matrix[53][226] * vector[53] +matrix[54][226] * vector[54] +matrix[55][226] * vector[55] +matrix[56][226] * vector[56] +matrix[57][226] * vector[57] +matrix[58][226] * vector[58] +matrix[59][226] * vector[59] +matrix[60][226] * vector[60] +matrix[61][226] * vector[61] +matrix[62][226] * vector[62] +matrix[63][226] * vector[63] +matrix[64][226] * vector[64] +matrix[65][226] * vector[65] +matrix[66][226] * vector[66] +matrix[67][226] * vector[67] +matrix[68][226] * vector[68] +matrix[69][226] * vector[69] +matrix[70][226] * vector[70] +matrix[71][226] * vector[71] +matrix[72][226] * vector[72] +matrix[73][226] * vector[73] +matrix[74][226] * vector[74] +matrix[75][226] * vector[75] +matrix[76][226] * vector[76] +matrix[77][226] * vector[77] +matrix[78][226] * vector[78] +matrix[79][226] * vector[79] +matrix[80][226] * vector[80] +matrix[81][226] * vector[81] +matrix[82][226] * vector[82] +matrix[83][226] * vector[83] +matrix[84][226] * vector[84] +matrix[85][226] * vector[85] +matrix[86][226] * vector[86] +matrix[87][226] * vector[87] +matrix[88][226] * vector[88] +matrix[89][226] * vector[89] +matrix[90][226] * vector[90] +matrix[91][226] * vector[91] +matrix[92][226] * vector[92] +matrix[93][226] * vector[93] +matrix[94][226] * vector[94] +matrix[95][226] * vector[95] +matrix[96][226] * vector[96] +matrix[97][226] * vector[97] +matrix[98][226] * vector[98] +matrix[99][226] * vector[99] +b[226];
assign result[227] = matrix[0][227] * vector[0] +matrix[1][227] * vector[1] +matrix[2][227] * vector[2] +matrix[3][227] * vector[3] +matrix[4][227] * vector[4] +matrix[5][227] * vector[5] +matrix[6][227] * vector[6] +matrix[7][227] * vector[7] +matrix[8][227] * vector[8] +matrix[9][227] * vector[9] +matrix[10][227] * vector[10] +matrix[11][227] * vector[11] +matrix[12][227] * vector[12] +matrix[13][227] * vector[13] +matrix[14][227] * vector[14] +matrix[15][227] * vector[15] +matrix[16][227] * vector[16] +matrix[17][227] * vector[17] +matrix[18][227] * vector[18] +matrix[19][227] * vector[19] +matrix[20][227] * vector[20] +matrix[21][227] * vector[21] +matrix[22][227] * vector[22] +matrix[23][227] * vector[23] +matrix[24][227] * vector[24] +matrix[25][227] * vector[25] +matrix[26][227] * vector[26] +matrix[27][227] * vector[27] +matrix[28][227] * vector[28] +matrix[29][227] * vector[29] +matrix[30][227] * vector[30] +matrix[31][227] * vector[31] +matrix[32][227] * vector[32] +matrix[33][227] * vector[33] +matrix[34][227] * vector[34] +matrix[35][227] * vector[35] +matrix[36][227] * vector[36] +matrix[37][227] * vector[37] +matrix[38][227] * vector[38] +matrix[39][227] * vector[39] +matrix[40][227] * vector[40] +matrix[41][227] * vector[41] +matrix[42][227] * vector[42] +matrix[43][227] * vector[43] +matrix[44][227] * vector[44] +matrix[45][227] * vector[45] +matrix[46][227] * vector[46] +matrix[47][227] * vector[47] +matrix[48][227] * vector[48] +matrix[49][227] * vector[49] +matrix[50][227] * vector[50] +matrix[51][227] * vector[51] +matrix[52][227] * vector[52] +matrix[53][227] * vector[53] +matrix[54][227] * vector[54] +matrix[55][227] * vector[55] +matrix[56][227] * vector[56] +matrix[57][227] * vector[57] +matrix[58][227] * vector[58] +matrix[59][227] * vector[59] +matrix[60][227] * vector[60] +matrix[61][227] * vector[61] +matrix[62][227] * vector[62] +matrix[63][227] * vector[63] +matrix[64][227] * vector[64] +matrix[65][227] * vector[65] +matrix[66][227] * vector[66] +matrix[67][227] * vector[67] +matrix[68][227] * vector[68] +matrix[69][227] * vector[69] +matrix[70][227] * vector[70] +matrix[71][227] * vector[71] +matrix[72][227] * vector[72] +matrix[73][227] * vector[73] +matrix[74][227] * vector[74] +matrix[75][227] * vector[75] +matrix[76][227] * vector[76] +matrix[77][227] * vector[77] +matrix[78][227] * vector[78] +matrix[79][227] * vector[79] +matrix[80][227] * vector[80] +matrix[81][227] * vector[81] +matrix[82][227] * vector[82] +matrix[83][227] * vector[83] +matrix[84][227] * vector[84] +matrix[85][227] * vector[85] +matrix[86][227] * vector[86] +matrix[87][227] * vector[87] +matrix[88][227] * vector[88] +matrix[89][227] * vector[89] +matrix[90][227] * vector[90] +matrix[91][227] * vector[91] +matrix[92][227] * vector[92] +matrix[93][227] * vector[93] +matrix[94][227] * vector[94] +matrix[95][227] * vector[95] +matrix[96][227] * vector[96] +matrix[97][227] * vector[97] +matrix[98][227] * vector[98] +matrix[99][227] * vector[99] +b[227];
assign result[228] = matrix[0][228] * vector[0] +matrix[1][228] * vector[1] +matrix[2][228] * vector[2] +matrix[3][228] * vector[3] +matrix[4][228] * vector[4] +matrix[5][228] * vector[5] +matrix[6][228] * vector[6] +matrix[7][228] * vector[7] +matrix[8][228] * vector[8] +matrix[9][228] * vector[9] +matrix[10][228] * vector[10] +matrix[11][228] * vector[11] +matrix[12][228] * vector[12] +matrix[13][228] * vector[13] +matrix[14][228] * vector[14] +matrix[15][228] * vector[15] +matrix[16][228] * vector[16] +matrix[17][228] * vector[17] +matrix[18][228] * vector[18] +matrix[19][228] * vector[19] +matrix[20][228] * vector[20] +matrix[21][228] * vector[21] +matrix[22][228] * vector[22] +matrix[23][228] * vector[23] +matrix[24][228] * vector[24] +matrix[25][228] * vector[25] +matrix[26][228] * vector[26] +matrix[27][228] * vector[27] +matrix[28][228] * vector[28] +matrix[29][228] * vector[29] +matrix[30][228] * vector[30] +matrix[31][228] * vector[31] +matrix[32][228] * vector[32] +matrix[33][228] * vector[33] +matrix[34][228] * vector[34] +matrix[35][228] * vector[35] +matrix[36][228] * vector[36] +matrix[37][228] * vector[37] +matrix[38][228] * vector[38] +matrix[39][228] * vector[39] +matrix[40][228] * vector[40] +matrix[41][228] * vector[41] +matrix[42][228] * vector[42] +matrix[43][228] * vector[43] +matrix[44][228] * vector[44] +matrix[45][228] * vector[45] +matrix[46][228] * vector[46] +matrix[47][228] * vector[47] +matrix[48][228] * vector[48] +matrix[49][228] * vector[49] +matrix[50][228] * vector[50] +matrix[51][228] * vector[51] +matrix[52][228] * vector[52] +matrix[53][228] * vector[53] +matrix[54][228] * vector[54] +matrix[55][228] * vector[55] +matrix[56][228] * vector[56] +matrix[57][228] * vector[57] +matrix[58][228] * vector[58] +matrix[59][228] * vector[59] +matrix[60][228] * vector[60] +matrix[61][228] * vector[61] +matrix[62][228] * vector[62] +matrix[63][228] * vector[63] +matrix[64][228] * vector[64] +matrix[65][228] * vector[65] +matrix[66][228] * vector[66] +matrix[67][228] * vector[67] +matrix[68][228] * vector[68] +matrix[69][228] * vector[69] +matrix[70][228] * vector[70] +matrix[71][228] * vector[71] +matrix[72][228] * vector[72] +matrix[73][228] * vector[73] +matrix[74][228] * vector[74] +matrix[75][228] * vector[75] +matrix[76][228] * vector[76] +matrix[77][228] * vector[77] +matrix[78][228] * vector[78] +matrix[79][228] * vector[79] +matrix[80][228] * vector[80] +matrix[81][228] * vector[81] +matrix[82][228] * vector[82] +matrix[83][228] * vector[83] +matrix[84][228] * vector[84] +matrix[85][228] * vector[85] +matrix[86][228] * vector[86] +matrix[87][228] * vector[87] +matrix[88][228] * vector[88] +matrix[89][228] * vector[89] +matrix[90][228] * vector[90] +matrix[91][228] * vector[91] +matrix[92][228] * vector[92] +matrix[93][228] * vector[93] +matrix[94][228] * vector[94] +matrix[95][228] * vector[95] +matrix[96][228] * vector[96] +matrix[97][228] * vector[97] +matrix[98][228] * vector[98] +matrix[99][228] * vector[99] +b[228];
assign result[229] = matrix[0][229] * vector[0] +matrix[1][229] * vector[1] +matrix[2][229] * vector[2] +matrix[3][229] * vector[3] +matrix[4][229] * vector[4] +matrix[5][229] * vector[5] +matrix[6][229] * vector[6] +matrix[7][229] * vector[7] +matrix[8][229] * vector[8] +matrix[9][229] * vector[9] +matrix[10][229] * vector[10] +matrix[11][229] * vector[11] +matrix[12][229] * vector[12] +matrix[13][229] * vector[13] +matrix[14][229] * vector[14] +matrix[15][229] * vector[15] +matrix[16][229] * vector[16] +matrix[17][229] * vector[17] +matrix[18][229] * vector[18] +matrix[19][229] * vector[19] +matrix[20][229] * vector[20] +matrix[21][229] * vector[21] +matrix[22][229] * vector[22] +matrix[23][229] * vector[23] +matrix[24][229] * vector[24] +matrix[25][229] * vector[25] +matrix[26][229] * vector[26] +matrix[27][229] * vector[27] +matrix[28][229] * vector[28] +matrix[29][229] * vector[29] +matrix[30][229] * vector[30] +matrix[31][229] * vector[31] +matrix[32][229] * vector[32] +matrix[33][229] * vector[33] +matrix[34][229] * vector[34] +matrix[35][229] * vector[35] +matrix[36][229] * vector[36] +matrix[37][229] * vector[37] +matrix[38][229] * vector[38] +matrix[39][229] * vector[39] +matrix[40][229] * vector[40] +matrix[41][229] * vector[41] +matrix[42][229] * vector[42] +matrix[43][229] * vector[43] +matrix[44][229] * vector[44] +matrix[45][229] * vector[45] +matrix[46][229] * vector[46] +matrix[47][229] * vector[47] +matrix[48][229] * vector[48] +matrix[49][229] * vector[49] +matrix[50][229] * vector[50] +matrix[51][229] * vector[51] +matrix[52][229] * vector[52] +matrix[53][229] * vector[53] +matrix[54][229] * vector[54] +matrix[55][229] * vector[55] +matrix[56][229] * vector[56] +matrix[57][229] * vector[57] +matrix[58][229] * vector[58] +matrix[59][229] * vector[59] +matrix[60][229] * vector[60] +matrix[61][229] * vector[61] +matrix[62][229] * vector[62] +matrix[63][229] * vector[63] +matrix[64][229] * vector[64] +matrix[65][229] * vector[65] +matrix[66][229] * vector[66] +matrix[67][229] * vector[67] +matrix[68][229] * vector[68] +matrix[69][229] * vector[69] +matrix[70][229] * vector[70] +matrix[71][229] * vector[71] +matrix[72][229] * vector[72] +matrix[73][229] * vector[73] +matrix[74][229] * vector[74] +matrix[75][229] * vector[75] +matrix[76][229] * vector[76] +matrix[77][229] * vector[77] +matrix[78][229] * vector[78] +matrix[79][229] * vector[79] +matrix[80][229] * vector[80] +matrix[81][229] * vector[81] +matrix[82][229] * vector[82] +matrix[83][229] * vector[83] +matrix[84][229] * vector[84] +matrix[85][229] * vector[85] +matrix[86][229] * vector[86] +matrix[87][229] * vector[87] +matrix[88][229] * vector[88] +matrix[89][229] * vector[89] +matrix[90][229] * vector[90] +matrix[91][229] * vector[91] +matrix[92][229] * vector[92] +matrix[93][229] * vector[93] +matrix[94][229] * vector[94] +matrix[95][229] * vector[95] +matrix[96][229] * vector[96] +matrix[97][229] * vector[97] +matrix[98][229] * vector[98] +matrix[99][229] * vector[99] +b[229];
assign result[230] = matrix[0][230] * vector[0] +matrix[1][230] * vector[1] +matrix[2][230] * vector[2] +matrix[3][230] * vector[3] +matrix[4][230] * vector[4] +matrix[5][230] * vector[5] +matrix[6][230] * vector[6] +matrix[7][230] * vector[7] +matrix[8][230] * vector[8] +matrix[9][230] * vector[9] +matrix[10][230] * vector[10] +matrix[11][230] * vector[11] +matrix[12][230] * vector[12] +matrix[13][230] * vector[13] +matrix[14][230] * vector[14] +matrix[15][230] * vector[15] +matrix[16][230] * vector[16] +matrix[17][230] * vector[17] +matrix[18][230] * vector[18] +matrix[19][230] * vector[19] +matrix[20][230] * vector[20] +matrix[21][230] * vector[21] +matrix[22][230] * vector[22] +matrix[23][230] * vector[23] +matrix[24][230] * vector[24] +matrix[25][230] * vector[25] +matrix[26][230] * vector[26] +matrix[27][230] * vector[27] +matrix[28][230] * vector[28] +matrix[29][230] * vector[29] +matrix[30][230] * vector[30] +matrix[31][230] * vector[31] +matrix[32][230] * vector[32] +matrix[33][230] * vector[33] +matrix[34][230] * vector[34] +matrix[35][230] * vector[35] +matrix[36][230] * vector[36] +matrix[37][230] * vector[37] +matrix[38][230] * vector[38] +matrix[39][230] * vector[39] +matrix[40][230] * vector[40] +matrix[41][230] * vector[41] +matrix[42][230] * vector[42] +matrix[43][230] * vector[43] +matrix[44][230] * vector[44] +matrix[45][230] * vector[45] +matrix[46][230] * vector[46] +matrix[47][230] * vector[47] +matrix[48][230] * vector[48] +matrix[49][230] * vector[49] +matrix[50][230] * vector[50] +matrix[51][230] * vector[51] +matrix[52][230] * vector[52] +matrix[53][230] * vector[53] +matrix[54][230] * vector[54] +matrix[55][230] * vector[55] +matrix[56][230] * vector[56] +matrix[57][230] * vector[57] +matrix[58][230] * vector[58] +matrix[59][230] * vector[59] +matrix[60][230] * vector[60] +matrix[61][230] * vector[61] +matrix[62][230] * vector[62] +matrix[63][230] * vector[63] +matrix[64][230] * vector[64] +matrix[65][230] * vector[65] +matrix[66][230] * vector[66] +matrix[67][230] * vector[67] +matrix[68][230] * vector[68] +matrix[69][230] * vector[69] +matrix[70][230] * vector[70] +matrix[71][230] * vector[71] +matrix[72][230] * vector[72] +matrix[73][230] * vector[73] +matrix[74][230] * vector[74] +matrix[75][230] * vector[75] +matrix[76][230] * vector[76] +matrix[77][230] * vector[77] +matrix[78][230] * vector[78] +matrix[79][230] * vector[79] +matrix[80][230] * vector[80] +matrix[81][230] * vector[81] +matrix[82][230] * vector[82] +matrix[83][230] * vector[83] +matrix[84][230] * vector[84] +matrix[85][230] * vector[85] +matrix[86][230] * vector[86] +matrix[87][230] * vector[87] +matrix[88][230] * vector[88] +matrix[89][230] * vector[89] +matrix[90][230] * vector[90] +matrix[91][230] * vector[91] +matrix[92][230] * vector[92] +matrix[93][230] * vector[93] +matrix[94][230] * vector[94] +matrix[95][230] * vector[95] +matrix[96][230] * vector[96] +matrix[97][230] * vector[97] +matrix[98][230] * vector[98] +matrix[99][230] * vector[99] +b[230];
assign result[231] = matrix[0][231] * vector[0] +matrix[1][231] * vector[1] +matrix[2][231] * vector[2] +matrix[3][231] * vector[3] +matrix[4][231] * vector[4] +matrix[5][231] * vector[5] +matrix[6][231] * vector[6] +matrix[7][231] * vector[7] +matrix[8][231] * vector[8] +matrix[9][231] * vector[9] +matrix[10][231] * vector[10] +matrix[11][231] * vector[11] +matrix[12][231] * vector[12] +matrix[13][231] * vector[13] +matrix[14][231] * vector[14] +matrix[15][231] * vector[15] +matrix[16][231] * vector[16] +matrix[17][231] * vector[17] +matrix[18][231] * vector[18] +matrix[19][231] * vector[19] +matrix[20][231] * vector[20] +matrix[21][231] * vector[21] +matrix[22][231] * vector[22] +matrix[23][231] * vector[23] +matrix[24][231] * vector[24] +matrix[25][231] * vector[25] +matrix[26][231] * vector[26] +matrix[27][231] * vector[27] +matrix[28][231] * vector[28] +matrix[29][231] * vector[29] +matrix[30][231] * vector[30] +matrix[31][231] * vector[31] +matrix[32][231] * vector[32] +matrix[33][231] * vector[33] +matrix[34][231] * vector[34] +matrix[35][231] * vector[35] +matrix[36][231] * vector[36] +matrix[37][231] * vector[37] +matrix[38][231] * vector[38] +matrix[39][231] * vector[39] +matrix[40][231] * vector[40] +matrix[41][231] * vector[41] +matrix[42][231] * vector[42] +matrix[43][231] * vector[43] +matrix[44][231] * vector[44] +matrix[45][231] * vector[45] +matrix[46][231] * vector[46] +matrix[47][231] * vector[47] +matrix[48][231] * vector[48] +matrix[49][231] * vector[49] +matrix[50][231] * vector[50] +matrix[51][231] * vector[51] +matrix[52][231] * vector[52] +matrix[53][231] * vector[53] +matrix[54][231] * vector[54] +matrix[55][231] * vector[55] +matrix[56][231] * vector[56] +matrix[57][231] * vector[57] +matrix[58][231] * vector[58] +matrix[59][231] * vector[59] +matrix[60][231] * vector[60] +matrix[61][231] * vector[61] +matrix[62][231] * vector[62] +matrix[63][231] * vector[63] +matrix[64][231] * vector[64] +matrix[65][231] * vector[65] +matrix[66][231] * vector[66] +matrix[67][231] * vector[67] +matrix[68][231] * vector[68] +matrix[69][231] * vector[69] +matrix[70][231] * vector[70] +matrix[71][231] * vector[71] +matrix[72][231] * vector[72] +matrix[73][231] * vector[73] +matrix[74][231] * vector[74] +matrix[75][231] * vector[75] +matrix[76][231] * vector[76] +matrix[77][231] * vector[77] +matrix[78][231] * vector[78] +matrix[79][231] * vector[79] +matrix[80][231] * vector[80] +matrix[81][231] * vector[81] +matrix[82][231] * vector[82] +matrix[83][231] * vector[83] +matrix[84][231] * vector[84] +matrix[85][231] * vector[85] +matrix[86][231] * vector[86] +matrix[87][231] * vector[87] +matrix[88][231] * vector[88] +matrix[89][231] * vector[89] +matrix[90][231] * vector[90] +matrix[91][231] * vector[91] +matrix[92][231] * vector[92] +matrix[93][231] * vector[93] +matrix[94][231] * vector[94] +matrix[95][231] * vector[95] +matrix[96][231] * vector[96] +matrix[97][231] * vector[97] +matrix[98][231] * vector[98] +matrix[99][231] * vector[99] +b[231];
assign result[232] = matrix[0][232] * vector[0] +matrix[1][232] * vector[1] +matrix[2][232] * vector[2] +matrix[3][232] * vector[3] +matrix[4][232] * vector[4] +matrix[5][232] * vector[5] +matrix[6][232] * vector[6] +matrix[7][232] * vector[7] +matrix[8][232] * vector[8] +matrix[9][232] * vector[9] +matrix[10][232] * vector[10] +matrix[11][232] * vector[11] +matrix[12][232] * vector[12] +matrix[13][232] * vector[13] +matrix[14][232] * vector[14] +matrix[15][232] * vector[15] +matrix[16][232] * vector[16] +matrix[17][232] * vector[17] +matrix[18][232] * vector[18] +matrix[19][232] * vector[19] +matrix[20][232] * vector[20] +matrix[21][232] * vector[21] +matrix[22][232] * vector[22] +matrix[23][232] * vector[23] +matrix[24][232] * vector[24] +matrix[25][232] * vector[25] +matrix[26][232] * vector[26] +matrix[27][232] * vector[27] +matrix[28][232] * vector[28] +matrix[29][232] * vector[29] +matrix[30][232] * vector[30] +matrix[31][232] * vector[31] +matrix[32][232] * vector[32] +matrix[33][232] * vector[33] +matrix[34][232] * vector[34] +matrix[35][232] * vector[35] +matrix[36][232] * vector[36] +matrix[37][232] * vector[37] +matrix[38][232] * vector[38] +matrix[39][232] * vector[39] +matrix[40][232] * vector[40] +matrix[41][232] * vector[41] +matrix[42][232] * vector[42] +matrix[43][232] * vector[43] +matrix[44][232] * vector[44] +matrix[45][232] * vector[45] +matrix[46][232] * vector[46] +matrix[47][232] * vector[47] +matrix[48][232] * vector[48] +matrix[49][232] * vector[49] +matrix[50][232] * vector[50] +matrix[51][232] * vector[51] +matrix[52][232] * vector[52] +matrix[53][232] * vector[53] +matrix[54][232] * vector[54] +matrix[55][232] * vector[55] +matrix[56][232] * vector[56] +matrix[57][232] * vector[57] +matrix[58][232] * vector[58] +matrix[59][232] * vector[59] +matrix[60][232] * vector[60] +matrix[61][232] * vector[61] +matrix[62][232] * vector[62] +matrix[63][232] * vector[63] +matrix[64][232] * vector[64] +matrix[65][232] * vector[65] +matrix[66][232] * vector[66] +matrix[67][232] * vector[67] +matrix[68][232] * vector[68] +matrix[69][232] * vector[69] +matrix[70][232] * vector[70] +matrix[71][232] * vector[71] +matrix[72][232] * vector[72] +matrix[73][232] * vector[73] +matrix[74][232] * vector[74] +matrix[75][232] * vector[75] +matrix[76][232] * vector[76] +matrix[77][232] * vector[77] +matrix[78][232] * vector[78] +matrix[79][232] * vector[79] +matrix[80][232] * vector[80] +matrix[81][232] * vector[81] +matrix[82][232] * vector[82] +matrix[83][232] * vector[83] +matrix[84][232] * vector[84] +matrix[85][232] * vector[85] +matrix[86][232] * vector[86] +matrix[87][232] * vector[87] +matrix[88][232] * vector[88] +matrix[89][232] * vector[89] +matrix[90][232] * vector[90] +matrix[91][232] * vector[91] +matrix[92][232] * vector[92] +matrix[93][232] * vector[93] +matrix[94][232] * vector[94] +matrix[95][232] * vector[95] +matrix[96][232] * vector[96] +matrix[97][232] * vector[97] +matrix[98][232] * vector[98] +matrix[99][232] * vector[99] +b[232];
assign result[233] = matrix[0][233] * vector[0] +matrix[1][233] * vector[1] +matrix[2][233] * vector[2] +matrix[3][233] * vector[3] +matrix[4][233] * vector[4] +matrix[5][233] * vector[5] +matrix[6][233] * vector[6] +matrix[7][233] * vector[7] +matrix[8][233] * vector[8] +matrix[9][233] * vector[9] +matrix[10][233] * vector[10] +matrix[11][233] * vector[11] +matrix[12][233] * vector[12] +matrix[13][233] * vector[13] +matrix[14][233] * vector[14] +matrix[15][233] * vector[15] +matrix[16][233] * vector[16] +matrix[17][233] * vector[17] +matrix[18][233] * vector[18] +matrix[19][233] * vector[19] +matrix[20][233] * vector[20] +matrix[21][233] * vector[21] +matrix[22][233] * vector[22] +matrix[23][233] * vector[23] +matrix[24][233] * vector[24] +matrix[25][233] * vector[25] +matrix[26][233] * vector[26] +matrix[27][233] * vector[27] +matrix[28][233] * vector[28] +matrix[29][233] * vector[29] +matrix[30][233] * vector[30] +matrix[31][233] * vector[31] +matrix[32][233] * vector[32] +matrix[33][233] * vector[33] +matrix[34][233] * vector[34] +matrix[35][233] * vector[35] +matrix[36][233] * vector[36] +matrix[37][233] * vector[37] +matrix[38][233] * vector[38] +matrix[39][233] * vector[39] +matrix[40][233] * vector[40] +matrix[41][233] * vector[41] +matrix[42][233] * vector[42] +matrix[43][233] * vector[43] +matrix[44][233] * vector[44] +matrix[45][233] * vector[45] +matrix[46][233] * vector[46] +matrix[47][233] * vector[47] +matrix[48][233] * vector[48] +matrix[49][233] * vector[49] +matrix[50][233] * vector[50] +matrix[51][233] * vector[51] +matrix[52][233] * vector[52] +matrix[53][233] * vector[53] +matrix[54][233] * vector[54] +matrix[55][233] * vector[55] +matrix[56][233] * vector[56] +matrix[57][233] * vector[57] +matrix[58][233] * vector[58] +matrix[59][233] * vector[59] +matrix[60][233] * vector[60] +matrix[61][233] * vector[61] +matrix[62][233] * vector[62] +matrix[63][233] * vector[63] +matrix[64][233] * vector[64] +matrix[65][233] * vector[65] +matrix[66][233] * vector[66] +matrix[67][233] * vector[67] +matrix[68][233] * vector[68] +matrix[69][233] * vector[69] +matrix[70][233] * vector[70] +matrix[71][233] * vector[71] +matrix[72][233] * vector[72] +matrix[73][233] * vector[73] +matrix[74][233] * vector[74] +matrix[75][233] * vector[75] +matrix[76][233] * vector[76] +matrix[77][233] * vector[77] +matrix[78][233] * vector[78] +matrix[79][233] * vector[79] +matrix[80][233] * vector[80] +matrix[81][233] * vector[81] +matrix[82][233] * vector[82] +matrix[83][233] * vector[83] +matrix[84][233] * vector[84] +matrix[85][233] * vector[85] +matrix[86][233] * vector[86] +matrix[87][233] * vector[87] +matrix[88][233] * vector[88] +matrix[89][233] * vector[89] +matrix[90][233] * vector[90] +matrix[91][233] * vector[91] +matrix[92][233] * vector[92] +matrix[93][233] * vector[93] +matrix[94][233] * vector[94] +matrix[95][233] * vector[95] +matrix[96][233] * vector[96] +matrix[97][233] * vector[97] +matrix[98][233] * vector[98] +matrix[99][233] * vector[99] +b[233];
assign result[234] = matrix[0][234] * vector[0] +matrix[1][234] * vector[1] +matrix[2][234] * vector[2] +matrix[3][234] * vector[3] +matrix[4][234] * vector[4] +matrix[5][234] * vector[5] +matrix[6][234] * vector[6] +matrix[7][234] * vector[7] +matrix[8][234] * vector[8] +matrix[9][234] * vector[9] +matrix[10][234] * vector[10] +matrix[11][234] * vector[11] +matrix[12][234] * vector[12] +matrix[13][234] * vector[13] +matrix[14][234] * vector[14] +matrix[15][234] * vector[15] +matrix[16][234] * vector[16] +matrix[17][234] * vector[17] +matrix[18][234] * vector[18] +matrix[19][234] * vector[19] +matrix[20][234] * vector[20] +matrix[21][234] * vector[21] +matrix[22][234] * vector[22] +matrix[23][234] * vector[23] +matrix[24][234] * vector[24] +matrix[25][234] * vector[25] +matrix[26][234] * vector[26] +matrix[27][234] * vector[27] +matrix[28][234] * vector[28] +matrix[29][234] * vector[29] +matrix[30][234] * vector[30] +matrix[31][234] * vector[31] +matrix[32][234] * vector[32] +matrix[33][234] * vector[33] +matrix[34][234] * vector[34] +matrix[35][234] * vector[35] +matrix[36][234] * vector[36] +matrix[37][234] * vector[37] +matrix[38][234] * vector[38] +matrix[39][234] * vector[39] +matrix[40][234] * vector[40] +matrix[41][234] * vector[41] +matrix[42][234] * vector[42] +matrix[43][234] * vector[43] +matrix[44][234] * vector[44] +matrix[45][234] * vector[45] +matrix[46][234] * vector[46] +matrix[47][234] * vector[47] +matrix[48][234] * vector[48] +matrix[49][234] * vector[49] +matrix[50][234] * vector[50] +matrix[51][234] * vector[51] +matrix[52][234] * vector[52] +matrix[53][234] * vector[53] +matrix[54][234] * vector[54] +matrix[55][234] * vector[55] +matrix[56][234] * vector[56] +matrix[57][234] * vector[57] +matrix[58][234] * vector[58] +matrix[59][234] * vector[59] +matrix[60][234] * vector[60] +matrix[61][234] * vector[61] +matrix[62][234] * vector[62] +matrix[63][234] * vector[63] +matrix[64][234] * vector[64] +matrix[65][234] * vector[65] +matrix[66][234] * vector[66] +matrix[67][234] * vector[67] +matrix[68][234] * vector[68] +matrix[69][234] * vector[69] +matrix[70][234] * vector[70] +matrix[71][234] * vector[71] +matrix[72][234] * vector[72] +matrix[73][234] * vector[73] +matrix[74][234] * vector[74] +matrix[75][234] * vector[75] +matrix[76][234] * vector[76] +matrix[77][234] * vector[77] +matrix[78][234] * vector[78] +matrix[79][234] * vector[79] +matrix[80][234] * vector[80] +matrix[81][234] * vector[81] +matrix[82][234] * vector[82] +matrix[83][234] * vector[83] +matrix[84][234] * vector[84] +matrix[85][234] * vector[85] +matrix[86][234] * vector[86] +matrix[87][234] * vector[87] +matrix[88][234] * vector[88] +matrix[89][234] * vector[89] +matrix[90][234] * vector[90] +matrix[91][234] * vector[91] +matrix[92][234] * vector[92] +matrix[93][234] * vector[93] +matrix[94][234] * vector[94] +matrix[95][234] * vector[95] +matrix[96][234] * vector[96] +matrix[97][234] * vector[97] +matrix[98][234] * vector[98] +matrix[99][234] * vector[99] +b[234];
assign result[235] = matrix[0][235] * vector[0] +matrix[1][235] * vector[1] +matrix[2][235] * vector[2] +matrix[3][235] * vector[3] +matrix[4][235] * vector[4] +matrix[5][235] * vector[5] +matrix[6][235] * vector[6] +matrix[7][235] * vector[7] +matrix[8][235] * vector[8] +matrix[9][235] * vector[9] +matrix[10][235] * vector[10] +matrix[11][235] * vector[11] +matrix[12][235] * vector[12] +matrix[13][235] * vector[13] +matrix[14][235] * vector[14] +matrix[15][235] * vector[15] +matrix[16][235] * vector[16] +matrix[17][235] * vector[17] +matrix[18][235] * vector[18] +matrix[19][235] * vector[19] +matrix[20][235] * vector[20] +matrix[21][235] * vector[21] +matrix[22][235] * vector[22] +matrix[23][235] * vector[23] +matrix[24][235] * vector[24] +matrix[25][235] * vector[25] +matrix[26][235] * vector[26] +matrix[27][235] * vector[27] +matrix[28][235] * vector[28] +matrix[29][235] * vector[29] +matrix[30][235] * vector[30] +matrix[31][235] * vector[31] +matrix[32][235] * vector[32] +matrix[33][235] * vector[33] +matrix[34][235] * vector[34] +matrix[35][235] * vector[35] +matrix[36][235] * vector[36] +matrix[37][235] * vector[37] +matrix[38][235] * vector[38] +matrix[39][235] * vector[39] +matrix[40][235] * vector[40] +matrix[41][235] * vector[41] +matrix[42][235] * vector[42] +matrix[43][235] * vector[43] +matrix[44][235] * vector[44] +matrix[45][235] * vector[45] +matrix[46][235] * vector[46] +matrix[47][235] * vector[47] +matrix[48][235] * vector[48] +matrix[49][235] * vector[49] +matrix[50][235] * vector[50] +matrix[51][235] * vector[51] +matrix[52][235] * vector[52] +matrix[53][235] * vector[53] +matrix[54][235] * vector[54] +matrix[55][235] * vector[55] +matrix[56][235] * vector[56] +matrix[57][235] * vector[57] +matrix[58][235] * vector[58] +matrix[59][235] * vector[59] +matrix[60][235] * vector[60] +matrix[61][235] * vector[61] +matrix[62][235] * vector[62] +matrix[63][235] * vector[63] +matrix[64][235] * vector[64] +matrix[65][235] * vector[65] +matrix[66][235] * vector[66] +matrix[67][235] * vector[67] +matrix[68][235] * vector[68] +matrix[69][235] * vector[69] +matrix[70][235] * vector[70] +matrix[71][235] * vector[71] +matrix[72][235] * vector[72] +matrix[73][235] * vector[73] +matrix[74][235] * vector[74] +matrix[75][235] * vector[75] +matrix[76][235] * vector[76] +matrix[77][235] * vector[77] +matrix[78][235] * vector[78] +matrix[79][235] * vector[79] +matrix[80][235] * vector[80] +matrix[81][235] * vector[81] +matrix[82][235] * vector[82] +matrix[83][235] * vector[83] +matrix[84][235] * vector[84] +matrix[85][235] * vector[85] +matrix[86][235] * vector[86] +matrix[87][235] * vector[87] +matrix[88][235] * vector[88] +matrix[89][235] * vector[89] +matrix[90][235] * vector[90] +matrix[91][235] * vector[91] +matrix[92][235] * vector[92] +matrix[93][235] * vector[93] +matrix[94][235] * vector[94] +matrix[95][235] * vector[95] +matrix[96][235] * vector[96] +matrix[97][235] * vector[97] +matrix[98][235] * vector[98] +matrix[99][235] * vector[99] +b[235];
assign result[236] = matrix[0][236] * vector[0] +matrix[1][236] * vector[1] +matrix[2][236] * vector[2] +matrix[3][236] * vector[3] +matrix[4][236] * vector[4] +matrix[5][236] * vector[5] +matrix[6][236] * vector[6] +matrix[7][236] * vector[7] +matrix[8][236] * vector[8] +matrix[9][236] * vector[9] +matrix[10][236] * vector[10] +matrix[11][236] * vector[11] +matrix[12][236] * vector[12] +matrix[13][236] * vector[13] +matrix[14][236] * vector[14] +matrix[15][236] * vector[15] +matrix[16][236] * vector[16] +matrix[17][236] * vector[17] +matrix[18][236] * vector[18] +matrix[19][236] * vector[19] +matrix[20][236] * vector[20] +matrix[21][236] * vector[21] +matrix[22][236] * vector[22] +matrix[23][236] * vector[23] +matrix[24][236] * vector[24] +matrix[25][236] * vector[25] +matrix[26][236] * vector[26] +matrix[27][236] * vector[27] +matrix[28][236] * vector[28] +matrix[29][236] * vector[29] +matrix[30][236] * vector[30] +matrix[31][236] * vector[31] +matrix[32][236] * vector[32] +matrix[33][236] * vector[33] +matrix[34][236] * vector[34] +matrix[35][236] * vector[35] +matrix[36][236] * vector[36] +matrix[37][236] * vector[37] +matrix[38][236] * vector[38] +matrix[39][236] * vector[39] +matrix[40][236] * vector[40] +matrix[41][236] * vector[41] +matrix[42][236] * vector[42] +matrix[43][236] * vector[43] +matrix[44][236] * vector[44] +matrix[45][236] * vector[45] +matrix[46][236] * vector[46] +matrix[47][236] * vector[47] +matrix[48][236] * vector[48] +matrix[49][236] * vector[49] +matrix[50][236] * vector[50] +matrix[51][236] * vector[51] +matrix[52][236] * vector[52] +matrix[53][236] * vector[53] +matrix[54][236] * vector[54] +matrix[55][236] * vector[55] +matrix[56][236] * vector[56] +matrix[57][236] * vector[57] +matrix[58][236] * vector[58] +matrix[59][236] * vector[59] +matrix[60][236] * vector[60] +matrix[61][236] * vector[61] +matrix[62][236] * vector[62] +matrix[63][236] * vector[63] +matrix[64][236] * vector[64] +matrix[65][236] * vector[65] +matrix[66][236] * vector[66] +matrix[67][236] * vector[67] +matrix[68][236] * vector[68] +matrix[69][236] * vector[69] +matrix[70][236] * vector[70] +matrix[71][236] * vector[71] +matrix[72][236] * vector[72] +matrix[73][236] * vector[73] +matrix[74][236] * vector[74] +matrix[75][236] * vector[75] +matrix[76][236] * vector[76] +matrix[77][236] * vector[77] +matrix[78][236] * vector[78] +matrix[79][236] * vector[79] +matrix[80][236] * vector[80] +matrix[81][236] * vector[81] +matrix[82][236] * vector[82] +matrix[83][236] * vector[83] +matrix[84][236] * vector[84] +matrix[85][236] * vector[85] +matrix[86][236] * vector[86] +matrix[87][236] * vector[87] +matrix[88][236] * vector[88] +matrix[89][236] * vector[89] +matrix[90][236] * vector[90] +matrix[91][236] * vector[91] +matrix[92][236] * vector[92] +matrix[93][236] * vector[93] +matrix[94][236] * vector[94] +matrix[95][236] * vector[95] +matrix[96][236] * vector[96] +matrix[97][236] * vector[97] +matrix[98][236] * vector[98] +matrix[99][236] * vector[99] +b[236];
assign result[237] = matrix[0][237] * vector[0] +matrix[1][237] * vector[1] +matrix[2][237] * vector[2] +matrix[3][237] * vector[3] +matrix[4][237] * vector[4] +matrix[5][237] * vector[5] +matrix[6][237] * vector[6] +matrix[7][237] * vector[7] +matrix[8][237] * vector[8] +matrix[9][237] * vector[9] +matrix[10][237] * vector[10] +matrix[11][237] * vector[11] +matrix[12][237] * vector[12] +matrix[13][237] * vector[13] +matrix[14][237] * vector[14] +matrix[15][237] * vector[15] +matrix[16][237] * vector[16] +matrix[17][237] * vector[17] +matrix[18][237] * vector[18] +matrix[19][237] * vector[19] +matrix[20][237] * vector[20] +matrix[21][237] * vector[21] +matrix[22][237] * vector[22] +matrix[23][237] * vector[23] +matrix[24][237] * vector[24] +matrix[25][237] * vector[25] +matrix[26][237] * vector[26] +matrix[27][237] * vector[27] +matrix[28][237] * vector[28] +matrix[29][237] * vector[29] +matrix[30][237] * vector[30] +matrix[31][237] * vector[31] +matrix[32][237] * vector[32] +matrix[33][237] * vector[33] +matrix[34][237] * vector[34] +matrix[35][237] * vector[35] +matrix[36][237] * vector[36] +matrix[37][237] * vector[37] +matrix[38][237] * vector[38] +matrix[39][237] * vector[39] +matrix[40][237] * vector[40] +matrix[41][237] * vector[41] +matrix[42][237] * vector[42] +matrix[43][237] * vector[43] +matrix[44][237] * vector[44] +matrix[45][237] * vector[45] +matrix[46][237] * vector[46] +matrix[47][237] * vector[47] +matrix[48][237] * vector[48] +matrix[49][237] * vector[49] +matrix[50][237] * vector[50] +matrix[51][237] * vector[51] +matrix[52][237] * vector[52] +matrix[53][237] * vector[53] +matrix[54][237] * vector[54] +matrix[55][237] * vector[55] +matrix[56][237] * vector[56] +matrix[57][237] * vector[57] +matrix[58][237] * vector[58] +matrix[59][237] * vector[59] +matrix[60][237] * vector[60] +matrix[61][237] * vector[61] +matrix[62][237] * vector[62] +matrix[63][237] * vector[63] +matrix[64][237] * vector[64] +matrix[65][237] * vector[65] +matrix[66][237] * vector[66] +matrix[67][237] * vector[67] +matrix[68][237] * vector[68] +matrix[69][237] * vector[69] +matrix[70][237] * vector[70] +matrix[71][237] * vector[71] +matrix[72][237] * vector[72] +matrix[73][237] * vector[73] +matrix[74][237] * vector[74] +matrix[75][237] * vector[75] +matrix[76][237] * vector[76] +matrix[77][237] * vector[77] +matrix[78][237] * vector[78] +matrix[79][237] * vector[79] +matrix[80][237] * vector[80] +matrix[81][237] * vector[81] +matrix[82][237] * vector[82] +matrix[83][237] * vector[83] +matrix[84][237] * vector[84] +matrix[85][237] * vector[85] +matrix[86][237] * vector[86] +matrix[87][237] * vector[87] +matrix[88][237] * vector[88] +matrix[89][237] * vector[89] +matrix[90][237] * vector[90] +matrix[91][237] * vector[91] +matrix[92][237] * vector[92] +matrix[93][237] * vector[93] +matrix[94][237] * vector[94] +matrix[95][237] * vector[95] +matrix[96][237] * vector[96] +matrix[97][237] * vector[97] +matrix[98][237] * vector[98] +matrix[99][237] * vector[99] +b[237];
assign result[238] = matrix[0][238] * vector[0] +matrix[1][238] * vector[1] +matrix[2][238] * vector[2] +matrix[3][238] * vector[3] +matrix[4][238] * vector[4] +matrix[5][238] * vector[5] +matrix[6][238] * vector[6] +matrix[7][238] * vector[7] +matrix[8][238] * vector[8] +matrix[9][238] * vector[9] +matrix[10][238] * vector[10] +matrix[11][238] * vector[11] +matrix[12][238] * vector[12] +matrix[13][238] * vector[13] +matrix[14][238] * vector[14] +matrix[15][238] * vector[15] +matrix[16][238] * vector[16] +matrix[17][238] * vector[17] +matrix[18][238] * vector[18] +matrix[19][238] * vector[19] +matrix[20][238] * vector[20] +matrix[21][238] * vector[21] +matrix[22][238] * vector[22] +matrix[23][238] * vector[23] +matrix[24][238] * vector[24] +matrix[25][238] * vector[25] +matrix[26][238] * vector[26] +matrix[27][238] * vector[27] +matrix[28][238] * vector[28] +matrix[29][238] * vector[29] +matrix[30][238] * vector[30] +matrix[31][238] * vector[31] +matrix[32][238] * vector[32] +matrix[33][238] * vector[33] +matrix[34][238] * vector[34] +matrix[35][238] * vector[35] +matrix[36][238] * vector[36] +matrix[37][238] * vector[37] +matrix[38][238] * vector[38] +matrix[39][238] * vector[39] +matrix[40][238] * vector[40] +matrix[41][238] * vector[41] +matrix[42][238] * vector[42] +matrix[43][238] * vector[43] +matrix[44][238] * vector[44] +matrix[45][238] * vector[45] +matrix[46][238] * vector[46] +matrix[47][238] * vector[47] +matrix[48][238] * vector[48] +matrix[49][238] * vector[49] +matrix[50][238] * vector[50] +matrix[51][238] * vector[51] +matrix[52][238] * vector[52] +matrix[53][238] * vector[53] +matrix[54][238] * vector[54] +matrix[55][238] * vector[55] +matrix[56][238] * vector[56] +matrix[57][238] * vector[57] +matrix[58][238] * vector[58] +matrix[59][238] * vector[59] +matrix[60][238] * vector[60] +matrix[61][238] * vector[61] +matrix[62][238] * vector[62] +matrix[63][238] * vector[63] +matrix[64][238] * vector[64] +matrix[65][238] * vector[65] +matrix[66][238] * vector[66] +matrix[67][238] * vector[67] +matrix[68][238] * vector[68] +matrix[69][238] * vector[69] +matrix[70][238] * vector[70] +matrix[71][238] * vector[71] +matrix[72][238] * vector[72] +matrix[73][238] * vector[73] +matrix[74][238] * vector[74] +matrix[75][238] * vector[75] +matrix[76][238] * vector[76] +matrix[77][238] * vector[77] +matrix[78][238] * vector[78] +matrix[79][238] * vector[79] +matrix[80][238] * vector[80] +matrix[81][238] * vector[81] +matrix[82][238] * vector[82] +matrix[83][238] * vector[83] +matrix[84][238] * vector[84] +matrix[85][238] * vector[85] +matrix[86][238] * vector[86] +matrix[87][238] * vector[87] +matrix[88][238] * vector[88] +matrix[89][238] * vector[89] +matrix[90][238] * vector[90] +matrix[91][238] * vector[91] +matrix[92][238] * vector[92] +matrix[93][238] * vector[93] +matrix[94][238] * vector[94] +matrix[95][238] * vector[95] +matrix[96][238] * vector[96] +matrix[97][238] * vector[97] +matrix[98][238] * vector[98] +matrix[99][238] * vector[99] +b[238];
assign result[239] = matrix[0][239] * vector[0] +matrix[1][239] * vector[1] +matrix[2][239] * vector[2] +matrix[3][239] * vector[3] +matrix[4][239] * vector[4] +matrix[5][239] * vector[5] +matrix[6][239] * vector[6] +matrix[7][239] * vector[7] +matrix[8][239] * vector[8] +matrix[9][239] * vector[9] +matrix[10][239] * vector[10] +matrix[11][239] * vector[11] +matrix[12][239] * vector[12] +matrix[13][239] * vector[13] +matrix[14][239] * vector[14] +matrix[15][239] * vector[15] +matrix[16][239] * vector[16] +matrix[17][239] * vector[17] +matrix[18][239] * vector[18] +matrix[19][239] * vector[19] +matrix[20][239] * vector[20] +matrix[21][239] * vector[21] +matrix[22][239] * vector[22] +matrix[23][239] * vector[23] +matrix[24][239] * vector[24] +matrix[25][239] * vector[25] +matrix[26][239] * vector[26] +matrix[27][239] * vector[27] +matrix[28][239] * vector[28] +matrix[29][239] * vector[29] +matrix[30][239] * vector[30] +matrix[31][239] * vector[31] +matrix[32][239] * vector[32] +matrix[33][239] * vector[33] +matrix[34][239] * vector[34] +matrix[35][239] * vector[35] +matrix[36][239] * vector[36] +matrix[37][239] * vector[37] +matrix[38][239] * vector[38] +matrix[39][239] * vector[39] +matrix[40][239] * vector[40] +matrix[41][239] * vector[41] +matrix[42][239] * vector[42] +matrix[43][239] * vector[43] +matrix[44][239] * vector[44] +matrix[45][239] * vector[45] +matrix[46][239] * vector[46] +matrix[47][239] * vector[47] +matrix[48][239] * vector[48] +matrix[49][239] * vector[49] +matrix[50][239] * vector[50] +matrix[51][239] * vector[51] +matrix[52][239] * vector[52] +matrix[53][239] * vector[53] +matrix[54][239] * vector[54] +matrix[55][239] * vector[55] +matrix[56][239] * vector[56] +matrix[57][239] * vector[57] +matrix[58][239] * vector[58] +matrix[59][239] * vector[59] +matrix[60][239] * vector[60] +matrix[61][239] * vector[61] +matrix[62][239] * vector[62] +matrix[63][239] * vector[63] +matrix[64][239] * vector[64] +matrix[65][239] * vector[65] +matrix[66][239] * vector[66] +matrix[67][239] * vector[67] +matrix[68][239] * vector[68] +matrix[69][239] * vector[69] +matrix[70][239] * vector[70] +matrix[71][239] * vector[71] +matrix[72][239] * vector[72] +matrix[73][239] * vector[73] +matrix[74][239] * vector[74] +matrix[75][239] * vector[75] +matrix[76][239] * vector[76] +matrix[77][239] * vector[77] +matrix[78][239] * vector[78] +matrix[79][239] * vector[79] +matrix[80][239] * vector[80] +matrix[81][239] * vector[81] +matrix[82][239] * vector[82] +matrix[83][239] * vector[83] +matrix[84][239] * vector[84] +matrix[85][239] * vector[85] +matrix[86][239] * vector[86] +matrix[87][239] * vector[87] +matrix[88][239] * vector[88] +matrix[89][239] * vector[89] +matrix[90][239] * vector[90] +matrix[91][239] * vector[91] +matrix[92][239] * vector[92] +matrix[93][239] * vector[93] +matrix[94][239] * vector[94] +matrix[95][239] * vector[95] +matrix[96][239] * vector[96] +matrix[97][239] * vector[97] +matrix[98][239] * vector[98] +matrix[99][239] * vector[99] +b[239];
assign result[240] = matrix[0][240] * vector[0] +matrix[1][240] * vector[1] +matrix[2][240] * vector[2] +matrix[3][240] * vector[3] +matrix[4][240] * vector[4] +matrix[5][240] * vector[5] +matrix[6][240] * vector[6] +matrix[7][240] * vector[7] +matrix[8][240] * vector[8] +matrix[9][240] * vector[9] +matrix[10][240] * vector[10] +matrix[11][240] * vector[11] +matrix[12][240] * vector[12] +matrix[13][240] * vector[13] +matrix[14][240] * vector[14] +matrix[15][240] * vector[15] +matrix[16][240] * vector[16] +matrix[17][240] * vector[17] +matrix[18][240] * vector[18] +matrix[19][240] * vector[19] +matrix[20][240] * vector[20] +matrix[21][240] * vector[21] +matrix[22][240] * vector[22] +matrix[23][240] * vector[23] +matrix[24][240] * vector[24] +matrix[25][240] * vector[25] +matrix[26][240] * vector[26] +matrix[27][240] * vector[27] +matrix[28][240] * vector[28] +matrix[29][240] * vector[29] +matrix[30][240] * vector[30] +matrix[31][240] * vector[31] +matrix[32][240] * vector[32] +matrix[33][240] * vector[33] +matrix[34][240] * vector[34] +matrix[35][240] * vector[35] +matrix[36][240] * vector[36] +matrix[37][240] * vector[37] +matrix[38][240] * vector[38] +matrix[39][240] * vector[39] +matrix[40][240] * vector[40] +matrix[41][240] * vector[41] +matrix[42][240] * vector[42] +matrix[43][240] * vector[43] +matrix[44][240] * vector[44] +matrix[45][240] * vector[45] +matrix[46][240] * vector[46] +matrix[47][240] * vector[47] +matrix[48][240] * vector[48] +matrix[49][240] * vector[49] +matrix[50][240] * vector[50] +matrix[51][240] * vector[51] +matrix[52][240] * vector[52] +matrix[53][240] * vector[53] +matrix[54][240] * vector[54] +matrix[55][240] * vector[55] +matrix[56][240] * vector[56] +matrix[57][240] * vector[57] +matrix[58][240] * vector[58] +matrix[59][240] * vector[59] +matrix[60][240] * vector[60] +matrix[61][240] * vector[61] +matrix[62][240] * vector[62] +matrix[63][240] * vector[63] +matrix[64][240] * vector[64] +matrix[65][240] * vector[65] +matrix[66][240] * vector[66] +matrix[67][240] * vector[67] +matrix[68][240] * vector[68] +matrix[69][240] * vector[69] +matrix[70][240] * vector[70] +matrix[71][240] * vector[71] +matrix[72][240] * vector[72] +matrix[73][240] * vector[73] +matrix[74][240] * vector[74] +matrix[75][240] * vector[75] +matrix[76][240] * vector[76] +matrix[77][240] * vector[77] +matrix[78][240] * vector[78] +matrix[79][240] * vector[79] +matrix[80][240] * vector[80] +matrix[81][240] * vector[81] +matrix[82][240] * vector[82] +matrix[83][240] * vector[83] +matrix[84][240] * vector[84] +matrix[85][240] * vector[85] +matrix[86][240] * vector[86] +matrix[87][240] * vector[87] +matrix[88][240] * vector[88] +matrix[89][240] * vector[89] +matrix[90][240] * vector[90] +matrix[91][240] * vector[91] +matrix[92][240] * vector[92] +matrix[93][240] * vector[93] +matrix[94][240] * vector[94] +matrix[95][240] * vector[95] +matrix[96][240] * vector[96] +matrix[97][240] * vector[97] +matrix[98][240] * vector[98] +matrix[99][240] * vector[99] +b[240];
assign result[241] = matrix[0][241] * vector[0] +matrix[1][241] * vector[1] +matrix[2][241] * vector[2] +matrix[3][241] * vector[3] +matrix[4][241] * vector[4] +matrix[5][241] * vector[5] +matrix[6][241] * vector[6] +matrix[7][241] * vector[7] +matrix[8][241] * vector[8] +matrix[9][241] * vector[9] +matrix[10][241] * vector[10] +matrix[11][241] * vector[11] +matrix[12][241] * vector[12] +matrix[13][241] * vector[13] +matrix[14][241] * vector[14] +matrix[15][241] * vector[15] +matrix[16][241] * vector[16] +matrix[17][241] * vector[17] +matrix[18][241] * vector[18] +matrix[19][241] * vector[19] +matrix[20][241] * vector[20] +matrix[21][241] * vector[21] +matrix[22][241] * vector[22] +matrix[23][241] * vector[23] +matrix[24][241] * vector[24] +matrix[25][241] * vector[25] +matrix[26][241] * vector[26] +matrix[27][241] * vector[27] +matrix[28][241] * vector[28] +matrix[29][241] * vector[29] +matrix[30][241] * vector[30] +matrix[31][241] * vector[31] +matrix[32][241] * vector[32] +matrix[33][241] * vector[33] +matrix[34][241] * vector[34] +matrix[35][241] * vector[35] +matrix[36][241] * vector[36] +matrix[37][241] * vector[37] +matrix[38][241] * vector[38] +matrix[39][241] * vector[39] +matrix[40][241] * vector[40] +matrix[41][241] * vector[41] +matrix[42][241] * vector[42] +matrix[43][241] * vector[43] +matrix[44][241] * vector[44] +matrix[45][241] * vector[45] +matrix[46][241] * vector[46] +matrix[47][241] * vector[47] +matrix[48][241] * vector[48] +matrix[49][241] * vector[49] +matrix[50][241] * vector[50] +matrix[51][241] * vector[51] +matrix[52][241] * vector[52] +matrix[53][241] * vector[53] +matrix[54][241] * vector[54] +matrix[55][241] * vector[55] +matrix[56][241] * vector[56] +matrix[57][241] * vector[57] +matrix[58][241] * vector[58] +matrix[59][241] * vector[59] +matrix[60][241] * vector[60] +matrix[61][241] * vector[61] +matrix[62][241] * vector[62] +matrix[63][241] * vector[63] +matrix[64][241] * vector[64] +matrix[65][241] * vector[65] +matrix[66][241] * vector[66] +matrix[67][241] * vector[67] +matrix[68][241] * vector[68] +matrix[69][241] * vector[69] +matrix[70][241] * vector[70] +matrix[71][241] * vector[71] +matrix[72][241] * vector[72] +matrix[73][241] * vector[73] +matrix[74][241] * vector[74] +matrix[75][241] * vector[75] +matrix[76][241] * vector[76] +matrix[77][241] * vector[77] +matrix[78][241] * vector[78] +matrix[79][241] * vector[79] +matrix[80][241] * vector[80] +matrix[81][241] * vector[81] +matrix[82][241] * vector[82] +matrix[83][241] * vector[83] +matrix[84][241] * vector[84] +matrix[85][241] * vector[85] +matrix[86][241] * vector[86] +matrix[87][241] * vector[87] +matrix[88][241] * vector[88] +matrix[89][241] * vector[89] +matrix[90][241] * vector[90] +matrix[91][241] * vector[91] +matrix[92][241] * vector[92] +matrix[93][241] * vector[93] +matrix[94][241] * vector[94] +matrix[95][241] * vector[95] +matrix[96][241] * vector[96] +matrix[97][241] * vector[97] +matrix[98][241] * vector[98] +matrix[99][241] * vector[99] +b[241];
assign result[242] = matrix[0][242] * vector[0] +matrix[1][242] * vector[1] +matrix[2][242] * vector[2] +matrix[3][242] * vector[3] +matrix[4][242] * vector[4] +matrix[5][242] * vector[5] +matrix[6][242] * vector[6] +matrix[7][242] * vector[7] +matrix[8][242] * vector[8] +matrix[9][242] * vector[9] +matrix[10][242] * vector[10] +matrix[11][242] * vector[11] +matrix[12][242] * vector[12] +matrix[13][242] * vector[13] +matrix[14][242] * vector[14] +matrix[15][242] * vector[15] +matrix[16][242] * vector[16] +matrix[17][242] * vector[17] +matrix[18][242] * vector[18] +matrix[19][242] * vector[19] +matrix[20][242] * vector[20] +matrix[21][242] * vector[21] +matrix[22][242] * vector[22] +matrix[23][242] * vector[23] +matrix[24][242] * vector[24] +matrix[25][242] * vector[25] +matrix[26][242] * vector[26] +matrix[27][242] * vector[27] +matrix[28][242] * vector[28] +matrix[29][242] * vector[29] +matrix[30][242] * vector[30] +matrix[31][242] * vector[31] +matrix[32][242] * vector[32] +matrix[33][242] * vector[33] +matrix[34][242] * vector[34] +matrix[35][242] * vector[35] +matrix[36][242] * vector[36] +matrix[37][242] * vector[37] +matrix[38][242] * vector[38] +matrix[39][242] * vector[39] +matrix[40][242] * vector[40] +matrix[41][242] * vector[41] +matrix[42][242] * vector[42] +matrix[43][242] * vector[43] +matrix[44][242] * vector[44] +matrix[45][242] * vector[45] +matrix[46][242] * vector[46] +matrix[47][242] * vector[47] +matrix[48][242] * vector[48] +matrix[49][242] * vector[49] +matrix[50][242] * vector[50] +matrix[51][242] * vector[51] +matrix[52][242] * vector[52] +matrix[53][242] * vector[53] +matrix[54][242] * vector[54] +matrix[55][242] * vector[55] +matrix[56][242] * vector[56] +matrix[57][242] * vector[57] +matrix[58][242] * vector[58] +matrix[59][242] * vector[59] +matrix[60][242] * vector[60] +matrix[61][242] * vector[61] +matrix[62][242] * vector[62] +matrix[63][242] * vector[63] +matrix[64][242] * vector[64] +matrix[65][242] * vector[65] +matrix[66][242] * vector[66] +matrix[67][242] * vector[67] +matrix[68][242] * vector[68] +matrix[69][242] * vector[69] +matrix[70][242] * vector[70] +matrix[71][242] * vector[71] +matrix[72][242] * vector[72] +matrix[73][242] * vector[73] +matrix[74][242] * vector[74] +matrix[75][242] * vector[75] +matrix[76][242] * vector[76] +matrix[77][242] * vector[77] +matrix[78][242] * vector[78] +matrix[79][242] * vector[79] +matrix[80][242] * vector[80] +matrix[81][242] * vector[81] +matrix[82][242] * vector[82] +matrix[83][242] * vector[83] +matrix[84][242] * vector[84] +matrix[85][242] * vector[85] +matrix[86][242] * vector[86] +matrix[87][242] * vector[87] +matrix[88][242] * vector[88] +matrix[89][242] * vector[89] +matrix[90][242] * vector[90] +matrix[91][242] * vector[91] +matrix[92][242] * vector[92] +matrix[93][242] * vector[93] +matrix[94][242] * vector[94] +matrix[95][242] * vector[95] +matrix[96][242] * vector[96] +matrix[97][242] * vector[97] +matrix[98][242] * vector[98] +matrix[99][242] * vector[99] +b[242];
assign result[243] = matrix[0][243] * vector[0] +matrix[1][243] * vector[1] +matrix[2][243] * vector[2] +matrix[3][243] * vector[3] +matrix[4][243] * vector[4] +matrix[5][243] * vector[5] +matrix[6][243] * vector[6] +matrix[7][243] * vector[7] +matrix[8][243] * vector[8] +matrix[9][243] * vector[9] +matrix[10][243] * vector[10] +matrix[11][243] * vector[11] +matrix[12][243] * vector[12] +matrix[13][243] * vector[13] +matrix[14][243] * vector[14] +matrix[15][243] * vector[15] +matrix[16][243] * vector[16] +matrix[17][243] * vector[17] +matrix[18][243] * vector[18] +matrix[19][243] * vector[19] +matrix[20][243] * vector[20] +matrix[21][243] * vector[21] +matrix[22][243] * vector[22] +matrix[23][243] * vector[23] +matrix[24][243] * vector[24] +matrix[25][243] * vector[25] +matrix[26][243] * vector[26] +matrix[27][243] * vector[27] +matrix[28][243] * vector[28] +matrix[29][243] * vector[29] +matrix[30][243] * vector[30] +matrix[31][243] * vector[31] +matrix[32][243] * vector[32] +matrix[33][243] * vector[33] +matrix[34][243] * vector[34] +matrix[35][243] * vector[35] +matrix[36][243] * vector[36] +matrix[37][243] * vector[37] +matrix[38][243] * vector[38] +matrix[39][243] * vector[39] +matrix[40][243] * vector[40] +matrix[41][243] * vector[41] +matrix[42][243] * vector[42] +matrix[43][243] * vector[43] +matrix[44][243] * vector[44] +matrix[45][243] * vector[45] +matrix[46][243] * vector[46] +matrix[47][243] * vector[47] +matrix[48][243] * vector[48] +matrix[49][243] * vector[49] +matrix[50][243] * vector[50] +matrix[51][243] * vector[51] +matrix[52][243] * vector[52] +matrix[53][243] * vector[53] +matrix[54][243] * vector[54] +matrix[55][243] * vector[55] +matrix[56][243] * vector[56] +matrix[57][243] * vector[57] +matrix[58][243] * vector[58] +matrix[59][243] * vector[59] +matrix[60][243] * vector[60] +matrix[61][243] * vector[61] +matrix[62][243] * vector[62] +matrix[63][243] * vector[63] +matrix[64][243] * vector[64] +matrix[65][243] * vector[65] +matrix[66][243] * vector[66] +matrix[67][243] * vector[67] +matrix[68][243] * vector[68] +matrix[69][243] * vector[69] +matrix[70][243] * vector[70] +matrix[71][243] * vector[71] +matrix[72][243] * vector[72] +matrix[73][243] * vector[73] +matrix[74][243] * vector[74] +matrix[75][243] * vector[75] +matrix[76][243] * vector[76] +matrix[77][243] * vector[77] +matrix[78][243] * vector[78] +matrix[79][243] * vector[79] +matrix[80][243] * vector[80] +matrix[81][243] * vector[81] +matrix[82][243] * vector[82] +matrix[83][243] * vector[83] +matrix[84][243] * vector[84] +matrix[85][243] * vector[85] +matrix[86][243] * vector[86] +matrix[87][243] * vector[87] +matrix[88][243] * vector[88] +matrix[89][243] * vector[89] +matrix[90][243] * vector[90] +matrix[91][243] * vector[91] +matrix[92][243] * vector[92] +matrix[93][243] * vector[93] +matrix[94][243] * vector[94] +matrix[95][243] * vector[95] +matrix[96][243] * vector[96] +matrix[97][243] * vector[97] +matrix[98][243] * vector[98] +matrix[99][243] * vector[99] +b[243];
assign result[244] = matrix[0][244] * vector[0] +matrix[1][244] * vector[1] +matrix[2][244] * vector[2] +matrix[3][244] * vector[3] +matrix[4][244] * vector[4] +matrix[5][244] * vector[5] +matrix[6][244] * vector[6] +matrix[7][244] * vector[7] +matrix[8][244] * vector[8] +matrix[9][244] * vector[9] +matrix[10][244] * vector[10] +matrix[11][244] * vector[11] +matrix[12][244] * vector[12] +matrix[13][244] * vector[13] +matrix[14][244] * vector[14] +matrix[15][244] * vector[15] +matrix[16][244] * vector[16] +matrix[17][244] * vector[17] +matrix[18][244] * vector[18] +matrix[19][244] * vector[19] +matrix[20][244] * vector[20] +matrix[21][244] * vector[21] +matrix[22][244] * vector[22] +matrix[23][244] * vector[23] +matrix[24][244] * vector[24] +matrix[25][244] * vector[25] +matrix[26][244] * vector[26] +matrix[27][244] * vector[27] +matrix[28][244] * vector[28] +matrix[29][244] * vector[29] +matrix[30][244] * vector[30] +matrix[31][244] * vector[31] +matrix[32][244] * vector[32] +matrix[33][244] * vector[33] +matrix[34][244] * vector[34] +matrix[35][244] * vector[35] +matrix[36][244] * vector[36] +matrix[37][244] * vector[37] +matrix[38][244] * vector[38] +matrix[39][244] * vector[39] +matrix[40][244] * vector[40] +matrix[41][244] * vector[41] +matrix[42][244] * vector[42] +matrix[43][244] * vector[43] +matrix[44][244] * vector[44] +matrix[45][244] * vector[45] +matrix[46][244] * vector[46] +matrix[47][244] * vector[47] +matrix[48][244] * vector[48] +matrix[49][244] * vector[49] +matrix[50][244] * vector[50] +matrix[51][244] * vector[51] +matrix[52][244] * vector[52] +matrix[53][244] * vector[53] +matrix[54][244] * vector[54] +matrix[55][244] * vector[55] +matrix[56][244] * vector[56] +matrix[57][244] * vector[57] +matrix[58][244] * vector[58] +matrix[59][244] * vector[59] +matrix[60][244] * vector[60] +matrix[61][244] * vector[61] +matrix[62][244] * vector[62] +matrix[63][244] * vector[63] +matrix[64][244] * vector[64] +matrix[65][244] * vector[65] +matrix[66][244] * vector[66] +matrix[67][244] * vector[67] +matrix[68][244] * vector[68] +matrix[69][244] * vector[69] +matrix[70][244] * vector[70] +matrix[71][244] * vector[71] +matrix[72][244] * vector[72] +matrix[73][244] * vector[73] +matrix[74][244] * vector[74] +matrix[75][244] * vector[75] +matrix[76][244] * vector[76] +matrix[77][244] * vector[77] +matrix[78][244] * vector[78] +matrix[79][244] * vector[79] +matrix[80][244] * vector[80] +matrix[81][244] * vector[81] +matrix[82][244] * vector[82] +matrix[83][244] * vector[83] +matrix[84][244] * vector[84] +matrix[85][244] * vector[85] +matrix[86][244] * vector[86] +matrix[87][244] * vector[87] +matrix[88][244] * vector[88] +matrix[89][244] * vector[89] +matrix[90][244] * vector[90] +matrix[91][244] * vector[91] +matrix[92][244] * vector[92] +matrix[93][244] * vector[93] +matrix[94][244] * vector[94] +matrix[95][244] * vector[95] +matrix[96][244] * vector[96] +matrix[97][244] * vector[97] +matrix[98][244] * vector[98] +matrix[99][244] * vector[99] +b[244];
assign result[245] = matrix[0][245] * vector[0] +matrix[1][245] * vector[1] +matrix[2][245] * vector[2] +matrix[3][245] * vector[3] +matrix[4][245] * vector[4] +matrix[5][245] * vector[5] +matrix[6][245] * vector[6] +matrix[7][245] * vector[7] +matrix[8][245] * vector[8] +matrix[9][245] * vector[9] +matrix[10][245] * vector[10] +matrix[11][245] * vector[11] +matrix[12][245] * vector[12] +matrix[13][245] * vector[13] +matrix[14][245] * vector[14] +matrix[15][245] * vector[15] +matrix[16][245] * vector[16] +matrix[17][245] * vector[17] +matrix[18][245] * vector[18] +matrix[19][245] * vector[19] +matrix[20][245] * vector[20] +matrix[21][245] * vector[21] +matrix[22][245] * vector[22] +matrix[23][245] * vector[23] +matrix[24][245] * vector[24] +matrix[25][245] * vector[25] +matrix[26][245] * vector[26] +matrix[27][245] * vector[27] +matrix[28][245] * vector[28] +matrix[29][245] * vector[29] +matrix[30][245] * vector[30] +matrix[31][245] * vector[31] +matrix[32][245] * vector[32] +matrix[33][245] * vector[33] +matrix[34][245] * vector[34] +matrix[35][245] * vector[35] +matrix[36][245] * vector[36] +matrix[37][245] * vector[37] +matrix[38][245] * vector[38] +matrix[39][245] * vector[39] +matrix[40][245] * vector[40] +matrix[41][245] * vector[41] +matrix[42][245] * vector[42] +matrix[43][245] * vector[43] +matrix[44][245] * vector[44] +matrix[45][245] * vector[45] +matrix[46][245] * vector[46] +matrix[47][245] * vector[47] +matrix[48][245] * vector[48] +matrix[49][245] * vector[49] +matrix[50][245] * vector[50] +matrix[51][245] * vector[51] +matrix[52][245] * vector[52] +matrix[53][245] * vector[53] +matrix[54][245] * vector[54] +matrix[55][245] * vector[55] +matrix[56][245] * vector[56] +matrix[57][245] * vector[57] +matrix[58][245] * vector[58] +matrix[59][245] * vector[59] +matrix[60][245] * vector[60] +matrix[61][245] * vector[61] +matrix[62][245] * vector[62] +matrix[63][245] * vector[63] +matrix[64][245] * vector[64] +matrix[65][245] * vector[65] +matrix[66][245] * vector[66] +matrix[67][245] * vector[67] +matrix[68][245] * vector[68] +matrix[69][245] * vector[69] +matrix[70][245] * vector[70] +matrix[71][245] * vector[71] +matrix[72][245] * vector[72] +matrix[73][245] * vector[73] +matrix[74][245] * vector[74] +matrix[75][245] * vector[75] +matrix[76][245] * vector[76] +matrix[77][245] * vector[77] +matrix[78][245] * vector[78] +matrix[79][245] * vector[79] +matrix[80][245] * vector[80] +matrix[81][245] * vector[81] +matrix[82][245] * vector[82] +matrix[83][245] * vector[83] +matrix[84][245] * vector[84] +matrix[85][245] * vector[85] +matrix[86][245] * vector[86] +matrix[87][245] * vector[87] +matrix[88][245] * vector[88] +matrix[89][245] * vector[89] +matrix[90][245] * vector[90] +matrix[91][245] * vector[91] +matrix[92][245] * vector[92] +matrix[93][245] * vector[93] +matrix[94][245] * vector[94] +matrix[95][245] * vector[95] +matrix[96][245] * vector[96] +matrix[97][245] * vector[97] +matrix[98][245] * vector[98] +matrix[99][245] * vector[99] +b[245];
assign result[246] = matrix[0][246] * vector[0] +matrix[1][246] * vector[1] +matrix[2][246] * vector[2] +matrix[3][246] * vector[3] +matrix[4][246] * vector[4] +matrix[5][246] * vector[5] +matrix[6][246] * vector[6] +matrix[7][246] * vector[7] +matrix[8][246] * vector[8] +matrix[9][246] * vector[9] +matrix[10][246] * vector[10] +matrix[11][246] * vector[11] +matrix[12][246] * vector[12] +matrix[13][246] * vector[13] +matrix[14][246] * vector[14] +matrix[15][246] * vector[15] +matrix[16][246] * vector[16] +matrix[17][246] * vector[17] +matrix[18][246] * vector[18] +matrix[19][246] * vector[19] +matrix[20][246] * vector[20] +matrix[21][246] * vector[21] +matrix[22][246] * vector[22] +matrix[23][246] * vector[23] +matrix[24][246] * vector[24] +matrix[25][246] * vector[25] +matrix[26][246] * vector[26] +matrix[27][246] * vector[27] +matrix[28][246] * vector[28] +matrix[29][246] * vector[29] +matrix[30][246] * vector[30] +matrix[31][246] * vector[31] +matrix[32][246] * vector[32] +matrix[33][246] * vector[33] +matrix[34][246] * vector[34] +matrix[35][246] * vector[35] +matrix[36][246] * vector[36] +matrix[37][246] * vector[37] +matrix[38][246] * vector[38] +matrix[39][246] * vector[39] +matrix[40][246] * vector[40] +matrix[41][246] * vector[41] +matrix[42][246] * vector[42] +matrix[43][246] * vector[43] +matrix[44][246] * vector[44] +matrix[45][246] * vector[45] +matrix[46][246] * vector[46] +matrix[47][246] * vector[47] +matrix[48][246] * vector[48] +matrix[49][246] * vector[49] +matrix[50][246] * vector[50] +matrix[51][246] * vector[51] +matrix[52][246] * vector[52] +matrix[53][246] * vector[53] +matrix[54][246] * vector[54] +matrix[55][246] * vector[55] +matrix[56][246] * vector[56] +matrix[57][246] * vector[57] +matrix[58][246] * vector[58] +matrix[59][246] * vector[59] +matrix[60][246] * vector[60] +matrix[61][246] * vector[61] +matrix[62][246] * vector[62] +matrix[63][246] * vector[63] +matrix[64][246] * vector[64] +matrix[65][246] * vector[65] +matrix[66][246] * vector[66] +matrix[67][246] * vector[67] +matrix[68][246] * vector[68] +matrix[69][246] * vector[69] +matrix[70][246] * vector[70] +matrix[71][246] * vector[71] +matrix[72][246] * vector[72] +matrix[73][246] * vector[73] +matrix[74][246] * vector[74] +matrix[75][246] * vector[75] +matrix[76][246] * vector[76] +matrix[77][246] * vector[77] +matrix[78][246] * vector[78] +matrix[79][246] * vector[79] +matrix[80][246] * vector[80] +matrix[81][246] * vector[81] +matrix[82][246] * vector[82] +matrix[83][246] * vector[83] +matrix[84][246] * vector[84] +matrix[85][246] * vector[85] +matrix[86][246] * vector[86] +matrix[87][246] * vector[87] +matrix[88][246] * vector[88] +matrix[89][246] * vector[89] +matrix[90][246] * vector[90] +matrix[91][246] * vector[91] +matrix[92][246] * vector[92] +matrix[93][246] * vector[93] +matrix[94][246] * vector[94] +matrix[95][246] * vector[95] +matrix[96][246] * vector[96] +matrix[97][246] * vector[97] +matrix[98][246] * vector[98] +matrix[99][246] * vector[99] +b[246];
assign result[247] = matrix[0][247] * vector[0] +matrix[1][247] * vector[1] +matrix[2][247] * vector[2] +matrix[3][247] * vector[3] +matrix[4][247] * vector[4] +matrix[5][247] * vector[5] +matrix[6][247] * vector[6] +matrix[7][247] * vector[7] +matrix[8][247] * vector[8] +matrix[9][247] * vector[9] +matrix[10][247] * vector[10] +matrix[11][247] * vector[11] +matrix[12][247] * vector[12] +matrix[13][247] * vector[13] +matrix[14][247] * vector[14] +matrix[15][247] * vector[15] +matrix[16][247] * vector[16] +matrix[17][247] * vector[17] +matrix[18][247] * vector[18] +matrix[19][247] * vector[19] +matrix[20][247] * vector[20] +matrix[21][247] * vector[21] +matrix[22][247] * vector[22] +matrix[23][247] * vector[23] +matrix[24][247] * vector[24] +matrix[25][247] * vector[25] +matrix[26][247] * vector[26] +matrix[27][247] * vector[27] +matrix[28][247] * vector[28] +matrix[29][247] * vector[29] +matrix[30][247] * vector[30] +matrix[31][247] * vector[31] +matrix[32][247] * vector[32] +matrix[33][247] * vector[33] +matrix[34][247] * vector[34] +matrix[35][247] * vector[35] +matrix[36][247] * vector[36] +matrix[37][247] * vector[37] +matrix[38][247] * vector[38] +matrix[39][247] * vector[39] +matrix[40][247] * vector[40] +matrix[41][247] * vector[41] +matrix[42][247] * vector[42] +matrix[43][247] * vector[43] +matrix[44][247] * vector[44] +matrix[45][247] * vector[45] +matrix[46][247] * vector[46] +matrix[47][247] * vector[47] +matrix[48][247] * vector[48] +matrix[49][247] * vector[49] +matrix[50][247] * vector[50] +matrix[51][247] * vector[51] +matrix[52][247] * vector[52] +matrix[53][247] * vector[53] +matrix[54][247] * vector[54] +matrix[55][247] * vector[55] +matrix[56][247] * vector[56] +matrix[57][247] * vector[57] +matrix[58][247] * vector[58] +matrix[59][247] * vector[59] +matrix[60][247] * vector[60] +matrix[61][247] * vector[61] +matrix[62][247] * vector[62] +matrix[63][247] * vector[63] +matrix[64][247] * vector[64] +matrix[65][247] * vector[65] +matrix[66][247] * vector[66] +matrix[67][247] * vector[67] +matrix[68][247] * vector[68] +matrix[69][247] * vector[69] +matrix[70][247] * vector[70] +matrix[71][247] * vector[71] +matrix[72][247] * vector[72] +matrix[73][247] * vector[73] +matrix[74][247] * vector[74] +matrix[75][247] * vector[75] +matrix[76][247] * vector[76] +matrix[77][247] * vector[77] +matrix[78][247] * vector[78] +matrix[79][247] * vector[79] +matrix[80][247] * vector[80] +matrix[81][247] * vector[81] +matrix[82][247] * vector[82] +matrix[83][247] * vector[83] +matrix[84][247] * vector[84] +matrix[85][247] * vector[85] +matrix[86][247] * vector[86] +matrix[87][247] * vector[87] +matrix[88][247] * vector[88] +matrix[89][247] * vector[89] +matrix[90][247] * vector[90] +matrix[91][247] * vector[91] +matrix[92][247] * vector[92] +matrix[93][247] * vector[93] +matrix[94][247] * vector[94] +matrix[95][247] * vector[95] +matrix[96][247] * vector[96] +matrix[97][247] * vector[97] +matrix[98][247] * vector[98] +matrix[99][247] * vector[99] +b[247];
assign result[248] = matrix[0][248] * vector[0] +matrix[1][248] * vector[1] +matrix[2][248] * vector[2] +matrix[3][248] * vector[3] +matrix[4][248] * vector[4] +matrix[5][248] * vector[5] +matrix[6][248] * vector[6] +matrix[7][248] * vector[7] +matrix[8][248] * vector[8] +matrix[9][248] * vector[9] +matrix[10][248] * vector[10] +matrix[11][248] * vector[11] +matrix[12][248] * vector[12] +matrix[13][248] * vector[13] +matrix[14][248] * vector[14] +matrix[15][248] * vector[15] +matrix[16][248] * vector[16] +matrix[17][248] * vector[17] +matrix[18][248] * vector[18] +matrix[19][248] * vector[19] +matrix[20][248] * vector[20] +matrix[21][248] * vector[21] +matrix[22][248] * vector[22] +matrix[23][248] * vector[23] +matrix[24][248] * vector[24] +matrix[25][248] * vector[25] +matrix[26][248] * vector[26] +matrix[27][248] * vector[27] +matrix[28][248] * vector[28] +matrix[29][248] * vector[29] +matrix[30][248] * vector[30] +matrix[31][248] * vector[31] +matrix[32][248] * vector[32] +matrix[33][248] * vector[33] +matrix[34][248] * vector[34] +matrix[35][248] * vector[35] +matrix[36][248] * vector[36] +matrix[37][248] * vector[37] +matrix[38][248] * vector[38] +matrix[39][248] * vector[39] +matrix[40][248] * vector[40] +matrix[41][248] * vector[41] +matrix[42][248] * vector[42] +matrix[43][248] * vector[43] +matrix[44][248] * vector[44] +matrix[45][248] * vector[45] +matrix[46][248] * vector[46] +matrix[47][248] * vector[47] +matrix[48][248] * vector[48] +matrix[49][248] * vector[49] +matrix[50][248] * vector[50] +matrix[51][248] * vector[51] +matrix[52][248] * vector[52] +matrix[53][248] * vector[53] +matrix[54][248] * vector[54] +matrix[55][248] * vector[55] +matrix[56][248] * vector[56] +matrix[57][248] * vector[57] +matrix[58][248] * vector[58] +matrix[59][248] * vector[59] +matrix[60][248] * vector[60] +matrix[61][248] * vector[61] +matrix[62][248] * vector[62] +matrix[63][248] * vector[63] +matrix[64][248] * vector[64] +matrix[65][248] * vector[65] +matrix[66][248] * vector[66] +matrix[67][248] * vector[67] +matrix[68][248] * vector[68] +matrix[69][248] * vector[69] +matrix[70][248] * vector[70] +matrix[71][248] * vector[71] +matrix[72][248] * vector[72] +matrix[73][248] * vector[73] +matrix[74][248] * vector[74] +matrix[75][248] * vector[75] +matrix[76][248] * vector[76] +matrix[77][248] * vector[77] +matrix[78][248] * vector[78] +matrix[79][248] * vector[79] +matrix[80][248] * vector[80] +matrix[81][248] * vector[81] +matrix[82][248] * vector[82] +matrix[83][248] * vector[83] +matrix[84][248] * vector[84] +matrix[85][248] * vector[85] +matrix[86][248] * vector[86] +matrix[87][248] * vector[87] +matrix[88][248] * vector[88] +matrix[89][248] * vector[89] +matrix[90][248] * vector[90] +matrix[91][248] * vector[91] +matrix[92][248] * vector[92] +matrix[93][248] * vector[93] +matrix[94][248] * vector[94] +matrix[95][248] * vector[95] +matrix[96][248] * vector[96] +matrix[97][248] * vector[97] +matrix[98][248] * vector[98] +matrix[99][248] * vector[99] +b[248];
assign result[249] = matrix[0][249] * vector[0] +matrix[1][249] * vector[1] +matrix[2][249] * vector[2] +matrix[3][249] * vector[3] +matrix[4][249] * vector[4] +matrix[5][249] * vector[5] +matrix[6][249] * vector[6] +matrix[7][249] * vector[7] +matrix[8][249] * vector[8] +matrix[9][249] * vector[9] +matrix[10][249] * vector[10] +matrix[11][249] * vector[11] +matrix[12][249] * vector[12] +matrix[13][249] * vector[13] +matrix[14][249] * vector[14] +matrix[15][249] * vector[15] +matrix[16][249] * vector[16] +matrix[17][249] * vector[17] +matrix[18][249] * vector[18] +matrix[19][249] * vector[19] +matrix[20][249] * vector[20] +matrix[21][249] * vector[21] +matrix[22][249] * vector[22] +matrix[23][249] * vector[23] +matrix[24][249] * vector[24] +matrix[25][249] * vector[25] +matrix[26][249] * vector[26] +matrix[27][249] * vector[27] +matrix[28][249] * vector[28] +matrix[29][249] * vector[29] +matrix[30][249] * vector[30] +matrix[31][249] * vector[31] +matrix[32][249] * vector[32] +matrix[33][249] * vector[33] +matrix[34][249] * vector[34] +matrix[35][249] * vector[35] +matrix[36][249] * vector[36] +matrix[37][249] * vector[37] +matrix[38][249] * vector[38] +matrix[39][249] * vector[39] +matrix[40][249] * vector[40] +matrix[41][249] * vector[41] +matrix[42][249] * vector[42] +matrix[43][249] * vector[43] +matrix[44][249] * vector[44] +matrix[45][249] * vector[45] +matrix[46][249] * vector[46] +matrix[47][249] * vector[47] +matrix[48][249] * vector[48] +matrix[49][249] * vector[49] +matrix[50][249] * vector[50] +matrix[51][249] * vector[51] +matrix[52][249] * vector[52] +matrix[53][249] * vector[53] +matrix[54][249] * vector[54] +matrix[55][249] * vector[55] +matrix[56][249] * vector[56] +matrix[57][249] * vector[57] +matrix[58][249] * vector[58] +matrix[59][249] * vector[59] +matrix[60][249] * vector[60] +matrix[61][249] * vector[61] +matrix[62][249] * vector[62] +matrix[63][249] * vector[63] +matrix[64][249] * vector[64] +matrix[65][249] * vector[65] +matrix[66][249] * vector[66] +matrix[67][249] * vector[67] +matrix[68][249] * vector[68] +matrix[69][249] * vector[69] +matrix[70][249] * vector[70] +matrix[71][249] * vector[71] +matrix[72][249] * vector[72] +matrix[73][249] * vector[73] +matrix[74][249] * vector[74] +matrix[75][249] * vector[75] +matrix[76][249] * vector[76] +matrix[77][249] * vector[77] +matrix[78][249] * vector[78] +matrix[79][249] * vector[79] +matrix[80][249] * vector[80] +matrix[81][249] * vector[81] +matrix[82][249] * vector[82] +matrix[83][249] * vector[83] +matrix[84][249] * vector[84] +matrix[85][249] * vector[85] +matrix[86][249] * vector[86] +matrix[87][249] * vector[87] +matrix[88][249] * vector[88] +matrix[89][249] * vector[89] +matrix[90][249] * vector[90] +matrix[91][249] * vector[91] +matrix[92][249] * vector[92] +matrix[93][249] * vector[93] +matrix[94][249] * vector[94] +matrix[95][249] * vector[95] +matrix[96][249] * vector[96] +matrix[97][249] * vector[97] +matrix[98][249] * vector[98] +matrix[99][249] * vector[99] +b[249];
assign result[250] = matrix[0][250] * vector[0] +matrix[1][250] * vector[1] +matrix[2][250] * vector[2] +matrix[3][250] * vector[3] +matrix[4][250] * vector[4] +matrix[5][250] * vector[5] +matrix[6][250] * vector[6] +matrix[7][250] * vector[7] +matrix[8][250] * vector[8] +matrix[9][250] * vector[9] +matrix[10][250] * vector[10] +matrix[11][250] * vector[11] +matrix[12][250] * vector[12] +matrix[13][250] * vector[13] +matrix[14][250] * vector[14] +matrix[15][250] * vector[15] +matrix[16][250] * vector[16] +matrix[17][250] * vector[17] +matrix[18][250] * vector[18] +matrix[19][250] * vector[19] +matrix[20][250] * vector[20] +matrix[21][250] * vector[21] +matrix[22][250] * vector[22] +matrix[23][250] * vector[23] +matrix[24][250] * vector[24] +matrix[25][250] * vector[25] +matrix[26][250] * vector[26] +matrix[27][250] * vector[27] +matrix[28][250] * vector[28] +matrix[29][250] * vector[29] +matrix[30][250] * vector[30] +matrix[31][250] * vector[31] +matrix[32][250] * vector[32] +matrix[33][250] * vector[33] +matrix[34][250] * vector[34] +matrix[35][250] * vector[35] +matrix[36][250] * vector[36] +matrix[37][250] * vector[37] +matrix[38][250] * vector[38] +matrix[39][250] * vector[39] +matrix[40][250] * vector[40] +matrix[41][250] * vector[41] +matrix[42][250] * vector[42] +matrix[43][250] * vector[43] +matrix[44][250] * vector[44] +matrix[45][250] * vector[45] +matrix[46][250] * vector[46] +matrix[47][250] * vector[47] +matrix[48][250] * vector[48] +matrix[49][250] * vector[49] +matrix[50][250] * vector[50] +matrix[51][250] * vector[51] +matrix[52][250] * vector[52] +matrix[53][250] * vector[53] +matrix[54][250] * vector[54] +matrix[55][250] * vector[55] +matrix[56][250] * vector[56] +matrix[57][250] * vector[57] +matrix[58][250] * vector[58] +matrix[59][250] * vector[59] +matrix[60][250] * vector[60] +matrix[61][250] * vector[61] +matrix[62][250] * vector[62] +matrix[63][250] * vector[63] +matrix[64][250] * vector[64] +matrix[65][250] * vector[65] +matrix[66][250] * vector[66] +matrix[67][250] * vector[67] +matrix[68][250] * vector[68] +matrix[69][250] * vector[69] +matrix[70][250] * vector[70] +matrix[71][250] * vector[71] +matrix[72][250] * vector[72] +matrix[73][250] * vector[73] +matrix[74][250] * vector[74] +matrix[75][250] * vector[75] +matrix[76][250] * vector[76] +matrix[77][250] * vector[77] +matrix[78][250] * vector[78] +matrix[79][250] * vector[79] +matrix[80][250] * vector[80] +matrix[81][250] * vector[81] +matrix[82][250] * vector[82] +matrix[83][250] * vector[83] +matrix[84][250] * vector[84] +matrix[85][250] * vector[85] +matrix[86][250] * vector[86] +matrix[87][250] * vector[87] +matrix[88][250] * vector[88] +matrix[89][250] * vector[89] +matrix[90][250] * vector[90] +matrix[91][250] * vector[91] +matrix[92][250] * vector[92] +matrix[93][250] * vector[93] +matrix[94][250] * vector[94] +matrix[95][250] * vector[95] +matrix[96][250] * vector[96] +matrix[97][250] * vector[97] +matrix[98][250] * vector[98] +matrix[99][250] * vector[99] +b[250];
assign result[251] = matrix[0][251] * vector[0] +matrix[1][251] * vector[1] +matrix[2][251] * vector[2] +matrix[3][251] * vector[3] +matrix[4][251] * vector[4] +matrix[5][251] * vector[5] +matrix[6][251] * vector[6] +matrix[7][251] * vector[7] +matrix[8][251] * vector[8] +matrix[9][251] * vector[9] +matrix[10][251] * vector[10] +matrix[11][251] * vector[11] +matrix[12][251] * vector[12] +matrix[13][251] * vector[13] +matrix[14][251] * vector[14] +matrix[15][251] * vector[15] +matrix[16][251] * vector[16] +matrix[17][251] * vector[17] +matrix[18][251] * vector[18] +matrix[19][251] * vector[19] +matrix[20][251] * vector[20] +matrix[21][251] * vector[21] +matrix[22][251] * vector[22] +matrix[23][251] * vector[23] +matrix[24][251] * vector[24] +matrix[25][251] * vector[25] +matrix[26][251] * vector[26] +matrix[27][251] * vector[27] +matrix[28][251] * vector[28] +matrix[29][251] * vector[29] +matrix[30][251] * vector[30] +matrix[31][251] * vector[31] +matrix[32][251] * vector[32] +matrix[33][251] * vector[33] +matrix[34][251] * vector[34] +matrix[35][251] * vector[35] +matrix[36][251] * vector[36] +matrix[37][251] * vector[37] +matrix[38][251] * vector[38] +matrix[39][251] * vector[39] +matrix[40][251] * vector[40] +matrix[41][251] * vector[41] +matrix[42][251] * vector[42] +matrix[43][251] * vector[43] +matrix[44][251] * vector[44] +matrix[45][251] * vector[45] +matrix[46][251] * vector[46] +matrix[47][251] * vector[47] +matrix[48][251] * vector[48] +matrix[49][251] * vector[49] +matrix[50][251] * vector[50] +matrix[51][251] * vector[51] +matrix[52][251] * vector[52] +matrix[53][251] * vector[53] +matrix[54][251] * vector[54] +matrix[55][251] * vector[55] +matrix[56][251] * vector[56] +matrix[57][251] * vector[57] +matrix[58][251] * vector[58] +matrix[59][251] * vector[59] +matrix[60][251] * vector[60] +matrix[61][251] * vector[61] +matrix[62][251] * vector[62] +matrix[63][251] * vector[63] +matrix[64][251] * vector[64] +matrix[65][251] * vector[65] +matrix[66][251] * vector[66] +matrix[67][251] * vector[67] +matrix[68][251] * vector[68] +matrix[69][251] * vector[69] +matrix[70][251] * vector[70] +matrix[71][251] * vector[71] +matrix[72][251] * vector[72] +matrix[73][251] * vector[73] +matrix[74][251] * vector[74] +matrix[75][251] * vector[75] +matrix[76][251] * vector[76] +matrix[77][251] * vector[77] +matrix[78][251] * vector[78] +matrix[79][251] * vector[79] +matrix[80][251] * vector[80] +matrix[81][251] * vector[81] +matrix[82][251] * vector[82] +matrix[83][251] * vector[83] +matrix[84][251] * vector[84] +matrix[85][251] * vector[85] +matrix[86][251] * vector[86] +matrix[87][251] * vector[87] +matrix[88][251] * vector[88] +matrix[89][251] * vector[89] +matrix[90][251] * vector[90] +matrix[91][251] * vector[91] +matrix[92][251] * vector[92] +matrix[93][251] * vector[93] +matrix[94][251] * vector[94] +matrix[95][251] * vector[95] +matrix[96][251] * vector[96] +matrix[97][251] * vector[97] +matrix[98][251] * vector[98] +matrix[99][251] * vector[99] +b[251];
assign result[252] = matrix[0][252] * vector[0] +matrix[1][252] * vector[1] +matrix[2][252] * vector[2] +matrix[3][252] * vector[3] +matrix[4][252] * vector[4] +matrix[5][252] * vector[5] +matrix[6][252] * vector[6] +matrix[7][252] * vector[7] +matrix[8][252] * vector[8] +matrix[9][252] * vector[9] +matrix[10][252] * vector[10] +matrix[11][252] * vector[11] +matrix[12][252] * vector[12] +matrix[13][252] * vector[13] +matrix[14][252] * vector[14] +matrix[15][252] * vector[15] +matrix[16][252] * vector[16] +matrix[17][252] * vector[17] +matrix[18][252] * vector[18] +matrix[19][252] * vector[19] +matrix[20][252] * vector[20] +matrix[21][252] * vector[21] +matrix[22][252] * vector[22] +matrix[23][252] * vector[23] +matrix[24][252] * vector[24] +matrix[25][252] * vector[25] +matrix[26][252] * vector[26] +matrix[27][252] * vector[27] +matrix[28][252] * vector[28] +matrix[29][252] * vector[29] +matrix[30][252] * vector[30] +matrix[31][252] * vector[31] +matrix[32][252] * vector[32] +matrix[33][252] * vector[33] +matrix[34][252] * vector[34] +matrix[35][252] * vector[35] +matrix[36][252] * vector[36] +matrix[37][252] * vector[37] +matrix[38][252] * vector[38] +matrix[39][252] * vector[39] +matrix[40][252] * vector[40] +matrix[41][252] * vector[41] +matrix[42][252] * vector[42] +matrix[43][252] * vector[43] +matrix[44][252] * vector[44] +matrix[45][252] * vector[45] +matrix[46][252] * vector[46] +matrix[47][252] * vector[47] +matrix[48][252] * vector[48] +matrix[49][252] * vector[49] +matrix[50][252] * vector[50] +matrix[51][252] * vector[51] +matrix[52][252] * vector[52] +matrix[53][252] * vector[53] +matrix[54][252] * vector[54] +matrix[55][252] * vector[55] +matrix[56][252] * vector[56] +matrix[57][252] * vector[57] +matrix[58][252] * vector[58] +matrix[59][252] * vector[59] +matrix[60][252] * vector[60] +matrix[61][252] * vector[61] +matrix[62][252] * vector[62] +matrix[63][252] * vector[63] +matrix[64][252] * vector[64] +matrix[65][252] * vector[65] +matrix[66][252] * vector[66] +matrix[67][252] * vector[67] +matrix[68][252] * vector[68] +matrix[69][252] * vector[69] +matrix[70][252] * vector[70] +matrix[71][252] * vector[71] +matrix[72][252] * vector[72] +matrix[73][252] * vector[73] +matrix[74][252] * vector[74] +matrix[75][252] * vector[75] +matrix[76][252] * vector[76] +matrix[77][252] * vector[77] +matrix[78][252] * vector[78] +matrix[79][252] * vector[79] +matrix[80][252] * vector[80] +matrix[81][252] * vector[81] +matrix[82][252] * vector[82] +matrix[83][252] * vector[83] +matrix[84][252] * vector[84] +matrix[85][252] * vector[85] +matrix[86][252] * vector[86] +matrix[87][252] * vector[87] +matrix[88][252] * vector[88] +matrix[89][252] * vector[89] +matrix[90][252] * vector[90] +matrix[91][252] * vector[91] +matrix[92][252] * vector[92] +matrix[93][252] * vector[93] +matrix[94][252] * vector[94] +matrix[95][252] * vector[95] +matrix[96][252] * vector[96] +matrix[97][252] * vector[97] +matrix[98][252] * vector[98] +matrix[99][252] * vector[99] +b[252];
assign result[253] = matrix[0][253] * vector[0] +matrix[1][253] * vector[1] +matrix[2][253] * vector[2] +matrix[3][253] * vector[3] +matrix[4][253] * vector[4] +matrix[5][253] * vector[5] +matrix[6][253] * vector[6] +matrix[7][253] * vector[7] +matrix[8][253] * vector[8] +matrix[9][253] * vector[9] +matrix[10][253] * vector[10] +matrix[11][253] * vector[11] +matrix[12][253] * vector[12] +matrix[13][253] * vector[13] +matrix[14][253] * vector[14] +matrix[15][253] * vector[15] +matrix[16][253] * vector[16] +matrix[17][253] * vector[17] +matrix[18][253] * vector[18] +matrix[19][253] * vector[19] +matrix[20][253] * vector[20] +matrix[21][253] * vector[21] +matrix[22][253] * vector[22] +matrix[23][253] * vector[23] +matrix[24][253] * vector[24] +matrix[25][253] * vector[25] +matrix[26][253] * vector[26] +matrix[27][253] * vector[27] +matrix[28][253] * vector[28] +matrix[29][253] * vector[29] +matrix[30][253] * vector[30] +matrix[31][253] * vector[31] +matrix[32][253] * vector[32] +matrix[33][253] * vector[33] +matrix[34][253] * vector[34] +matrix[35][253] * vector[35] +matrix[36][253] * vector[36] +matrix[37][253] * vector[37] +matrix[38][253] * vector[38] +matrix[39][253] * vector[39] +matrix[40][253] * vector[40] +matrix[41][253] * vector[41] +matrix[42][253] * vector[42] +matrix[43][253] * vector[43] +matrix[44][253] * vector[44] +matrix[45][253] * vector[45] +matrix[46][253] * vector[46] +matrix[47][253] * vector[47] +matrix[48][253] * vector[48] +matrix[49][253] * vector[49] +matrix[50][253] * vector[50] +matrix[51][253] * vector[51] +matrix[52][253] * vector[52] +matrix[53][253] * vector[53] +matrix[54][253] * vector[54] +matrix[55][253] * vector[55] +matrix[56][253] * vector[56] +matrix[57][253] * vector[57] +matrix[58][253] * vector[58] +matrix[59][253] * vector[59] +matrix[60][253] * vector[60] +matrix[61][253] * vector[61] +matrix[62][253] * vector[62] +matrix[63][253] * vector[63] +matrix[64][253] * vector[64] +matrix[65][253] * vector[65] +matrix[66][253] * vector[66] +matrix[67][253] * vector[67] +matrix[68][253] * vector[68] +matrix[69][253] * vector[69] +matrix[70][253] * vector[70] +matrix[71][253] * vector[71] +matrix[72][253] * vector[72] +matrix[73][253] * vector[73] +matrix[74][253] * vector[74] +matrix[75][253] * vector[75] +matrix[76][253] * vector[76] +matrix[77][253] * vector[77] +matrix[78][253] * vector[78] +matrix[79][253] * vector[79] +matrix[80][253] * vector[80] +matrix[81][253] * vector[81] +matrix[82][253] * vector[82] +matrix[83][253] * vector[83] +matrix[84][253] * vector[84] +matrix[85][253] * vector[85] +matrix[86][253] * vector[86] +matrix[87][253] * vector[87] +matrix[88][253] * vector[88] +matrix[89][253] * vector[89] +matrix[90][253] * vector[90] +matrix[91][253] * vector[91] +matrix[92][253] * vector[92] +matrix[93][253] * vector[93] +matrix[94][253] * vector[94] +matrix[95][253] * vector[95] +matrix[96][253] * vector[96] +matrix[97][253] * vector[97] +matrix[98][253] * vector[98] +matrix[99][253] * vector[99] +b[253];
assign result[254] = matrix[0][254] * vector[0] +matrix[1][254] * vector[1] +matrix[2][254] * vector[2] +matrix[3][254] * vector[3] +matrix[4][254] * vector[4] +matrix[5][254] * vector[5] +matrix[6][254] * vector[6] +matrix[7][254] * vector[7] +matrix[8][254] * vector[8] +matrix[9][254] * vector[9] +matrix[10][254] * vector[10] +matrix[11][254] * vector[11] +matrix[12][254] * vector[12] +matrix[13][254] * vector[13] +matrix[14][254] * vector[14] +matrix[15][254] * vector[15] +matrix[16][254] * vector[16] +matrix[17][254] * vector[17] +matrix[18][254] * vector[18] +matrix[19][254] * vector[19] +matrix[20][254] * vector[20] +matrix[21][254] * vector[21] +matrix[22][254] * vector[22] +matrix[23][254] * vector[23] +matrix[24][254] * vector[24] +matrix[25][254] * vector[25] +matrix[26][254] * vector[26] +matrix[27][254] * vector[27] +matrix[28][254] * vector[28] +matrix[29][254] * vector[29] +matrix[30][254] * vector[30] +matrix[31][254] * vector[31] +matrix[32][254] * vector[32] +matrix[33][254] * vector[33] +matrix[34][254] * vector[34] +matrix[35][254] * vector[35] +matrix[36][254] * vector[36] +matrix[37][254] * vector[37] +matrix[38][254] * vector[38] +matrix[39][254] * vector[39] +matrix[40][254] * vector[40] +matrix[41][254] * vector[41] +matrix[42][254] * vector[42] +matrix[43][254] * vector[43] +matrix[44][254] * vector[44] +matrix[45][254] * vector[45] +matrix[46][254] * vector[46] +matrix[47][254] * vector[47] +matrix[48][254] * vector[48] +matrix[49][254] * vector[49] +matrix[50][254] * vector[50] +matrix[51][254] * vector[51] +matrix[52][254] * vector[52] +matrix[53][254] * vector[53] +matrix[54][254] * vector[54] +matrix[55][254] * vector[55] +matrix[56][254] * vector[56] +matrix[57][254] * vector[57] +matrix[58][254] * vector[58] +matrix[59][254] * vector[59] +matrix[60][254] * vector[60] +matrix[61][254] * vector[61] +matrix[62][254] * vector[62] +matrix[63][254] * vector[63] +matrix[64][254] * vector[64] +matrix[65][254] * vector[65] +matrix[66][254] * vector[66] +matrix[67][254] * vector[67] +matrix[68][254] * vector[68] +matrix[69][254] * vector[69] +matrix[70][254] * vector[70] +matrix[71][254] * vector[71] +matrix[72][254] * vector[72] +matrix[73][254] * vector[73] +matrix[74][254] * vector[74] +matrix[75][254] * vector[75] +matrix[76][254] * vector[76] +matrix[77][254] * vector[77] +matrix[78][254] * vector[78] +matrix[79][254] * vector[79] +matrix[80][254] * vector[80] +matrix[81][254] * vector[81] +matrix[82][254] * vector[82] +matrix[83][254] * vector[83] +matrix[84][254] * vector[84] +matrix[85][254] * vector[85] +matrix[86][254] * vector[86] +matrix[87][254] * vector[87] +matrix[88][254] * vector[88] +matrix[89][254] * vector[89] +matrix[90][254] * vector[90] +matrix[91][254] * vector[91] +matrix[92][254] * vector[92] +matrix[93][254] * vector[93] +matrix[94][254] * vector[94] +matrix[95][254] * vector[95] +matrix[96][254] * vector[96] +matrix[97][254] * vector[97] +matrix[98][254] * vector[98] +matrix[99][254] * vector[99] +b[254];
assign result[255] = matrix[0][255] * vector[0] +matrix[1][255] * vector[1] +matrix[2][255] * vector[2] +matrix[3][255] * vector[3] +matrix[4][255] * vector[4] +matrix[5][255] * vector[5] +matrix[6][255] * vector[6] +matrix[7][255] * vector[7] +matrix[8][255] * vector[8] +matrix[9][255] * vector[9] +matrix[10][255] * vector[10] +matrix[11][255] * vector[11] +matrix[12][255] * vector[12] +matrix[13][255] * vector[13] +matrix[14][255] * vector[14] +matrix[15][255] * vector[15] +matrix[16][255] * vector[16] +matrix[17][255] * vector[17] +matrix[18][255] * vector[18] +matrix[19][255] * vector[19] +matrix[20][255] * vector[20] +matrix[21][255] * vector[21] +matrix[22][255] * vector[22] +matrix[23][255] * vector[23] +matrix[24][255] * vector[24] +matrix[25][255] * vector[25] +matrix[26][255] * vector[26] +matrix[27][255] * vector[27] +matrix[28][255] * vector[28] +matrix[29][255] * vector[29] +matrix[30][255] * vector[30] +matrix[31][255] * vector[31] +matrix[32][255] * vector[32] +matrix[33][255] * vector[33] +matrix[34][255] * vector[34] +matrix[35][255] * vector[35] +matrix[36][255] * vector[36] +matrix[37][255] * vector[37] +matrix[38][255] * vector[38] +matrix[39][255] * vector[39] +matrix[40][255] * vector[40] +matrix[41][255] * vector[41] +matrix[42][255] * vector[42] +matrix[43][255] * vector[43] +matrix[44][255] * vector[44] +matrix[45][255] * vector[45] +matrix[46][255] * vector[46] +matrix[47][255] * vector[47] +matrix[48][255] * vector[48] +matrix[49][255] * vector[49] +matrix[50][255] * vector[50] +matrix[51][255] * vector[51] +matrix[52][255] * vector[52] +matrix[53][255] * vector[53] +matrix[54][255] * vector[54] +matrix[55][255] * vector[55] +matrix[56][255] * vector[56] +matrix[57][255] * vector[57] +matrix[58][255] * vector[58] +matrix[59][255] * vector[59] +matrix[60][255] * vector[60] +matrix[61][255] * vector[61] +matrix[62][255] * vector[62] +matrix[63][255] * vector[63] +matrix[64][255] * vector[64] +matrix[65][255] * vector[65] +matrix[66][255] * vector[66] +matrix[67][255] * vector[67] +matrix[68][255] * vector[68] +matrix[69][255] * vector[69] +matrix[70][255] * vector[70] +matrix[71][255] * vector[71] +matrix[72][255] * vector[72] +matrix[73][255] * vector[73] +matrix[74][255] * vector[74] +matrix[75][255] * vector[75] +matrix[76][255] * vector[76] +matrix[77][255] * vector[77] +matrix[78][255] * vector[78] +matrix[79][255] * vector[79] +matrix[80][255] * vector[80] +matrix[81][255] * vector[81] +matrix[82][255] * vector[82] +matrix[83][255] * vector[83] +matrix[84][255] * vector[84] +matrix[85][255] * vector[85] +matrix[86][255] * vector[86] +matrix[87][255] * vector[87] +matrix[88][255] * vector[88] +matrix[89][255] * vector[89] +matrix[90][255] * vector[90] +matrix[91][255] * vector[91] +matrix[92][255] * vector[92] +matrix[93][255] * vector[93] +matrix[94][255] * vector[94] +matrix[95][255] * vector[95] +matrix[96][255] * vector[96] +matrix[97][255] * vector[97] +matrix[98][255] * vector[98] +matrix[99][255] * vector[99] +b[255];
assign result[256] = matrix[0][256] * vector[0] +matrix[1][256] * vector[1] +matrix[2][256] * vector[2] +matrix[3][256] * vector[3] +matrix[4][256] * vector[4] +matrix[5][256] * vector[5] +matrix[6][256] * vector[6] +matrix[7][256] * vector[7] +matrix[8][256] * vector[8] +matrix[9][256] * vector[9] +matrix[10][256] * vector[10] +matrix[11][256] * vector[11] +matrix[12][256] * vector[12] +matrix[13][256] * vector[13] +matrix[14][256] * vector[14] +matrix[15][256] * vector[15] +matrix[16][256] * vector[16] +matrix[17][256] * vector[17] +matrix[18][256] * vector[18] +matrix[19][256] * vector[19] +matrix[20][256] * vector[20] +matrix[21][256] * vector[21] +matrix[22][256] * vector[22] +matrix[23][256] * vector[23] +matrix[24][256] * vector[24] +matrix[25][256] * vector[25] +matrix[26][256] * vector[26] +matrix[27][256] * vector[27] +matrix[28][256] * vector[28] +matrix[29][256] * vector[29] +matrix[30][256] * vector[30] +matrix[31][256] * vector[31] +matrix[32][256] * vector[32] +matrix[33][256] * vector[33] +matrix[34][256] * vector[34] +matrix[35][256] * vector[35] +matrix[36][256] * vector[36] +matrix[37][256] * vector[37] +matrix[38][256] * vector[38] +matrix[39][256] * vector[39] +matrix[40][256] * vector[40] +matrix[41][256] * vector[41] +matrix[42][256] * vector[42] +matrix[43][256] * vector[43] +matrix[44][256] * vector[44] +matrix[45][256] * vector[45] +matrix[46][256] * vector[46] +matrix[47][256] * vector[47] +matrix[48][256] * vector[48] +matrix[49][256] * vector[49] +matrix[50][256] * vector[50] +matrix[51][256] * vector[51] +matrix[52][256] * vector[52] +matrix[53][256] * vector[53] +matrix[54][256] * vector[54] +matrix[55][256] * vector[55] +matrix[56][256] * vector[56] +matrix[57][256] * vector[57] +matrix[58][256] * vector[58] +matrix[59][256] * vector[59] +matrix[60][256] * vector[60] +matrix[61][256] * vector[61] +matrix[62][256] * vector[62] +matrix[63][256] * vector[63] +matrix[64][256] * vector[64] +matrix[65][256] * vector[65] +matrix[66][256] * vector[66] +matrix[67][256] * vector[67] +matrix[68][256] * vector[68] +matrix[69][256] * vector[69] +matrix[70][256] * vector[70] +matrix[71][256] * vector[71] +matrix[72][256] * vector[72] +matrix[73][256] * vector[73] +matrix[74][256] * vector[74] +matrix[75][256] * vector[75] +matrix[76][256] * vector[76] +matrix[77][256] * vector[77] +matrix[78][256] * vector[78] +matrix[79][256] * vector[79] +matrix[80][256] * vector[80] +matrix[81][256] * vector[81] +matrix[82][256] * vector[82] +matrix[83][256] * vector[83] +matrix[84][256] * vector[84] +matrix[85][256] * vector[85] +matrix[86][256] * vector[86] +matrix[87][256] * vector[87] +matrix[88][256] * vector[88] +matrix[89][256] * vector[89] +matrix[90][256] * vector[90] +matrix[91][256] * vector[91] +matrix[92][256] * vector[92] +matrix[93][256] * vector[93] +matrix[94][256] * vector[94] +matrix[95][256] * vector[95] +matrix[96][256] * vector[96] +matrix[97][256] * vector[97] +matrix[98][256] * vector[98] +matrix[99][256] * vector[99] +b[256];
assign result[257] = matrix[0][257] * vector[0] +matrix[1][257] * vector[1] +matrix[2][257] * vector[2] +matrix[3][257] * vector[3] +matrix[4][257] * vector[4] +matrix[5][257] * vector[5] +matrix[6][257] * vector[6] +matrix[7][257] * vector[7] +matrix[8][257] * vector[8] +matrix[9][257] * vector[9] +matrix[10][257] * vector[10] +matrix[11][257] * vector[11] +matrix[12][257] * vector[12] +matrix[13][257] * vector[13] +matrix[14][257] * vector[14] +matrix[15][257] * vector[15] +matrix[16][257] * vector[16] +matrix[17][257] * vector[17] +matrix[18][257] * vector[18] +matrix[19][257] * vector[19] +matrix[20][257] * vector[20] +matrix[21][257] * vector[21] +matrix[22][257] * vector[22] +matrix[23][257] * vector[23] +matrix[24][257] * vector[24] +matrix[25][257] * vector[25] +matrix[26][257] * vector[26] +matrix[27][257] * vector[27] +matrix[28][257] * vector[28] +matrix[29][257] * vector[29] +matrix[30][257] * vector[30] +matrix[31][257] * vector[31] +matrix[32][257] * vector[32] +matrix[33][257] * vector[33] +matrix[34][257] * vector[34] +matrix[35][257] * vector[35] +matrix[36][257] * vector[36] +matrix[37][257] * vector[37] +matrix[38][257] * vector[38] +matrix[39][257] * vector[39] +matrix[40][257] * vector[40] +matrix[41][257] * vector[41] +matrix[42][257] * vector[42] +matrix[43][257] * vector[43] +matrix[44][257] * vector[44] +matrix[45][257] * vector[45] +matrix[46][257] * vector[46] +matrix[47][257] * vector[47] +matrix[48][257] * vector[48] +matrix[49][257] * vector[49] +matrix[50][257] * vector[50] +matrix[51][257] * vector[51] +matrix[52][257] * vector[52] +matrix[53][257] * vector[53] +matrix[54][257] * vector[54] +matrix[55][257] * vector[55] +matrix[56][257] * vector[56] +matrix[57][257] * vector[57] +matrix[58][257] * vector[58] +matrix[59][257] * vector[59] +matrix[60][257] * vector[60] +matrix[61][257] * vector[61] +matrix[62][257] * vector[62] +matrix[63][257] * vector[63] +matrix[64][257] * vector[64] +matrix[65][257] * vector[65] +matrix[66][257] * vector[66] +matrix[67][257] * vector[67] +matrix[68][257] * vector[68] +matrix[69][257] * vector[69] +matrix[70][257] * vector[70] +matrix[71][257] * vector[71] +matrix[72][257] * vector[72] +matrix[73][257] * vector[73] +matrix[74][257] * vector[74] +matrix[75][257] * vector[75] +matrix[76][257] * vector[76] +matrix[77][257] * vector[77] +matrix[78][257] * vector[78] +matrix[79][257] * vector[79] +matrix[80][257] * vector[80] +matrix[81][257] * vector[81] +matrix[82][257] * vector[82] +matrix[83][257] * vector[83] +matrix[84][257] * vector[84] +matrix[85][257] * vector[85] +matrix[86][257] * vector[86] +matrix[87][257] * vector[87] +matrix[88][257] * vector[88] +matrix[89][257] * vector[89] +matrix[90][257] * vector[90] +matrix[91][257] * vector[91] +matrix[92][257] * vector[92] +matrix[93][257] * vector[93] +matrix[94][257] * vector[94] +matrix[95][257] * vector[95] +matrix[96][257] * vector[96] +matrix[97][257] * vector[97] +matrix[98][257] * vector[98] +matrix[99][257] * vector[99] +b[257];
assign result[258] = matrix[0][258] * vector[0] +matrix[1][258] * vector[1] +matrix[2][258] * vector[2] +matrix[3][258] * vector[3] +matrix[4][258] * vector[4] +matrix[5][258] * vector[5] +matrix[6][258] * vector[6] +matrix[7][258] * vector[7] +matrix[8][258] * vector[8] +matrix[9][258] * vector[9] +matrix[10][258] * vector[10] +matrix[11][258] * vector[11] +matrix[12][258] * vector[12] +matrix[13][258] * vector[13] +matrix[14][258] * vector[14] +matrix[15][258] * vector[15] +matrix[16][258] * vector[16] +matrix[17][258] * vector[17] +matrix[18][258] * vector[18] +matrix[19][258] * vector[19] +matrix[20][258] * vector[20] +matrix[21][258] * vector[21] +matrix[22][258] * vector[22] +matrix[23][258] * vector[23] +matrix[24][258] * vector[24] +matrix[25][258] * vector[25] +matrix[26][258] * vector[26] +matrix[27][258] * vector[27] +matrix[28][258] * vector[28] +matrix[29][258] * vector[29] +matrix[30][258] * vector[30] +matrix[31][258] * vector[31] +matrix[32][258] * vector[32] +matrix[33][258] * vector[33] +matrix[34][258] * vector[34] +matrix[35][258] * vector[35] +matrix[36][258] * vector[36] +matrix[37][258] * vector[37] +matrix[38][258] * vector[38] +matrix[39][258] * vector[39] +matrix[40][258] * vector[40] +matrix[41][258] * vector[41] +matrix[42][258] * vector[42] +matrix[43][258] * vector[43] +matrix[44][258] * vector[44] +matrix[45][258] * vector[45] +matrix[46][258] * vector[46] +matrix[47][258] * vector[47] +matrix[48][258] * vector[48] +matrix[49][258] * vector[49] +matrix[50][258] * vector[50] +matrix[51][258] * vector[51] +matrix[52][258] * vector[52] +matrix[53][258] * vector[53] +matrix[54][258] * vector[54] +matrix[55][258] * vector[55] +matrix[56][258] * vector[56] +matrix[57][258] * vector[57] +matrix[58][258] * vector[58] +matrix[59][258] * vector[59] +matrix[60][258] * vector[60] +matrix[61][258] * vector[61] +matrix[62][258] * vector[62] +matrix[63][258] * vector[63] +matrix[64][258] * vector[64] +matrix[65][258] * vector[65] +matrix[66][258] * vector[66] +matrix[67][258] * vector[67] +matrix[68][258] * vector[68] +matrix[69][258] * vector[69] +matrix[70][258] * vector[70] +matrix[71][258] * vector[71] +matrix[72][258] * vector[72] +matrix[73][258] * vector[73] +matrix[74][258] * vector[74] +matrix[75][258] * vector[75] +matrix[76][258] * vector[76] +matrix[77][258] * vector[77] +matrix[78][258] * vector[78] +matrix[79][258] * vector[79] +matrix[80][258] * vector[80] +matrix[81][258] * vector[81] +matrix[82][258] * vector[82] +matrix[83][258] * vector[83] +matrix[84][258] * vector[84] +matrix[85][258] * vector[85] +matrix[86][258] * vector[86] +matrix[87][258] * vector[87] +matrix[88][258] * vector[88] +matrix[89][258] * vector[89] +matrix[90][258] * vector[90] +matrix[91][258] * vector[91] +matrix[92][258] * vector[92] +matrix[93][258] * vector[93] +matrix[94][258] * vector[94] +matrix[95][258] * vector[95] +matrix[96][258] * vector[96] +matrix[97][258] * vector[97] +matrix[98][258] * vector[98] +matrix[99][258] * vector[99] +b[258];
assign result[259] = matrix[0][259] * vector[0] +matrix[1][259] * vector[1] +matrix[2][259] * vector[2] +matrix[3][259] * vector[3] +matrix[4][259] * vector[4] +matrix[5][259] * vector[5] +matrix[6][259] * vector[6] +matrix[7][259] * vector[7] +matrix[8][259] * vector[8] +matrix[9][259] * vector[9] +matrix[10][259] * vector[10] +matrix[11][259] * vector[11] +matrix[12][259] * vector[12] +matrix[13][259] * vector[13] +matrix[14][259] * vector[14] +matrix[15][259] * vector[15] +matrix[16][259] * vector[16] +matrix[17][259] * vector[17] +matrix[18][259] * vector[18] +matrix[19][259] * vector[19] +matrix[20][259] * vector[20] +matrix[21][259] * vector[21] +matrix[22][259] * vector[22] +matrix[23][259] * vector[23] +matrix[24][259] * vector[24] +matrix[25][259] * vector[25] +matrix[26][259] * vector[26] +matrix[27][259] * vector[27] +matrix[28][259] * vector[28] +matrix[29][259] * vector[29] +matrix[30][259] * vector[30] +matrix[31][259] * vector[31] +matrix[32][259] * vector[32] +matrix[33][259] * vector[33] +matrix[34][259] * vector[34] +matrix[35][259] * vector[35] +matrix[36][259] * vector[36] +matrix[37][259] * vector[37] +matrix[38][259] * vector[38] +matrix[39][259] * vector[39] +matrix[40][259] * vector[40] +matrix[41][259] * vector[41] +matrix[42][259] * vector[42] +matrix[43][259] * vector[43] +matrix[44][259] * vector[44] +matrix[45][259] * vector[45] +matrix[46][259] * vector[46] +matrix[47][259] * vector[47] +matrix[48][259] * vector[48] +matrix[49][259] * vector[49] +matrix[50][259] * vector[50] +matrix[51][259] * vector[51] +matrix[52][259] * vector[52] +matrix[53][259] * vector[53] +matrix[54][259] * vector[54] +matrix[55][259] * vector[55] +matrix[56][259] * vector[56] +matrix[57][259] * vector[57] +matrix[58][259] * vector[58] +matrix[59][259] * vector[59] +matrix[60][259] * vector[60] +matrix[61][259] * vector[61] +matrix[62][259] * vector[62] +matrix[63][259] * vector[63] +matrix[64][259] * vector[64] +matrix[65][259] * vector[65] +matrix[66][259] * vector[66] +matrix[67][259] * vector[67] +matrix[68][259] * vector[68] +matrix[69][259] * vector[69] +matrix[70][259] * vector[70] +matrix[71][259] * vector[71] +matrix[72][259] * vector[72] +matrix[73][259] * vector[73] +matrix[74][259] * vector[74] +matrix[75][259] * vector[75] +matrix[76][259] * vector[76] +matrix[77][259] * vector[77] +matrix[78][259] * vector[78] +matrix[79][259] * vector[79] +matrix[80][259] * vector[80] +matrix[81][259] * vector[81] +matrix[82][259] * vector[82] +matrix[83][259] * vector[83] +matrix[84][259] * vector[84] +matrix[85][259] * vector[85] +matrix[86][259] * vector[86] +matrix[87][259] * vector[87] +matrix[88][259] * vector[88] +matrix[89][259] * vector[89] +matrix[90][259] * vector[90] +matrix[91][259] * vector[91] +matrix[92][259] * vector[92] +matrix[93][259] * vector[93] +matrix[94][259] * vector[94] +matrix[95][259] * vector[95] +matrix[96][259] * vector[96] +matrix[97][259] * vector[97] +matrix[98][259] * vector[98] +matrix[99][259] * vector[99] +b[259];
assign result[260] = matrix[0][260] * vector[0] +matrix[1][260] * vector[1] +matrix[2][260] * vector[2] +matrix[3][260] * vector[3] +matrix[4][260] * vector[4] +matrix[5][260] * vector[5] +matrix[6][260] * vector[6] +matrix[7][260] * vector[7] +matrix[8][260] * vector[8] +matrix[9][260] * vector[9] +matrix[10][260] * vector[10] +matrix[11][260] * vector[11] +matrix[12][260] * vector[12] +matrix[13][260] * vector[13] +matrix[14][260] * vector[14] +matrix[15][260] * vector[15] +matrix[16][260] * vector[16] +matrix[17][260] * vector[17] +matrix[18][260] * vector[18] +matrix[19][260] * vector[19] +matrix[20][260] * vector[20] +matrix[21][260] * vector[21] +matrix[22][260] * vector[22] +matrix[23][260] * vector[23] +matrix[24][260] * vector[24] +matrix[25][260] * vector[25] +matrix[26][260] * vector[26] +matrix[27][260] * vector[27] +matrix[28][260] * vector[28] +matrix[29][260] * vector[29] +matrix[30][260] * vector[30] +matrix[31][260] * vector[31] +matrix[32][260] * vector[32] +matrix[33][260] * vector[33] +matrix[34][260] * vector[34] +matrix[35][260] * vector[35] +matrix[36][260] * vector[36] +matrix[37][260] * vector[37] +matrix[38][260] * vector[38] +matrix[39][260] * vector[39] +matrix[40][260] * vector[40] +matrix[41][260] * vector[41] +matrix[42][260] * vector[42] +matrix[43][260] * vector[43] +matrix[44][260] * vector[44] +matrix[45][260] * vector[45] +matrix[46][260] * vector[46] +matrix[47][260] * vector[47] +matrix[48][260] * vector[48] +matrix[49][260] * vector[49] +matrix[50][260] * vector[50] +matrix[51][260] * vector[51] +matrix[52][260] * vector[52] +matrix[53][260] * vector[53] +matrix[54][260] * vector[54] +matrix[55][260] * vector[55] +matrix[56][260] * vector[56] +matrix[57][260] * vector[57] +matrix[58][260] * vector[58] +matrix[59][260] * vector[59] +matrix[60][260] * vector[60] +matrix[61][260] * vector[61] +matrix[62][260] * vector[62] +matrix[63][260] * vector[63] +matrix[64][260] * vector[64] +matrix[65][260] * vector[65] +matrix[66][260] * vector[66] +matrix[67][260] * vector[67] +matrix[68][260] * vector[68] +matrix[69][260] * vector[69] +matrix[70][260] * vector[70] +matrix[71][260] * vector[71] +matrix[72][260] * vector[72] +matrix[73][260] * vector[73] +matrix[74][260] * vector[74] +matrix[75][260] * vector[75] +matrix[76][260] * vector[76] +matrix[77][260] * vector[77] +matrix[78][260] * vector[78] +matrix[79][260] * vector[79] +matrix[80][260] * vector[80] +matrix[81][260] * vector[81] +matrix[82][260] * vector[82] +matrix[83][260] * vector[83] +matrix[84][260] * vector[84] +matrix[85][260] * vector[85] +matrix[86][260] * vector[86] +matrix[87][260] * vector[87] +matrix[88][260] * vector[88] +matrix[89][260] * vector[89] +matrix[90][260] * vector[90] +matrix[91][260] * vector[91] +matrix[92][260] * vector[92] +matrix[93][260] * vector[93] +matrix[94][260] * vector[94] +matrix[95][260] * vector[95] +matrix[96][260] * vector[96] +matrix[97][260] * vector[97] +matrix[98][260] * vector[98] +matrix[99][260] * vector[99] +b[260];
assign result[261] = matrix[0][261] * vector[0] +matrix[1][261] * vector[1] +matrix[2][261] * vector[2] +matrix[3][261] * vector[3] +matrix[4][261] * vector[4] +matrix[5][261] * vector[5] +matrix[6][261] * vector[6] +matrix[7][261] * vector[7] +matrix[8][261] * vector[8] +matrix[9][261] * vector[9] +matrix[10][261] * vector[10] +matrix[11][261] * vector[11] +matrix[12][261] * vector[12] +matrix[13][261] * vector[13] +matrix[14][261] * vector[14] +matrix[15][261] * vector[15] +matrix[16][261] * vector[16] +matrix[17][261] * vector[17] +matrix[18][261] * vector[18] +matrix[19][261] * vector[19] +matrix[20][261] * vector[20] +matrix[21][261] * vector[21] +matrix[22][261] * vector[22] +matrix[23][261] * vector[23] +matrix[24][261] * vector[24] +matrix[25][261] * vector[25] +matrix[26][261] * vector[26] +matrix[27][261] * vector[27] +matrix[28][261] * vector[28] +matrix[29][261] * vector[29] +matrix[30][261] * vector[30] +matrix[31][261] * vector[31] +matrix[32][261] * vector[32] +matrix[33][261] * vector[33] +matrix[34][261] * vector[34] +matrix[35][261] * vector[35] +matrix[36][261] * vector[36] +matrix[37][261] * vector[37] +matrix[38][261] * vector[38] +matrix[39][261] * vector[39] +matrix[40][261] * vector[40] +matrix[41][261] * vector[41] +matrix[42][261] * vector[42] +matrix[43][261] * vector[43] +matrix[44][261] * vector[44] +matrix[45][261] * vector[45] +matrix[46][261] * vector[46] +matrix[47][261] * vector[47] +matrix[48][261] * vector[48] +matrix[49][261] * vector[49] +matrix[50][261] * vector[50] +matrix[51][261] * vector[51] +matrix[52][261] * vector[52] +matrix[53][261] * vector[53] +matrix[54][261] * vector[54] +matrix[55][261] * vector[55] +matrix[56][261] * vector[56] +matrix[57][261] * vector[57] +matrix[58][261] * vector[58] +matrix[59][261] * vector[59] +matrix[60][261] * vector[60] +matrix[61][261] * vector[61] +matrix[62][261] * vector[62] +matrix[63][261] * vector[63] +matrix[64][261] * vector[64] +matrix[65][261] * vector[65] +matrix[66][261] * vector[66] +matrix[67][261] * vector[67] +matrix[68][261] * vector[68] +matrix[69][261] * vector[69] +matrix[70][261] * vector[70] +matrix[71][261] * vector[71] +matrix[72][261] * vector[72] +matrix[73][261] * vector[73] +matrix[74][261] * vector[74] +matrix[75][261] * vector[75] +matrix[76][261] * vector[76] +matrix[77][261] * vector[77] +matrix[78][261] * vector[78] +matrix[79][261] * vector[79] +matrix[80][261] * vector[80] +matrix[81][261] * vector[81] +matrix[82][261] * vector[82] +matrix[83][261] * vector[83] +matrix[84][261] * vector[84] +matrix[85][261] * vector[85] +matrix[86][261] * vector[86] +matrix[87][261] * vector[87] +matrix[88][261] * vector[88] +matrix[89][261] * vector[89] +matrix[90][261] * vector[90] +matrix[91][261] * vector[91] +matrix[92][261] * vector[92] +matrix[93][261] * vector[93] +matrix[94][261] * vector[94] +matrix[95][261] * vector[95] +matrix[96][261] * vector[96] +matrix[97][261] * vector[97] +matrix[98][261] * vector[98] +matrix[99][261] * vector[99] +b[261];
assign result[262] = matrix[0][262] * vector[0] +matrix[1][262] * vector[1] +matrix[2][262] * vector[2] +matrix[3][262] * vector[3] +matrix[4][262] * vector[4] +matrix[5][262] * vector[5] +matrix[6][262] * vector[6] +matrix[7][262] * vector[7] +matrix[8][262] * vector[8] +matrix[9][262] * vector[9] +matrix[10][262] * vector[10] +matrix[11][262] * vector[11] +matrix[12][262] * vector[12] +matrix[13][262] * vector[13] +matrix[14][262] * vector[14] +matrix[15][262] * vector[15] +matrix[16][262] * vector[16] +matrix[17][262] * vector[17] +matrix[18][262] * vector[18] +matrix[19][262] * vector[19] +matrix[20][262] * vector[20] +matrix[21][262] * vector[21] +matrix[22][262] * vector[22] +matrix[23][262] * vector[23] +matrix[24][262] * vector[24] +matrix[25][262] * vector[25] +matrix[26][262] * vector[26] +matrix[27][262] * vector[27] +matrix[28][262] * vector[28] +matrix[29][262] * vector[29] +matrix[30][262] * vector[30] +matrix[31][262] * vector[31] +matrix[32][262] * vector[32] +matrix[33][262] * vector[33] +matrix[34][262] * vector[34] +matrix[35][262] * vector[35] +matrix[36][262] * vector[36] +matrix[37][262] * vector[37] +matrix[38][262] * vector[38] +matrix[39][262] * vector[39] +matrix[40][262] * vector[40] +matrix[41][262] * vector[41] +matrix[42][262] * vector[42] +matrix[43][262] * vector[43] +matrix[44][262] * vector[44] +matrix[45][262] * vector[45] +matrix[46][262] * vector[46] +matrix[47][262] * vector[47] +matrix[48][262] * vector[48] +matrix[49][262] * vector[49] +matrix[50][262] * vector[50] +matrix[51][262] * vector[51] +matrix[52][262] * vector[52] +matrix[53][262] * vector[53] +matrix[54][262] * vector[54] +matrix[55][262] * vector[55] +matrix[56][262] * vector[56] +matrix[57][262] * vector[57] +matrix[58][262] * vector[58] +matrix[59][262] * vector[59] +matrix[60][262] * vector[60] +matrix[61][262] * vector[61] +matrix[62][262] * vector[62] +matrix[63][262] * vector[63] +matrix[64][262] * vector[64] +matrix[65][262] * vector[65] +matrix[66][262] * vector[66] +matrix[67][262] * vector[67] +matrix[68][262] * vector[68] +matrix[69][262] * vector[69] +matrix[70][262] * vector[70] +matrix[71][262] * vector[71] +matrix[72][262] * vector[72] +matrix[73][262] * vector[73] +matrix[74][262] * vector[74] +matrix[75][262] * vector[75] +matrix[76][262] * vector[76] +matrix[77][262] * vector[77] +matrix[78][262] * vector[78] +matrix[79][262] * vector[79] +matrix[80][262] * vector[80] +matrix[81][262] * vector[81] +matrix[82][262] * vector[82] +matrix[83][262] * vector[83] +matrix[84][262] * vector[84] +matrix[85][262] * vector[85] +matrix[86][262] * vector[86] +matrix[87][262] * vector[87] +matrix[88][262] * vector[88] +matrix[89][262] * vector[89] +matrix[90][262] * vector[90] +matrix[91][262] * vector[91] +matrix[92][262] * vector[92] +matrix[93][262] * vector[93] +matrix[94][262] * vector[94] +matrix[95][262] * vector[95] +matrix[96][262] * vector[96] +matrix[97][262] * vector[97] +matrix[98][262] * vector[98] +matrix[99][262] * vector[99] +b[262];
assign result[263] = matrix[0][263] * vector[0] +matrix[1][263] * vector[1] +matrix[2][263] * vector[2] +matrix[3][263] * vector[3] +matrix[4][263] * vector[4] +matrix[5][263] * vector[5] +matrix[6][263] * vector[6] +matrix[7][263] * vector[7] +matrix[8][263] * vector[8] +matrix[9][263] * vector[9] +matrix[10][263] * vector[10] +matrix[11][263] * vector[11] +matrix[12][263] * vector[12] +matrix[13][263] * vector[13] +matrix[14][263] * vector[14] +matrix[15][263] * vector[15] +matrix[16][263] * vector[16] +matrix[17][263] * vector[17] +matrix[18][263] * vector[18] +matrix[19][263] * vector[19] +matrix[20][263] * vector[20] +matrix[21][263] * vector[21] +matrix[22][263] * vector[22] +matrix[23][263] * vector[23] +matrix[24][263] * vector[24] +matrix[25][263] * vector[25] +matrix[26][263] * vector[26] +matrix[27][263] * vector[27] +matrix[28][263] * vector[28] +matrix[29][263] * vector[29] +matrix[30][263] * vector[30] +matrix[31][263] * vector[31] +matrix[32][263] * vector[32] +matrix[33][263] * vector[33] +matrix[34][263] * vector[34] +matrix[35][263] * vector[35] +matrix[36][263] * vector[36] +matrix[37][263] * vector[37] +matrix[38][263] * vector[38] +matrix[39][263] * vector[39] +matrix[40][263] * vector[40] +matrix[41][263] * vector[41] +matrix[42][263] * vector[42] +matrix[43][263] * vector[43] +matrix[44][263] * vector[44] +matrix[45][263] * vector[45] +matrix[46][263] * vector[46] +matrix[47][263] * vector[47] +matrix[48][263] * vector[48] +matrix[49][263] * vector[49] +matrix[50][263] * vector[50] +matrix[51][263] * vector[51] +matrix[52][263] * vector[52] +matrix[53][263] * vector[53] +matrix[54][263] * vector[54] +matrix[55][263] * vector[55] +matrix[56][263] * vector[56] +matrix[57][263] * vector[57] +matrix[58][263] * vector[58] +matrix[59][263] * vector[59] +matrix[60][263] * vector[60] +matrix[61][263] * vector[61] +matrix[62][263] * vector[62] +matrix[63][263] * vector[63] +matrix[64][263] * vector[64] +matrix[65][263] * vector[65] +matrix[66][263] * vector[66] +matrix[67][263] * vector[67] +matrix[68][263] * vector[68] +matrix[69][263] * vector[69] +matrix[70][263] * vector[70] +matrix[71][263] * vector[71] +matrix[72][263] * vector[72] +matrix[73][263] * vector[73] +matrix[74][263] * vector[74] +matrix[75][263] * vector[75] +matrix[76][263] * vector[76] +matrix[77][263] * vector[77] +matrix[78][263] * vector[78] +matrix[79][263] * vector[79] +matrix[80][263] * vector[80] +matrix[81][263] * vector[81] +matrix[82][263] * vector[82] +matrix[83][263] * vector[83] +matrix[84][263] * vector[84] +matrix[85][263] * vector[85] +matrix[86][263] * vector[86] +matrix[87][263] * vector[87] +matrix[88][263] * vector[88] +matrix[89][263] * vector[89] +matrix[90][263] * vector[90] +matrix[91][263] * vector[91] +matrix[92][263] * vector[92] +matrix[93][263] * vector[93] +matrix[94][263] * vector[94] +matrix[95][263] * vector[95] +matrix[96][263] * vector[96] +matrix[97][263] * vector[97] +matrix[98][263] * vector[98] +matrix[99][263] * vector[99] +b[263];
assign result[264] = matrix[0][264] * vector[0] +matrix[1][264] * vector[1] +matrix[2][264] * vector[2] +matrix[3][264] * vector[3] +matrix[4][264] * vector[4] +matrix[5][264] * vector[5] +matrix[6][264] * vector[6] +matrix[7][264] * vector[7] +matrix[8][264] * vector[8] +matrix[9][264] * vector[9] +matrix[10][264] * vector[10] +matrix[11][264] * vector[11] +matrix[12][264] * vector[12] +matrix[13][264] * vector[13] +matrix[14][264] * vector[14] +matrix[15][264] * vector[15] +matrix[16][264] * vector[16] +matrix[17][264] * vector[17] +matrix[18][264] * vector[18] +matrix[19][264] * vector[19] +matrix[20][264] * vector[20] +matrix[21][264] * vector[21] +matrix[22][264] * vector[22] +matrix[23][264] * vector[23] +matrix[24][264] * vector[24] +matrix[25][264] * vector[25] +matrix[26][264] * vector[26] +matrix[27][264] * vector[27] +matrix[28][264] * vector[28] +matrix[29][264] * vector[29] +matrix[30][264] * vector[30] +matrix[31][264] * vector[31] +matrix[32][264] * vector[32] +matrix[33][264] * vector[33] +matrix[34][264] * vector[34] +matrix[35][264] * vector[35] +matrix[36][264] * vector[36] +matrix[37][264] * vector[37] +matrix[38][264] * vector[38] +matrix[39][264] * vector[39] +matrix[40][264] * vector[40] +matrix[41][264] * vector[41] +matrix[42][264] * vector[42] +matrix[43][264] * vector[43] +matrix[44][264] * vector[44] +matrix[45][264] * vector[45] +matrix[46][264] * vector[46] +matrix[47][264] * vector[47] +matrix[48][264] * vector[48] +matrix[49][264] * vector[49] +matrix[50][264] * vector[50] +matrix[51][264] * vector[51] +matrix[52][264] * vector[52] +matrix[53][264] * vector[53] +matrix[54][264] * vector[54] +matrix[55][264] * vector[55] +matrix[56][264] * vector[56] +matrix[57][264] * vector[57] +matrix[58][264] * vector[58] +matrix[59][264] * vector[59] +matrix[60][264] * vector[60] +matrix[61][264] * vector[61] +matrix[62][264] * vector[62] +matrix[63][264] * vector[63] +matrix[64][264] * vector[64] +matrix[65][264] * vector[65] +matrix[66][264] * vector[66] +matrix[67][264] * vector[67] +matrix[68][264] * vector[68] +matrix[69][264] * vector[69] +matrix[70][264] * vector[70] +matrix[71][264] * vector[71] +matrix[72][264] * vector[72] +matrix[73][264] * vector[73] +matrix[74][264] * vector[74] +matrix[75][264] * vector[75] +matrix[76][264] * vector[76] +matrix[77][264] * vector[77] +matrix[78][264] * vector[78] +matrix[79][264] * vector[79] +matrix[80][264] * vector[80] +matrix[81][264] * vector[81] +matrix[82][264] * vector[82] +matrix[83][264] * vector[83] +matrix[84][264] * vector[84] +matrix[85][264] * vector[85] +matrix[86][264] * vector[86] +matrix[87][264] * vector[87] +matrix[88][264] * vector[88] +matrix[89][264] * vector[89] +matrix[90][264] * vector[90] +matrix[91][264] * vector[91] +matrix[92][264] * vector[92] +matrix[93][264] * vector[93] +matrix[94][264] * vector[94] +matrix[95][264] * vector[95] +matrix[96][264] * vector[96] +matrix[97][264] * vector[97] +matrix[98][264] * vector[98] +matrix[99][264] * vector[99] +b[264];
assign result[265] = matrix[0][265] * vector[0] +matrix[1][265] * vector[1] +matrix[2][265] * vector[2] +matrix[3][265] * vector[3] +matrix[4][265] * vector[4] +matrix[5][265] * vector[5] +matrix[6][265] * vector[6] +matrix[7][265] * vector[7] +matrix[8][265] * vector[8] +matrix[9][265] * vector[9] +matrix[10][265] * vector[10] +matrix[11][265] * vector[11] +matrix[12][265] * vector[12] +matrix[13][265] * vector[13] +matrix[14][265] * vector[14] +matrix[15][265] * vector[15] +matrix[16][265] * vector[16] +matrix[17][265] * vector[17] +matrix[18][265] * vector[18] +matrix[19][265] * vector[19] +matrix[20][265] * vector[20] +matrix[21][265] * vector[21] +matrix[22][265] * vector[22] +matrix[23][265] * vector[23] +matrix[24][265] * vector[24] +matrix[25][265] * vector[25] +matrix[26][265] * vector[26] +matrix[27][265] * vector[27] +matrix[28][265] * vector[28] +matrix[29][265] * vector[29] +matrix[30][265] * vector[30] +matrix[31][265] * vector[31] +matrix[32][265] * vector[32] +matrix[33][265] * vector[33] +matrix[34][265] * vector[34] +matrix[35][265] * vector[35] +matrix[36][265] * vector[36] +matrix[37][265] * vector[37] +matrix[38][265] * vector[38] +matrix[39][265] * vector[39] +matrix[40][265] * vector[40] +matrix[41][265] * vector[41] +matrix[42][265] * vector[42] +matrix[43][265] * vector[43] +matrix[44][265] * vector[44] +matrix[45][265] * vector[45] +matrix[46][265] * vector[46] +matrix[47][265] * vector[47] +matrix[48][265] * vector[48] +matrix[49][265] * vector[49] +matrix[50][265] * vector[50] +matrix[51][265] * vector[51] +matrix[52][265] * vector[52] +matrix[53][265] * vector[53] +matrix[54][265] * vector[54] +matrix[55][265] * vector[55] +matrix[56][265] * vector[56] +matrix[57][265] * vector[57] +matrix[58][265] * vector[58] +matrix[59][265] * vector[59] +matrix[60][265] * vector[60] +matrix[61][265] * vector[61] +matrix[62][265] * vector[62] +matrix[63][265] * vector[63] +matrix[64][265] * vector[64] +matrix[65][265] * vector[65] +matrix[66][265] * vector[66] +matrix[67][265] * vector[67] +matrix[68][265] * vector[68] +matrix[69][265] * vector[69] +matrix[70][265] * vector[70] +matrix[71][265] * vector[71] +matrix[72][265] * vector[72] +matrix[73][265] * vector[73] +matrix[74][265] * vector[74] +matrix[75][265] * vector[75] +matrix[76][265] * vector[76] +matrix[77][265] * vector[77] +matrix[78][265] * vector[78] +matrix[79][265] * vector[79] +matrix[80][265] * vector[80] +matrix[81][265] * vector[81] +matrix[82][265] * vector[82] +matrix[83][265] * vector[83] +matrix[84][265] * vector[84] +matrix[85][265] * vector[85] +matrix[86][265] * vector[86] +matrix[87][265] * vector[87] +matrix[88][265] * vector[88] +matrix[89][265] * vector[89] +matrix[90][265] * vector[90] +matrix[91][265] * vector[91] +matrix[92][265] * vector[92] +matrix[93][265] * vector[93] +matrix[94][265] * vector[94] +matrix[95][265] * vector[95] +matrix[96][265] * vector[96] +matrix[97][265] * vector[97] +matrix[98][265] * vector[98] +matrix[99][265] * vector[99] +b[265];
assign result[266] = matrix[0][266] * vector[0] +matrix[1][266] * vector[1] +matrix[2][266] * vector[2] +matrix[3][266] * vector[3] +matrix[4][266] * vector[4] +matrix[5][266] * vector[5] +matrix[6][266] * vector[6] +matrix[7][266] * vector[7] +matrix[8][266] * vector[8] +matrix[9][266] * vector[9] +matrix[10][266] * vector[10] +matrix[11][266] * vector[11] +matrix[12][266] * vector[12] +matrix[13][266] * vector[13] +matrix[14][266] * vector[14] +matrix[15][266] * vector[15] +matrix[16][266] * vector[16] +matrix[17][266] * vector[17] +matrix[18][266] * vector[18] +matrix[19][266] * vector[19] +matrix[20][266] * vector[20] +matrix[21][266] * vector[21] +matrix[22][266] * vector[22] +matrix[23][266] * vector[23] +matrix[24][266] * vector[24] +matrix[25][266] * vector[25] +matrix[26][266] * vector[26] +matrix[27][266] * vector[27] +matrix[28][266] * vector[28] +matrix[29][266] * vector[29] +matrix[30][266] * vector[30] +matrix[31][266] * vector[31] +matrix[32][266] * vector[32] +matrix[33][266] * vector[33] +matrix[34][266] * vector[34] +matrix[35][266] * vector[35] +matrix[36][266] * vector[36] +matrix[37][266] * vector[37] +matrix[38][266] * vector[38] +matrix[39][266] * vector[39] +matrix[40][266] * vector[40] +matrix[41][266] * vector[41] +matrix[42][266] * vector[42] +matrix[43][266] * vector[43] +matrix[44][266] * vector[44] +matrix[45][266] * vector[45] +matrix[46][266] * vector[46] +matrix[47][266] * vector[47] +matrix[48][266] * vector[48] +matrix[49][266] * vector[49] +matrix[50][266] * vector[50] +matrix[51][266] * vector[51] +matrix[52][266] * vector[52] +matrix[53][266] * vector[53] +matrix[54][266] * vector[54] +matrix[55][266] * vector[55] +matrix[56][266] * vector[56] +matrix[57][266] * vector[57] +matrix[58][266] * vector[58] +matrix[59][266] * vector[59] +matrix[60][266] * vector[60] +matrix[61][266] * vector[61] +matrix[62][266] * vector[62] +matrix[63][266] * vector[63] +matrix[64][266] * vector[64] +matrix[65][266] * vector[65] +matrix[66][266] * vector[66] +matrix[67][266] * vector[67] +matrix[68][266] * vector[68] +matrix[69][266] * vector[69] +matrix[70][266] * vector[70] +matrix[71][266] * vector[71] +matrix[72][266] * vector[72] +matrix[73][266] * vector[73] +matrix[74][266] * vector[74] +matrix[75][266] * vector[75] +matrix[76][266] * vector[76] +matrix[77][266] * vector[77] +matrix[78][266] * vector[78] +matrix[79][266] * vector[79] +matrix[80][266] * vector[80] +matrix[81][266] * vector[81] +matrix[82][266] * vector[82] +matrix[83][266] * vector[83] +matrix[84][266] * vector[84] +matrix[85][266] * vector[85] +matrix[86][266] * vector[86] +matrix[87][266] * vector[87] +matrix[88][266] * vector[88] +matrix[89][266] * vector[89] +matrix[90][266] * vector[90] +matrix[91][266] * vector[91] +matrix[92][266] * vector[92] +matrix[93][266] * vector[93] +matrix[94][266] * vector[94] +matrix[95][266] * vector[95] +matrix[96][266] * vector[96] +matrix[97][266] * vector[97] +matrix[98][266] * vector[98] +matrix[99][266] * vector[99] +b[266];
assign result[267] = matrix[0][267] * vector[0] +matrix[1][267] * vector[1] +matrix[2][267] * vector[2] +matrix[3][267] * vector[3] +matrix[4][267] * vector[4] +matrix[5][267] * vector[5] +matrix[6][267] * vector[6] +matrix[7][267] * vector[7] +matrix[8][267] * vector[8] +matrix[9][267] * vector[9] +matrix[10][267] * vector[10] +matrix[11][267] * vector[11] +matrix[12][267] * vector[12] +matrix[13][267] * vector[13] +matrix[14][267] * vector[14] +matrix[15][267] * vector[15] +matrix[16][267] * vector[16] +matrix[17][267] * vector[17] +matrix[18][267] * vector[18] +matrix[19][267] * vector[19] +matrix[20][267] * vector[20] +matrix[21][267] * vector[21] +matrix[22][267] * vector[22] +matrix[23][267] * vector[23] +matrix[24][267] * vector[24] +matrix[25][267] * vector[25] +matrix[26][267] * vector[26] +matrix[27][267] * vector[27] +matrix[28][267] * vector[28] +matrix[29][267] * vector[29] +matrix[30][267] * vector[30] +matrix[31][267] * vector[31] +matrix[32][267] * vector[32] +matrix[33][267] * vector[33] +matrix[34][267] * vector[34] +matrix[35][267] * vector[35] +matrix[36][267] * vector[36] +matrix[37][267] * vector[37] +matrix[38][267] * vector[38] +matrix[39][267] * vector[39] +matrix[40][267] * vector[40] +matrix[41][267] * vector[41] +matrix[42][267] * vector[42] +matrix[43][267] * vector[43] +matrix[44][267] * vector[44] +matrix[45][267] * vector[45] +matrix[46][267] * vector[46] +matrix[47][267] * vector[47] +matrix[48][267] * vector[48] +matrix[49][267] * vector[49] +matrix[50][267] * vector[50] +matrix[51][267] * vector[51] +matrix[52][267] * vector[52] +matrix[53][267] * vector[53] +matrix[54][267] * vector[54] +matrix[55][267] * vector[55] +matrix[56][267] * vector[56] +matrix[57][267] * vector[57] +matrix[58][267] * vector[58] +matrix[59][267] * vector[59] +matrix[60][267] * vector[60] +matrix[61][267] * vector[61] +matrix[62][267] * vector[62] +matrix[63][267] * vector[63] +matrix[64][267] * vector[64] +matrix[65][267] * vector[65] +matrix[66][267] * vector[66] +matrix[67][267] * vector[67] +matrix[68][267] * vector[68] +matrix[69][267] * vector[69] +matrix[70][267] * vector[70] +matrix[71][267] * vector[71] +matrix[72][267] * vector[72] +matrix[73][267] * vector[73] +matrix[74][267] * vector[74] +matrix[75][267] * vector[75] +matrix[76][267] * vector[76] +matrix[77][267] * vector[77] +matrix[78][267] * vector[78] +matrix[79][267] * vector[79] +matrix[80][267] * vector[80] +matrix[81][267] * vector[81] +matrix[82][267] * vector[82] +matrix[83][267] * vector[83] +matrix[84][267] * vector[84] +matrix[85][267] * vector[85] +matrix[86][267] * vector[86] +matrix[87][267] * vector[87] +matrix[88][267] * vector[88] +matrix[89][267] * vector[89] +matrix[90][267] * vector[90] +matrix[91][267] * vector[91] +matrix[92][267] * vector[92] +matrix[93][267] * vector[93] +matrix[94][267] * vector[94] +matrix[95][267] * vector[95] +matrix[96][267] * vector[96] +matrix[97][267] * vector[97] +matrix[98][267] * vector[98] +matrix[99][267] * vector[99] +b[267];
assign result[268] = matrix[0][268] * vector[0] +matrix[1][268] * vector[1] +matrix[2][268] * vector[2] +matrix[3][268] * vector[3] +matrix[4][268] * vector[4] +matrix[5][268] * vector[5] +matrix[6][268] * vector[6] +matrix[7][268] * vector[7] +matrix[8][268] * vector[8] +matrix[9][268] * vector[9] +matrix[10][268] * vector[10] +matrix[11][268] * vector[11] +matrix[12][268] * vector[12] +matrix[13][268] * vector[13] +matrix[14][268] * vector[14] +matrix[15][268] * vector[15] +matrix[16][268] * vector[16] +matrix[17][268] * vector[17] +matrix[18][268] * vector[18] +matrix[19][268] * vector[19] +matrix[20][268] * vector[20] +matrix[21][268] * vector[21] +matrix[22][268] * vector[22] +matrix[23][268] * vector[23] +matrix[24][268] * vector[24] +matrix[25][268] * vector[25] +matrix[26][268] * vector[26] +matrix[27][268] * vector[27] +matrix[28][268] * vector[28] +matrix[29][268] * vector[29] +matrix[30][268] * vector[30] +matrix[31][268] * vector[31] +matrix[32][268] * vector[32] +matrix[33][268] * vector[33] +matrix[34][268] * vector[34] +matrix[35][268] * vector[35] +matrix[36][268] * vector[36] +matrix[37][268] * vector[37] +matrix[38][268] * vector[38] +matrix[39][268] * vector[39] +matrix[40][268] * vector[40] +matrix[41][268] * vector[41] +matrix[42][268] * vector[42] +matrix[43][268] * vector[43] +matrix[44][268] * vector[44] +matrix[45][268] * vector[45] +matrix[46][268] * vector[46] +matrix[47][268] * vector[47] +matrix[48][268] * vector[48] +matrix[49][268] * vector[49] +matrix[50][268] * vector[50] +matrix[51][268] * vector[51] +matrix[52][268] * vector[52] +matrix[53][268] * vector[53] +matrix[54][268] * vector[54] +matrix[55][268] * vector[55] +matrix[56][268] * vector[56] +matrix[57][268] * vector[57] +matrix[58][268] * vector[58] +matrix[59][268] * vector[59] +matrix[60][268] * vector[60] +matrix[61][268] * vector[61] +matrix[62][268] * vector[62] +matrix[63][268] * vector[63] +matrix[64][268] * vector[64] +matrix[65][268] * vector[65] +matrix[66][268] * vector[66] +matrix[67][268] * vector[67] +matrix[68][268] * vector[68] +matrix[69][268] * vector[69] +matrix[70][268] * vector[70] +matrix[71][268] * vector[71] +matrix[72][268] * vector[72] +matrix[73][268] * vector[73] +matrix[74][268] * vector[74] +matrix[75][268] * vector[75] +matrix[76][268] * vector[76] +matrix[77][268] * vector[77] +matrix[78][268] * vector[78] +matrix[79][268] * vector[79] +matrix[80][268] * vector[80] +matrix[81][268] * vector[81] +matrix[82][268] * vector[82] +matrix[83][268] * vector[83] +matrix[84][268] * vector[84] +matrix[85][268] * vector[85] +matrix[86][268] * vector[86] +matrix[87][268] * vector[87] +matrix[88][268] * vector[88] +matrix[89][268] * vector[89] +matrix[90][268] * vector[90] +matrix[91][268] * vector[91] +matrix[92][268] * vector[92] +matrix[93][268] * vector[93] +matrix[94][268] * vector[94] +matrix[95][268] * vector[95] +matrix[96][268] * vector[96] +matrix[97][268] * vector[97] +matrix[98][268] * vector[98] +matrix[99][268] * vector[99] +b[268];
assign result[269] = matrix[0][269] * vector[0] +matrix[1][269] * vector[1] +matrix[2][269] * vector[2] +matrix[3][269] * vector[3] +matrix[4][269] * vector[4] +matrix[5][269] * vector[5] +matrix[6][269] * vector[6] +matrix[7][269] * vector[7] +matrix[8][269] * vector[8] +matrix[9][269] * vector[9] +matrix[10][269] * vector[10] +matrix[11][269] * vector[11] +matrix[12][269] * vector[12] +matrix[13][269] * vector[13] +matrix[14][269] * vector[14] +matrix[15][269] * vector[15] +matrix[16][269] * vector[16] +matrix[17][269] * vector[17] +matrix[18][269] * vector[18] +matrix[19][269] * vector[19] +matrix[20][269] * vector[20] +matrix[21][269] * vector[21] +matrix[22][269] * vector[22] +matrix[23][269] * vector[23] +matrix[24][269] * vector[24] +matrix[25][269] * vector[25] +matrix[26][269] * vector[26] +matrix[27][269] * vector[27] +matrix[28][269] * vector[28] +matrix[29][269] * vector[29] +matrix[30][269] * vector[30] +matrix[31][269] * vector[31] +matrix[32][269] * vector[32] +matrix[33][269] * vector[33] +matrix[34][269] * vector[34] +matrix[35][269] * vector[35] +matrix[36][269] * vector[36] +matrix[37][269] * vector[37] +matrix[38][269] * vector[38] +matrix[39][269] * vector[39] +matrix[40][269] * vector[40] +matrix[41][269] * vector[41] +matrix[42][269] * vector[42] +matrix[43][269] * vector[43] +matrix[44][269] * vector[44] +matrix[45][269] * vector[45] +matrix[46][269] * vector[46] +matrix[47][269] * vector[47] +matrix[48][269] * vector[48] +matrix[49][269] * vector[49] +matrix[50][269] * vector[50] +matrix[51][269] * vector[51] +matrix[52][269] * vector[52] +matrix[53][269] * vector[53] +matrix[54][269] * vector[54] +matrix[55][269] * vector[55] +matrix[56][269] * vector[56] +matrix[57][269] * vector[57] +matrix[58][269] * vector[58] +matrix[59][269] * vector[59] +matrix[60][269] * vector[60] +matrix[61][269] * vector[61] +matrix[62][269] * vector[62] +matrix[63][269] * vector[63] +matrix[64][269] * vector[64] +matrix[65][269] * vector[65] +matrix[66][269] * vector[66] +matrix[67][269] * vector[67] +matrix[68][269] * vector[68] +matrix[69][269] * vector[69] +matrix[70][269] * vector[70] +matrix[71][269] * vector[71] +matrix[72][269] * vector[72] +matrix[73][269] * vector[73] +matrix[74][269] * vector[74] +matrix[75][269] * vector[75] +matrix[76][269] * vector[76] +matrix[77][269] * vector[77] +matrix[78][269] * vector[78] +matrix[79][269] * vector[79] +matrix[80][269] * vector[80] +matrix[81][269] * vector[81] +matrix[82][269] * vector[82] +matrix[83][269] * vector[83] +matrix[84][269] * vector[84] +matrix[85][269] * vector[85] +matrix[86][269] * vector[86] +matrix[87][269] * vector[87] +matrix[88][269] * vector[88] +matrix[89][269] * vector[89] +matrix[90][269] * vector[90] +matrix[91][269] * vector[91] +matrix[92][269] * vector[92] +matrix[93][269] * vector[93] +matrix[94][269] * vector[94] +matrix[95][269] * vector[95] +matrix[96][269] * vector[96] +matrix[97][269] * vector[97] +matrix[98][269] * vector[98] +matrix[99][269] * vector[99] +b[269];
assign result[270] = matrix[0][270] * vector[0] +matrix[1][270] * vector[1] +matrix[2][270] * vector[2] +matrix[3][270] * vector[3] +matrix[4][270] * vector[4] +matrix[5][270] * vector[5] +matrix[6][270] * vector[6] +matrix[7][270] * vector[7] +matrix[8][270] * vector[8] +matrix[9][270] * vector[9] +matrix[10][270] * vector[10] +matrix[11][270] * vector[11] +matrix[12][270] * vector[12] +matrix[13][270] * vector[13] +matrix[14][270] * vector[14] +matrix[15][270] * vector[15] +matrix[16][270] * vector[16] +matrix[17][270] * vector[17] +matrix[18][270] * vector[18] +matrix[19][270] * vector[19] +matrix[20][270] * vector[20] +matrix[21][270] * vector[21] +matrix[22][270] * vector[22] +matrix[23][270] * vector[23] +matrix[24][270] * vector[24] +matrix[25][270] * vector[25] +matrix[26][270] * vector[26] +matrix[27][270] * vector[27] +matrix[28][270] * vector[28] +matrix[29][270] * vector[29] +matrix[30][270] * vector[30] +matrix[31][270] * vector[31] +matrix[32][270] * vector[32] +matrix[33][270] * vector[33] +matrix[34][270] * vector[34] +matrix[35][270] * vector[35] +matrix[36][270] * vector[36] +matrix[37][270] * vector[37] +matrix[38][270] * vector[38] +matrix[39][270] * vector[39] +matrix[40][270] * vector[40] +matrix[41][270] * vector[41] +matrix[42][270] * vector[42] +matrix[43][270] * vector[43] +matrix[44][270] * vector[44] +matrix[45][270] * vector[45] +matrix[46][270] * vector[46] +matrix[47][270] * vector[47] +matrix[48][270] * vector[48] +matrix[49][270] * vector[49] +matrix[50][270] * vector[50] +matrix[51][270] * vector[51] +matrix[52][270] * vector[52] +matrix[53][270] * vector[53] +matrix[54][270] * vector[54] +matrix[55][270] * vector[55] +matrix[56][270] * vector[56] +matrix[57][270] * vector[57] +matrix[58][270] * vector[58] +matrix[59][270] * vector[59] +matrix[60][270] * vector[60] +matrix[61][270] * vector[61] +matrix[62][270] * vector[62] +matrix[63][270] * vector[63] +matrix[64][270] * vector[64] +matrix[65][270] * vector[65] +matrix[66][270] * vector[66] +matrix[67][270] * vector[67] +matrix[68][270] * vector[68] +matrix[69][270] * vector[69] +matrix[70][270] * vector[70] +matrix[71][270] * vector[71] +matrix[72][270] * vector[72] +matrix[73][270] * vector[73] +matrix[74][270] * vector[74] +matrix[75][270] * vector[75] +matrix[76][270] * vector[76] +matrix[77][270] * vector[77] +matrix[78][270] * vector[78] +matrix[79][270] * vector[79] +matrix[80][270] * vector[80] +matrix[81][270] * vector[81] +matrix[82][270] * vector[82] +matrix[83][270] * vector[83] +matrix[84][270] * vector[84] +matrix[85][270] * vector[85] +matrix[86][270] * vector[86] +matrix[87][270] * vector[87] +matrix[88][270] * vector[88] +matrix[89][270] * vector[89] +matrix[90][270] * vector[90] +matrix[91][270] * vector[91] +matrix[92][270] * vector[92] +matrix[93][270] * vector[93] +matrix[94][270] * vector[94] +matrix[95][270] * vector[95] +matrix[96][270] * vector[96] +matrix[97][270] * vector[97] +matrix[98][270] * vector[98] +matrix[99][270] * vector[99] +b[270];
assign result[271] = matrix[0][271] * vector[0] +matrix[1][271] * vector[1] +matrix[2][271] * vector[2] +matrix[3][271] * vector[3] +matrix[4][271] * vector[4] +matrix[5][271] * vector[5] +matrix[6][271] * vector[6] +matrix[7][271] * vector[7] +matrix[8][271] * vector[8] +matrix[9][271] * vector[9] +matrix[10][271] * vector[10] +matrix[11][271] * vector[11] +matrix[12][271] * vector[12] +matrix[13][271] * vector[13] +matrix[14][271] * vector[14] +matrix[15][271] * vector[15] +matrix[16][271] * vector[16] +matrix[17][271] * vector[17] +matrix[18][271] * vector[18] +matrix[19][271] * vector[19] +matrix[20][271] * vector[20] +matrix[21][271] * vector[21] +matrix[22][271] * vector[22] +matrix[23][271] * vector[23] +matrix[24][271] * vector[24] +matrix[25][271] * vector[25] +matrix[26][271] * vector[26] +matrix[27][271] * vector[27] +matrix[28][271] * vector[28] +matrix[29][271] * vector[29] +matrix[30][271] * vector[30] +matrix[31][271] * vector[31] +matrix[32][271] * vector[32] +matrix[33][271] * vector[33] +matrix[34][271] * vector[34] +matrix[35][271] * vector[35] +matrix[36][271] * vector[36] +matrix[37][271] * vector[37] +matrix[38][271] * vector[38] +matrix[39][271] * vector[39] +matrix[40][271] * vector[40] +matrix[41][271] * vector[41] +matrix[42][271] * vector[42] +matrix[43][271] * vector[43] +matrix[44][271] * vector[44] +matrix[45][271] * vector[45] +matrix[46][271] * vector[46] +matrix[47][271] * vector[47] +matrix[48][271] * vector[48] +matrix[49][271] * vector[49] +matrix[50][271] * vector[50] +matrix[51][271] * vector[51] +matrix[52][271] * vector[52] +matrix[53][271] * vector[53] +matrix[54][271] * vector[54] +matrix[55][271] * vector[55] +matrix[56][271] * vector[56] +matrix[57][271] * vector[57] +matrix[58][271] * vector[58] +matrix[59][271] * vector[59] +matrix[60][271] * vector[60] +matrix[61][271] * vector[61] +matrix[62][271] * vector[62] +matrix[63][271] * vector[63] +matrix[64][271] * vector[64] +matrix[65][271] * vector[65] +matrix[66][271] * vector[66] +matrix[67][271] * vector[67] +matrix[68][271] * vector[68] +matrix[69][271] * vector[69] +matrix[70][271] * vector[70] +matrix[71][271] * vector[71] +matrix[72][271] * vector[72] +matrix[73][271] * vector[73] +matrix[74][271] * vector[74] +matrix[75][271] * vector[75] +matrix[76][271] * vector[76] +matrix[77][271] * vector[77] +matrix[78][271] * vector[78] +matrix[79][271] * vector[79] +matrix[80][271] * vector[80] +matrix[81][271] * vector[81] +matrix[82][271] * vector[82] +matrix[83][271] * vector[83] +matrix[84][271] * vector[84] +matrix[85][271] * vector[85] +matrix[86][271] * vector[86] +matrix[87][271] * vector[87] +matrix[88][271] * vector[88] +matrix[89][271] * vector[89] +matrix[90][271] * vector[90] +matrix[91][271] * vector[91] +matrix[92][271] * vector[92] +matrix[93][271] * vector[93] +matrix[94][271] * vector[94] +matrix[95][271] * vector[95] +matrix[96][271] * vector[96] +matrix[97][271] * vector[97] +matrix[98][271] * vector[98] +matrix[99][271] * vector[99] +b[271];
assign result[272] = matrix[0][272] * vector[0] +matrix[1][272] * vector[1] +matrix[2][272] * vector[2] +matrix[3][272] * vector[3] +matrix[4][272] * vector[4] +matrix[5][272] * vector[5] +matrix[6][272] * vector[6] +matrix[7][272] * vector[7] +matrix[8][272] * vector[8] +matrix[9][272] * vector[9] +matrix[10][272] * vector[10] +matrix[11][272] * vector[11] +matrix[12][272] * vector[12] +matrix[13][272] * vector[13] +matrix[14][272] * vector[14] +matrix[15][272] * vector[15] +matrix[16][272] * vector[16] +matrix[17][272] * vector[17] +matrix[18][272] * vector[18] +matrix[19][272] * vector[19] +matrix[20][272] * vector[20] +matrix[21][272] * vector[21] +matrix[22][272] * vector[22] +matrix[23][272] * vector[23] +matrix[24][272] * vector[24] +matrix[25][272] * vector[25] +matrix[26][272] * vector[26] +matrix[27][272] * vector[27] +matrix[28][272] * vector[28] +matrix[29][272] * vector[29] +matrix[30][272] * vector[30] +matrix[31][272] * vector[31] +matrix[32][272] * vector[32] +matrix[33][272] * vector[33] +matrix[34][272] * vector[34] +matrix[35][272] * vector[35] +matrix[36][272] * vector[36] +matrix[37][272] * vector[37] +matrix[38][272] * vector[38] +matrix[39][272] * vector[39] +matrix[40][272] * vector[40] +matrix[41][272] * vector[41] +matrix[42][272] * vector[42] +matrix[43][272] * vector[43] +matrix[44][272] * vector[44] +matrix[45][272] * vector[45] +matrix[46][272] * vector[46] +matrix[47][272] * vector[47] +matrix[48][272] * vector[48] +matrix[49][272] * vector[49] +matrix[50][272] * vector[50] +matrix[51][272] * vector[51] +matrix[52][272] * vector[52] +matrix[53][272] * vector[53] +matrix[54][272] * vector[54] +matrix[55][272] * vector[55] +matrix[56][272] * vector[56] +matrix[57][272] * vector[57] +matrix[58][272] * vector[58] +matrix[59][272] * vector[59] +matrix[60][272] * vector[60] +matrix[61][272] * vector[61] +matrix[62][272] * vector[62] +matrix[63][272] * vector[63] +matrix[64][272] * vector[64] +matrix[65][272] * vector[65] +matrix[66][272] * vector[66] +matrix[67][272] * vector[67] +matrix[68][272] * vector[68] +matrix[69][272] * vector[69] +matrix[70][272] * vector[70] +matrix[71][272] * vector[71] +matrix[72][272] * vector[72] +matrix[73][272] * vector[73] +matrix[74][272] * vector[74] +matrix[75][272] * vector[75] +matrix[76][272] * vector[76] +matrix[77][272] * vector[77] +matrix[78][272] * vector[78] +matrix[79][272] * vector[79] +matrix[80][272] * vector[80] +matrix[81][272] * vector[81] +matrix[82][272] * vector[82] +matrix[83][272] * vector[83] +matrix[84][272] * vector[84] +matrix[85][272] * vector[85] +matrix[86][272] * vector[86] +matrix[87][272] * vector[87] +matrix[88][272] * vector[88] +matrix[89][272] * vector[89] +matrix[90][272] * vector[90] +matrix[91][272] * vector[91] +matrix[92][272] * vector[92] +matrix[93][272] * vector[93] +matrix[94][272] * vector[94] +matrix[95][272] * vector[95] +matrix[96][272] * vector[96] +matrix[97][272] * vector[97] +matrix[98][272] * vector[98] +matrix[99][272] * vector[99] +b[272];
assign result[273] = matrix[0][273] * vector[0] +matrix[1][273] * vector[1] +matrix[2][273] * vector[2] +matrix[3][273] * vector[3] +matrix[4][273] * vector[4] +matrix[5][273] * vector[5] +matrix[6][273] * vector[6] +matrix[7][273] * vector[7] +matrix[8][273] * vector[8] +matrix[9][273] * vector[9] +matrix[10][273] * vector[10] +matrix[11][273] * vector[11] +matrix[12][273] * vector[12] +matrix[13][273] * vector[13] +matrix[14][273] * vector[14] +matrix[15][273] * vector[15] +matrix[16][273] * vector[16] +matrix[17][273] * vector[17] +matrix[18][273] * vector[18] +matrix[19][273] * vector[19] +matrix[20][273] * vector[20] +matrix[21][273] * vector[21] +matrix[22][273] * vector[22] +matrix[23][273] * vector[23] +matrix[24][273] * vector[24] +matrix[25][273] * vector[25] +matrix[26][273] * vector[26] +matrix[27][273] * vector[27] +matrix[28][273] * vector[28] +matrix[29][273] * vector[29] +matrix[30][273] * vector[30] +matrix[31][273] * vector[31] +matrix[32][273] * vector[32] +matrix[33][273] * vector[33] +matrix[34][273] * vector[34] +matrix[35][273] * vector[35] +matrix[36][273] * vector[36] +matrix[37][273] * vector[37] +matrix[38][273] * vector[38] +matrix[39][273] * vector[39] +matrix[40][273] * vector[40] +matrix[41][273] * vector[41] +matrix[42][273] * vector[42] +matrix[43][273] * vector[43] +matrix[44][273] * vector[44] +matrix[45][273] * vector[45] +matrix[46][273] * vector[46] +matrix[47][273] * vector[47] +matrix[48][273] * vector[48] +matrix[49][273] * vector[49] +matrix[50][273] * vector[50] +matrix[51][273] * vector[51] +matrix[52][273] * vector[52] +matrix[53][273] * vector[53] +matrix[54][273] * vector[54] +matrix[55][273] * vector[55] +matrix[56][273] * vector[56] +matrix[57][273] * vector[57] +matrix[58][273] * vector[58] +matrix[59][273] * vector[59] +matrix[60][273] * vector[60] +matrix[61][273] * vector[61] +matrix[62][273] * vector[62] +matrix[63][273] * vector[63] +matrix[64][273] * vector[64] +matrix[65][273] * vector[65] +matrix[66][273] * vector[66] +matrix[67][273] * vector[67] +matrix[68][273] * vector[68] +matrix[69][273] * vector[69] +matrix[70][273] * vector[70] +matrix[71][273] * vector[71] +matrix[72][273] * vector[72] +matrix[73][273] * vector[73] +matrix[74][273] * vector[74] +matrix[75][273] * vector[75] +matrix[76][273] * vector[76] +matrix[77][273] * vector[77] +matrix[78][273] * vector[78] +matrix[79][273] * vector[79] +matrix[80][273] * vector[80] +matrix[81][273] * vector[81] +matrix[82][273] * vector[82] +matrix[83][273] * vector[83] +matrix[84][273] * vector[84] +matrix[85][273] * vector[85] +matrix[86][273] * vector[86] +matrix[87][273] * vector[87] +matrix[88][273] * vector[88] +matrix[89][273] * vector[89] +matrix[90][273] * vector[90] +matrix[91][273] * vector[91] +matrix[92][273] * vector[92] +matrix[93][273] * vector[93] +matrix[94][273] * vector[94] +matrix[95][273] * vector[95] +matrix[96][273] * vector[96] +matrix[97][273] * vector[97] +matrix[98][273] * vector[98] +matrix[99][273] * vector[99] +b[273];
assign result[274] = matrix[0][274] * vector[0] +matrix[1][274] * vector[1] +matrix[2][274] * vector[2] +matrix[3][274] * vector[3] +matrix[4][274] * vector[4] +matrix[5][274] * vector[5] +matrix[6][274] * vector[6] +matrix[7][274] * vector[7] +matrix[8][274] * vector[8] +matrix[9][274] * vector[9] +matrix[10][274] * vector[10] +matrix[11][274] * vector[11] +matrix[12][274] * vector[12] +matrix[13][274] * vector[13] +matrix[14][274] * vector[14] +matrix[15][274] * vector[15] +matrix[16][274] * vector[16] +matrix[17][274] * vector[17] +matrix[18][274] * vector[18] +matrix[19][274] * vector[19] +matrix[20][274] * vector[20] +matrix[21][274] * vector[21] +matrix[22][274] * vector[22] +matrix[23][274] * vector[23] +matrix[24][274] * vector[24] +matrix[25][274] * vector[25] +matrix[26][274] * vector[26] +matrix[27][274] * vector[27] +matrix[28][274] * vector[28] +matrix[29][274] * vector[29] +matrix[30][274] * vector[30] +matrix[31][274] * vector[31] +matrix[32][274] * vector[32] +matrix[33][274] * vector[33] +matrix[34][274] * vector[34] +matrix[35][274] * vector[35] +matrix[36][274] * vector[36] +matrix[37][274] * vector[37] +matrix[38][274] * vector[38] +matrix[39][274] * vector[39] +matrix[40][274] * vector[40] +matrix[41][274] * vector[41] +matrix[42][274] * vector[42] +matrix[43][274] * vector[43] +matrix[44][274] * vector[44] +matrix[45][274] * vector[45] +matrix[46][274] * vector[46] +matrix[47][274] * vector[47] +matrix[48][274] * vector[48] +matrix[49][274] * vector[49] +matrix[50][274] * vector[50] +matrix[51][274] * vector[51] +matrix[52][274] * vector[52] +matrix[53][274] * vector[53] +matrix[54][274] * vector[54] +matrix[55][274] * vector[55] +matrix[56][274] * vector[56] +matrix[57][274] * vector[57] +matrix[58][274] * vector[58] +matrix[59][274] * vector[59] +matrix[60][274] * vector[60] +matrix[61][274] * vector[61] +matrix[62][274] * vector[62] +matrix[63][274] * vector[63] +matrix[64][274] * vector[64] +matrix[65][274] * vector[65] +matrix[66][274] * vector[66] +matrix[67][274] * vector[67] +matrix[68][274] * vector[68] +matrix[69][274] * vector[69] +matrix[70][274] * vector[70] +matrix[71][274] * vector[71] +matrix[72][274] * vector[72] +matrix[73][274] * vector[73] +matrix[74][274] * vector[74] +matrix[75][274] * vector[75] +matrix[76][274] * vector[76] +matrix[77][274] * vector[77] +matrix[78][274] * vector[78] +matrix[79][274] * vector[79] +matrix[80][274] * vector[80] +matrix[81][274] * vector[81] +matrix[82][274] * vector[82] +matrix[83][274] * vector[83] +matrix[84][274] * vector[84] +matrix[85][274] * vector[85] +matrix[86][274] * vector[86] +matrix[87][274] * vector[87] +matrix[88][274] * vector[88] +matrix[89][274] * vector[89] +matrix[90][274] * vector[90] +matrix[91][274] * vector[91] +matrix[92][274] * vector[92] +matrix[93][274] * vector[93] +matrix[94][274] * vector[94] +matrix[95][274] * vector[95] +matrix[96][274] * vector[96] +matrix[97][274] * vector[97] +matrix[98][274] * vector[98] +matrix[99][274] * vector[99] +b[274];
assign result[275] = matrix[0][275] * vector[0] +matrix[1][275] * vector[1] +matrix[2][275] * vector[2] +matrix[3][275] * vector[3] +matrix[4][275] * vector[4] +matrix[5][275] * vector[5] +matrix[6][275] * vector[6] +matrix[7][275] * vector[7] +matrix[8][275] * vector[8] +matrix[9][275] * vector[9] +matrix[10][275] * vector[10] +matrix[11][275] * vector[11] +matrix[12][275] * vector[12] +matrix[13][275] * vector[13] +matrix[14][275] * vector[14] +matrix[15][275] * vector[15] +matrix[16][275] * vector[16] +matrix[17][275] * vector[17] +matrix[18][275] * vector[18] +matrix[19][275] * vector[19] +matrix[20][275] * vector[20] +matrix[21][275] * vector[21] +matrix[22][275] * vector[22] +matrix[23][275] * vector[23] +matrix[24][275] * vector[24] +matrix[25][275] * vector[25] +matrix[26][275] * vector[26] +matrix[27][275] * vector[27] +matrix[28][275] * vector[28] +matrix[29][275] * vector[29] +matrix[30][275] * vector[30] +matrix[31][275] * vector[31] +matrix[32][275] * vector[32] +matrix[33][275] * vector[33] +matrix[34][275] * vector[34] +matrix[35][275] * vector[35] +matrix[36][275] * vector[36] +matrix[37][275] * vector[37] +matrix[38][275] * vector[38] +matrix[39][275] * vector[39] +matrix[40][275] * vector[40] +matrix[41][275] * vector[41] +matrix[42][275] * vector[42] +matrix[43][275] * vector[43] +matrix[44][275] * vector[44] +matrix[45][275] * vector[45] +matrix[46][275] * vector[46] +matrix[47][275] * vector[47] +matrix[48][275] * vector[48] +matrix[49][275] * vector[49] +matrix[50][275] * vector[50] +matrix[51][275] * vector[51] +matrix[52][275] * vector[52] +matrix[53][275] * vector[53] +matrix[54][275] * vector[54] +matrix[55][275] * vector[55] +matrix[56][275] * vector[56] +matrix[57][275] * vector[57] +matrix[58][275] * vector[58] +matrix[59][275] * vector[59] +matrix[60][275] * vector[60] +matrix[61][275] * vector[61] +matrix[62][275] * vector[62] +matrix[63][275] * vector[63] +matrix[64][275] * vector[64] +matrix[65][275] * vector[65] +matrix[66][275] * vector[66] +matrix[67][275] * vector[67] +matrix[68][275] * vector[68] +matrix[69][275] * vector[69] +matrix[70][275] * vector[70] +matrix[71][275] * vector[71] +matrix[72][275] * vector[72] +matrix[73][275] * vector[73] +matrix[74][275] * vector[74] +matrix[75][275] * vector[75] +matrix[76][275] * vector[76] +matrix[77][275] * vector[77] +matrix[78][275] * vector[78] +matrix[79][275] * vector[79] +matrix[80][275] * vector[80] +matrix[81][275] * vector[81] +matrix[82][275] * vector[82] +matrix[83][275] * vector[83] +matrix[84][275] * vector[84] +matrix[85][275] * vector[85] +matrix[86][275] * vector[86] +matrix[87][275] * vector[87] +matrix[88][275] * vector[88] +matrix[89][275] * vector[89] +matrix[90][275] * vector[90] +matrix[91][275] * vector[91] +matrix[92][275] * vector[92] +matrix[93][275] * vector[93] +matrix[94][275] * vector[94] +matrix[95][275] * vector[95] +matrix[96][275] * vector[96] +matrix[97][275] * vector[97] +matrix[98][275] * vector[98] +matrix[99][275] * vector[99] +b[275];
assign result[276] = matrix[0][276] * vector[0] +matrix[1][276] * vector[1] +matrix[2][276] * vector[2] +matrix[3][276] * vector[3] +matrix[4][276] * vector[4] +matrix[5][276] * vector[5] +matrix[6][276] * vector[6] +matrix[7][276] * vector[7] +matrix[8][276] * vector[8] +matrix[9][276] * vector[9] +matrix[10][276] * vector[10] +matrix[11][276] * vector[11] +matrix[12][276] * vector[12] +matrix[13][276] * vector[13] +matrix[14][276] * vector[14] +matrix[15][276] * vector[15] +matrix[16][276] * vector[16] +matrix[17][276] * vector[17] +matrix[18][276] * vector[18] +matrix[19][276] * vector[19] +matrix[20][276] * vector[20] +matrix[21][276] * vector[21] +matrix[22][276] * vector[22] +matrix[23][276] * vector[23] +matrix[24][276] * vector[24] +matrix[25][276] * vector[25] +matrix[26][276] * vector[26] +matrix[27][276] * vector[27] +matrix[28][276] * vector[28] +matrix[29][276] * vector[29] +matrix[30][276] * vector[30] +matrix[31][276] * vector[31] +matrix[32][276] * vector[32] +matrix[33][276] * vector[33] +matrix[34][276] * vector[34] +matrix[35][276] * vector[35] +matrix[36][276] * vector[36] +matrix[37][276] * vector[37] +matrix[38][276] * vector[38] +matrix[39][276] * vector[39] +matrix[40][276] * vector[40] +matrix[41][276] * vector[41] +matrix[42][276] * vector[42] +matrix[43][276] * vector[43] +matrix[44][276] * vector[44] +matrix[45][276] * vector[45] +matrix[46][276] * vector[46] +matrix[47][276] * vector[47] +matrix[48][276] * vector[48] +matrix[49][276] * vector[49] +matrix[50][276] * vector[50] +matrix[51][276] * vector[51] +matrix[52][276] * vector[52] +matrix[53][276] * vector[53] +matrix[54][276] * vector[54] +matrix[55][276] * vector[55] +matrix[56][276] * vector[56] +matrix[57][276] * vector[57] +matrix[58][276] * vector[58] +matrix[59][276] * vector[59] +matrix[60][276] * vector[60] +matrix[61][276] * vector[61] +matrix[62][276] * vector[62] +matrix[63][276] * vector[63] +matrix[64][276] * vector[64] +matrix[65][276] * vector[65] +matrix[66][276] * vector[66] +matrix[67][276] * vector[67] +matrix[68][276] * vector[68] +matrix[69][276] * vector[69] +matrix[70][276] * vector[70] +matrix[71][276] * vector[71] +matrix[72][276] * vector[72] +matrix[73][276] * vector[73] +matrix[74][276] * vector[74] +matrix[75][276] * vector[75] +matrix[76][276] * vector[76] +matrix[77][276] * vector[77] +matrix[78][276] * vector[78] +matrix[79][276] * vector[79] +matrix[80][276] * vector[80] +matrix[81][276] * vector[81] +matrix[82][276] * vector[82] +matrix[83][276] * vector[83] +matrix[84][276] * vector[84] +matrix[85][276] * vector[85] +matrix[86][276] * vector[86] +matrix[87][276] * vector[87] +matrix[88][276] * vector[88] +matrix[89][276] * vector[89] +matrix[90][276] * vector[90] +matrix[91][276] * vector[91] +matrix[92][276] * vector[92] +matrix[93][276] * vector[93] +matrix[94][276] * vector[94] +matrix[95][276] * vector[95] +matrix[96][276] * vector[96] +matrix[97][276] * vector[97] +matrix[98][276] * vector[98] +matrix[99][276] * vector[99] +b[276];
assign result[277] = matrix[0][277] * vector[0] +matrix[1][277] * vector[1] +matrix[2][277] * vector[2] +matrix[3][277] * vector[3] +matrix[4][277] * vector[4] +matrix[5][277] * vector[5] +matrix[6][277] * vector[6] +matrix[7][277] * vector[7] +matrix[8][277] * vector[8] +matrix[9][277] * vector[9] +matrix[10][277] * vector[10] +matrix[11][277] * vector[11] +matrix[12][277] * vector[12] +matrix[13][277] * vector[13] +matrix[14][277] * vector[14] +matrix[15][277] * vector[15] +matrix[16][277] * vector[16] +matrix[17][277] * vector[17] +matrix[18][277] * vector[18] +matrix[19][277] * vector[19] +matrix[20][277] * vector[20] +matrix[21][277] * vector[21] +matrix[22][277] * vector[22] +matrix[23][277] * vector[23] +matrix[24][277] * vector[24] +matrix[25][277] * vector[25] +matrix[26][277] * vector[26] +matrix[27][277] * vector[27] +matrix[28][277] * vector[28] +matrix[29][277] * vector[29] +matrix[30][277] * vector[30] +matrix[31][277] * vector[31] +matrix[32][277] * vector[32] +matrix[33][277] * vector[33] +matrix[34][277] * vector[34] +matrix[35][277] * vector[35] +matrix[36][277] * vector[36] +matrix[37][277] * vector[37] +matrix[38][277] * vector[38] +matrix[39][277] * vector[39] +matrix[40][277] * vector[40] +matrix[41][277] * vector[41] +matrix[42][277] * vector[42] +matrix[43][277] * vector[43] +matrix[44][277] * vector[44] +matrix[45][277] * vector[45] +matrix[46][277] * vector[46] +matrix[47][277] * vector[47] +matrix[48][277] * vector[48] +matrix[49][277] * vector[49] +matrix[50][277] * vector[50] +matrix[51][277] * vector[51] +matrix[52][277] * vector[52] +matrix[53][277] * vector[53] +matrix[54][277] * vector[54] +matrix[55][277] * vector[55] +matrix[56][277] * vector[56] +matrix[57][277] * vector[57] +matrix[58][277] * vector[58] +matrix[59][277] * vector[59] +matrix[60][277] * vector[60] +matrix[61][277] * vector[61] +matrix[62][277] * vector[62] +matrix[63][277] * vector[63] +matrix[64][277] * vector[64] +matrix[65][277] * vector[65] +matrix[66][277] * vector[66] +matrix[67][277] * vector[67] +matrix[68][277] * vector[68] +matrix[69][277] * vector[69] +matrix[70][277] * vector[70] +matrix[71][277] * vector[71] +matrix[72][277] * vector[72] +matrix[73][277] * vector[73] +matrix[74][277] * vector[74] +matrix[75][277] * vector[75] +matrix[76][277] * vector[76] +matrix[77][277] * vector[77] +matrix[78][277] * vector[78] +matrix[79][277] * vector[79] +matrix[80][277] * vector[80] +matrix[81][277] * vector[81] +matrix[82][277] * vector[82] +matrix[83][277] * vector[83] +matrix[84][277] * vector[84] +matrix[85][277] * vector[85] +matrix[86][277] * vector[86] +matrix[87][277] * vector[87] +matrix[88][277] * vector[88] +matrix[89][277] * vector[89] +matrix[90][277] * vector[90] +matrix[91][277] * vector[91] +matrix[92][277] * vector[92] +matrix[93][277] * vector[93] +matrix[94][277] * vector[94] +matrix[95][277] * vector[95] +matrix[96][277] * vector[96] +matrix[97][277] * vector[97] +matrix[98][277] * vector[98] +matrix[99][277] * vector[99] +b[277];
assign result[278] = matrix[0][278] * vector[0] +matrix[1][278] * vector[1] +matrix[2][278] * vector[2] +matrix[3][278] * vector[3] +matrix[4][278] * vector[4] +matrix[5][278] * vector[5] +matrix[6][278] * vector[6] +matrix[7][278] * vector[7] +matrix[8][278] * vector[8] +matrix[9][278] * vector[9] +matrix[10][278] * vector[10] +matrix[11][278] * vector[11] +matrix[12][278] * vector[12] +matrix[13][278] * vector[13] +matrix[14][278] * vector[14] +matrix[15][278] * vector[15] +matrix[16][278] * vector[16] +matrix[17][278] * vector[17] +matrix[18][278] * vector[18] +matrix[19][278] * vector[19] +matrix[20][278] * vector[20] +matrix[21][278] * vector[21] +matrix[22][278] * vector[22] +matrix[23][278] * vector[23] +matrix[24][278] * vector[24] +matrix[25][278] * vector[25] +matrix[26][278] * vector[26] +matrix[27][278] * vector[27] +matrix[28][278] * vector[28] +matrix[29][278] * vector[29] +matrix[30][278] * vector[30] +matrix[31][278] * vector[31] +matrix[32][278] * vector[32] +matrix[33][278] * vector[33] +matrix[34][278] * vector[34] +matrix[35][278] * vector[35] +matrix[36][278] * vector[36] +matrix[37][278] * vector[37] +matrix[38][278] * vector[38] +matrix[39][278] * vector[39] +matrix[40][278] * vector[40] +matrix[41][278] * vector[41] +matrix[42][278] * vector[42] +matrix[43][278] * vector[43] +matrix[44][278] * vector[44] +matrix[45][278] * vector[45] +matrix[46][278] * vector[46] +matrix[47][278] * vector[47] +matrix[48][278] * vector[48] +matrix[49][278] * vector[49] +matrix[50][278] * vector[50] +matrix[51][278] * vector[51] +matrix[52][278] * vector[52] +matrix[53][278] * vector[53] +matrix[54][278] * vector[54] +matrix[55][278] * vector[55] +matrix[56][278] * vector[56] +matrix[57][278] * vector[57] +matrix[58][278] * vector[58] +matrix[59][278] * vector[59] +matrix[60][278] * vector[60] +matrix[61][278] * vector[61] +matrix[62][278] * vector[62] +matrix[63][278] * vector[63] +matrix[64][278] * vector[64] +matrix[65][278] * vector[65] +matrix[66][278] * vector[66] +matrix[67][278] * vector[67] +matrix[68][278] * vector[68] +matrix[69][278] * vector[69] +matrix[70][278] * vector[70] +matrix[71][278] * vector[71] +matrix[72][278] * vector[72] +matrix[73][278] * vector[73] +matrix[74][278] * vector[74] +matrix[75][278] * vector[75] +matrix[76][278] * vector[76] +matrix[77][278] * vector[77] +matrix[78][278] * vector[78] +matrix[79][278] * vector[79] +matrix[80][278] * vector[80] +matrix[81][278] * vector[81] +matrix[82][278] * vector[82] +matrix[83][278] * vector[83] +matrix[84][278] * vector[84] +matrix[85][278] * vector[85] +matrix[86][278] * vector[86] +matrix[87][278] * vector[87] +matrix[88][278] * vector[88] +matrix[89][278] * vector[89] +matrix[90][278] * vector[90] +matrix[91][278] * vector[91] +matrix[92][278] * vector[92] +matrix[93][278] * vector[93] +matrix[94][278] * vector[94] +matrix[95][278] * vector[95] +matrix[96][278] * vector[96] +matrix[97][278] * vector[97] +matrix[98][278] * vector[98] +matrix[99][278] * vector[99] +b[278];
assign result[279] = matrix[0][279] * vector[0] +matrix[1][279] * vector[1] +matrix[2][279] * vector[2] +matrix[3][279] * vector[3] +matrix[4][279] * vector[4] +matrix[5][279] * vector[5] +matrix[6][279] * vector[6] +matrix[7][279] * vector[7] +matrix[8][279] * vector[8] +matrix[9][279] * vector[9] +matrix[10][279] * vector[10] +matrix[11][279] * vector[11] +matrix[12][279] * vector[12] +matrix[13][279] * vector[13] +matrix[14][279] * vector[14] +matrix[15][279] * vector[15] +matrix[16][279] * vector[16] +matrix[17][279] * vector[17] +matrix[18][279] * vector[18] +matrix[19][279] * vector[19] +matrix[20][279] * vector[20] +matrix[21][279] * vector[21] +matrix[22][279] * vector[22] +matrix[23][279] * vector[23] +matrix[24][279] * vector[24] +matrix[25][279] * vector[25] +matrix[26][279] * vector[26] +matrix[27][279] * vector[27] +matrix[28][279] * vector[28] +matrix[29][279] * vector[29] +matrix[30][279] * vector[30] +matrix[31][279] * vector[31] +matrix[32][279] * vector[32] +matrix[33][279] * vector[33] +matrix[34][279] * vector[34] +matrix[35][279] * vector[35] +matrix[36][279] * vector[36] +matrix[37][279] * vector[37] +matrix[38][279] * vector[38] +matrix[39][279] * vector[39] +matrix[40][279] * vector[40] +matrix[41][279] * vector[41] +matrix[42][279] * vector[42] +matrix[43][279] * vector[43] +matrix[44][279] * vector[44] +matrix[45][279] * vector[45] +matrix[46][279] * vector[46] +matrix[47][279] * vector[47] +matrix[48][279] * vector[48] +matrix[49][279] * vector[49] +matrix[50][279] * vector[50] +matrix[51][279] * vector[51] +matrix[52][279] * vector[52] +matrix[53][279] * vector[53] +matrix[54][279] * vector[54] +matrix[55][279] * vector[55] +matrix[56][279] * vector[56] +matrix[57][279] * vector[57] +matrix[58][279] * vector[58] +matrix[59][279] * vector[59] +matrix[60][279] * vector[60] +matrix[61][279] * vector[61] +matrix[62][279] * vector[62] +matrix[63][279] * vector[63] +matrix[64][279] * vector[64] +matrix[65][279] * vector[65] +matrix[66][279] * vector[66] +matrix[67][279] * vector[67] +matrix[68][279] * vector[68] +matrix[69][279] * vector[69] +matrix[70][279] * vector[70] +matrix[71][279] * vector[71] +matrix[72][279] * vector[72] +matrix[73][279] * vector[73] +matrix[74][279] * vector[74] +matrix[75][279] * vector[75] +matrix[76][279] * vector[76] +matrix[77][279] * vector[77] +matrix[78][279] * vector[78] +matrix[79][279] * vector[79] +matrix[80][279] * vector[80] +matrix[81][279] * vector[81] +matrix[82][279] * vector[82] +matrix[83][279] * vector[83] +matrix[84][279] * vector[84] +matrix[85][279] * vector[85] +matrix[86][279] * vector[86] +matrix[87][279] * vector[87] +matrix[88][279] * vector[88] +matrix[89][279] * vector[89] +matrix[90][279] * vector[90] +matrix[91][279] * vector[91] +matrix[92][279] * vector[92] +matrix[93][279] * vector[93] +matrix[94][279] * vector[94] +matrix[95][279] * vector[95] +matrix[96][279] * vector[96] +matrix[97][279] * vector[97] +matrix[98][279] * vector[98] +matrix[99][279] * vector[99] +b[279];
assign result[280] = matrix[0][280] * vector[0] +matrix[1][280] * vector[1] +matrix[2][280] * vector[2] +matrix[3][280] * vector[3] +matrix[4][280] * vector[4] +matrix[5][280] * vector[5] +matrix[6][280] * vector[6] +matrix[7][280] * vector[7] +matrix[8][280] * vector[8] +matrix[9][280] * vector[9] +matrix[10][280] * vector[10] +matrix[11][280] * vector[11] +matrix[12][280] * vector[12] +matrix[13][280] * vector[13] +matrix[14][280] * vector[14] +matrix[15][280] * vector[15] +matrix[16][280] * vector[16] +matrix[17][280] * vector[17] +matrix[18][280] * vector[18] +matrix[19][280] * vector[19] +matrix[20][280] * vector[20] +matrix[21][280] * vector[21] +matrix[22][280] * vector[22] +matrix[23][280] * vector[23] +matrix[24][280] * vector[24] +matrix[25][280] * vector[25] +matrix[26][280] * vector[26] +matrix[27][280] * vector[27] +matrix[28][280] * vector[28] +matrix[29][280] * vector[29] +matrix[30][280] * vector[30] +matrix[31][280] * vector[31] +matrix[32][280] * vector[32] +matrix[33][280] * vector[33] +matrix[34][280] * vector[34] +matrix[35][280] * vector[35] +matrix[36][280] * vector[36] +matrix[37][280] * vector[37] +matrix[38][280] * vector[38] +matrix[39][280] * vector[39] +matrix[40][280] * vector[40] +matrix[41][280] * vector[41] +matrix[42][280] * vector[42] +matrix[43][280] * vector[43] +matrix[44][280] * vector[44] +matrix[45][280] * vector[45] +matrix[46][280] * vector[46] +matrix[47][280] * vector[47] +matrix[48][280] * vector[48] +matrix[49][280] * vector[49] +matrix[50][280] * vector[50] +matrix[51][280] * vector[51] +matrix[52][280] * vector[52] +matrix[53][280] * vector[53] +matrix[54][280] * vector[54] +matrix[55][280] * vector[55] +matrix[56][280] * vector[56] +matrix[57][280] * vector[57] +matrix[58][280] * vector[58] +matrix[59][280] * vector[59] +matrix[60][280] * vector[60] +matrix[61][280] * vector[61] +matrix[62][280] * vector[62] +matrix[63][280] * vector[63] +matrix[64][280] * vector[64] +matrix[65][280] * vector[65] +matrix[66][280] * vector[66] +matrix[67][280] * vector[67] +matrix[68][280] * vector[68] +matrix[69][280] * vector[69] +matrix[70][280] * vector[70] +matrix[71][280] * vector[71] +matrix[72][280] * vector[72] +matrix[73][280] * vector[73] +matrix[74][280] * vector[74] +matrix[75][280] * vector[75] +matrix[76][280] * vector[76] +matrix[77][280] * vector[77] +matrix[78][280] * vector[78] +matrix[79][280] * vector[79] +matrix[80][280] * vector[80] +matrix[81][280] * vector[81] +matrix[82][280] * vector[82] +matrix[83][280] * vector[83] +matrix[84][280] * vector[84] +matrix[85][280] * vector[85] +matrix[86][280] * vector[86] +matrix[87][280] * vector[87] +matrix[88][280] * vector[88] +matrix[89][280] * vector[89] +matrix[90][280] * vector[90] +matrix[91][280] * vector[91] +matrix[92][280] * vector[92] +matrix[93][280] * vector[93] +matrix[94][280] * vector[94] +matrix[95][280] * vector[95] +matrix[96][280] * vector[96] +matrix[97][280] * vector[97] +matrix[98][280] * vector[98] +matrix[99][280] * vector[99] +b[280];
assign result[281] = matrix[0][281] * vector[0] +matrix[1][281] * vector[1] +matrix[2][281] * vector[2] +matrix[3][281] * vector[3] +matrix[4][281] * vector[4] +matrix[5][281] * vector[5] +matrix[6][281] * vector[6] +matrix[7][281] * vector[7] +matrix[8][281] * vector[8] +matrix[9][281] * vector[9] +matrix[10][281] * vector[10] +matrix[11][281] * vector[11] +matrix[12][281] * vector[12] +matrix[13][281] * vector[13] +matrix[14][281] * vector[14] +matrix[15][281] * vector[15] +matrix[16][281] * vector[16] +matrix[17][281] * vector[17] +matrix[18][281] * vector[18] +matrix[19][281] * vector[19] +matrix[20][281] * vector[20] +matrix[21][281] * vector[21] +matrix[22][281] * vector[22] +matrix[23][281] * vector[23] +matrix[24][281] * vector[24] +matrix[25][281] * vector[25] +matrix[26][281] * vector[26] +matrix[27][281] * vector[27] +matrix[28][281] * vector[28] +matrix[29][281] * vector[29] +matrix[30][281] * vector[30] +matrix[31][281] * vector[31] +matrix[32][281] * vector[32] +matrix[33][281] * vector[33] +matrix[34][281] * vector[34] +matrix[35][281] * vector[35] +matrix[36][281] * vector[36] +matrix[37][281] * vector[37] +matrix[38][281] * vector[38] +matrix[39][281] * vector[39] +matrix[40][281] * vector[40] +matrix[41][281] * vector[41] +matrix[42][281] * vector[42] +matrix[43][281] * vector[43] +matrix[44][281] * vector[44] +matrix[45][281] * vector[45] +matrix[46][281] * vector[46] +matrix[47][281] * vector[47] +matrix[48][281] * vector[48] +matrix[49][281] * vector[49] +matrix[50][281] * vector[50] +matrix[51][281] * vector[51] +matrix[52][281] * vector[52] +matrix[53][281] * vector[53] +matrix[54][281] * vector[54] +matrix[55][281] * vector[55] +matrix[56][281] * vector[56] +matrix[57][281] * vector[57] +matrix[58][281] * vector[58] +matrix[59][281] * vector[59] +matrix[60][281] * vector[60] +matrix[61][281] * vector[61] +matrix[62][281] * vector[62] +matrix[63][281] * vector[63] +matrix[64][281] * vector[64] +matrix[65][281] * vector[65] +matrix[66][281] * vector[66] +matrix[67][281] * vector[67] +matrix[68][281] * vector[68] +matrix[69][281] * vector[69] +matrix[70][281] * vector[70] +matrix[71][281] * vector[71] +matrix[72][281] * vector[72] +matrix[73][281] * vector[73] +matrix[74][281] * vector[74] +matrix[75][281] * vector[75] +matrix[76][281] * vector[76] +matrix[77][281] * vector[77] +matrix[78][281] * vector[78] +matrix[79][281] * vector[79] +matrix[80][281] * vector[80] +matrix[81][281] * vector[81] +matrix[82][281] * vector[82] +matrix[83][281] * vector[83] +matrix[84][281] * vector[84] +matrix[85][281] * vector[85] +matrix[86][281] * vector[86] +matrix[87][281] * vector[87] +matrix[88][281] * vector[88] +matrix[89][281] * vector[89] +matrix[90][281] * vector[90] +matrix[91][281] * vector[91] +matrix[92][281] * vector[92] +matrix[93][281] * vector[93] +matrix[94][281] * vector[94] +matrix[95][281] * vector[95] +matrix[96][281] * vector[96] +matrix[97][281] * vector[97] +matrix[98][281] * vector[98] +matrix[99][281] * vector[99] +b[281];
assign result[282] = matrix[0][282] * vector[0] +matrix[1][282] * vector[1] +matrix[2][282] * vector[2] +matrix[3][282] * vector[3] +matrix[4][282] * vector[4] +matrix[5][282] * vector[5] +matrix[6][282] * vector[6] +matrix[7][282] * vector[7] +matrix[8][282] * vector[8] +matrix[9][282] * vector[9] +matrix[10][282] * vector[10] +matrix[11][282] * vector[11] +matrix[12][282] * vector[12] +matrix[13][282] * vector[13] +matrix[14][282] * vector[14] +matrix[15][282] * vector[15] +matrix[16][282] * vector[16] +matrix[17][282] * vector[17] +matrix[18][282] * vector[18] +matrix[19][282] * vector[19] +matrix[20][282] * vector[20] +matrix[21][282] * vector[21] +matrix[22][282] * vector[22] +matrix[23][282] * vector[23] +matrix[24][282] * vector[24] +matrix[25][282] * vector[25] +matrix[26][282] * vector[26] +matrix[27][282] * vector[27] +matrix[28][282] * vector[28] +matrix[29][282] * vector[29] +matrix[30][282] * vector[30] +matrix[31][282] * vector[31] +matrix[32][282] * vector[32] +matrix[33][282] * vector[33] +matrix[34][282] * vector[34] +matrix[35][282] * vector[35] +matrix[36][282] * vector[36] +matrix[37][282] * vector[37] +matrix[38][282] * vector[38] +matrix[39][282] * vector[39] +matrix[40][282] * vector[40] +matrix[41][282] * vector[41] +matrix[42][282] * vector[42] +matrix[43][282] * vector[43] +matrix[44][282] * vector[44] +matrix[45][282] * vector[45] +matrix[46][282] * vector[46] +matrix[47][282] * vector[47] +matrix[48][282] * vector[48] +matrix[49][282] * vector[49] +matrix[50][282] * vector[50] +matrix[51][282] * vector[51] +matrix[52][282] * vector[52] +matrix[53][282] * vector[53] +matrix[54][282] * vector[54] +matrix[55][282] * vector[55] +matrix[56][282] * vector[56] +matrix[57][282] * vector[57] +matrix[58][282] * vector[58] +matrix[59][282] * vector[59] +matrix[60][282] * vector[60] +matrix[61][282] * vector[61] +matrix[62][282] * vector[62] +matrix[63][282] * vector[63] +matrix[64][282] * vector[64] +matrix[65][282] * vector[65] +matrix[66][282] * vector[66] +matrix[67][282] * vector[67] +matrix[68][282] * vector[68] +matrix[69][282] * vector[69] +matrix[70][282] * vector[70] +matrix[71][282] * vector[71] +matrix[72][282] * vector[72] +matrix[73][282] * vector[73] +matrix[74][282] * vector[74] +matrix[75][282] * vector[75] +matrix[76][282] * vector[76] +matrix[77][282] * vector[77] +matrix[78][282] * vector[78] +matrix[79][282] * vector[79] +matrix[80][282] * vector[80] +matrix[81][282] * vector[81] +matrix[82][282] * vector[82] +matrix[83][282] * vector[83] +matrix[84][282] * vector[84] +matrix[85][282] * vector[85] +matrix[86][282] * vector[86] +matrix[87][282] * vector[87] +matrix[88][282] * vector[88] +matrix[89][282] * vector[89] +matrix[90][282] * vector[90] +matrix[91][282] * vector[91] +matrix[92][282] * vector[92] +matrix[93][282] * vector[93] +matrix[94][282] * vector[94] +matrix[95][282] * vector[95] +matrix[96][282] * vector[96] +matrix[97][282] * vector[97] +matrix[98][282] * vector[98] +matrix[99][282] * vector[99] +b[282];
assign result[283] = matrix[0][283] * vector[0] +matrix[1][283] * vector[1] +matrix[2][283] * vector[2] +matrix[3][283] * vector[3] +matrix[4][283] * vector[4] +matrix[5][283] * vector[5] +matrix[6][283] * vector[6] +matrix[7][283] * vector[7] +matrix[8][283] * vector[8] +matrix[9][283] * vector[9] +matrix[10][283] * vector[10] +matrix[11][283] * vector[11] +matrix[12][283] * vector[12] +matrix[13][283] * vector[13] +matrix[14][283] * vector[14] +matrix[15][283] * vector[15] +matrix[16][283] * vector[16] +matrix[17][283] * vector[17] +matrix[18][283] * vector[18] +matrix[19][283] * vector[19] +matrix[20][283] * vector[20] +matrix[21][283] * vector[21] +matrix[22][283] * vector[22] +matrix[23][283] * vector[23] +matrix[24][283] * vector[24] +matrix[25][283] * vector[25] +matrix[26][283] * vector[26] +matrix[27][283] * vector[27] +matrix[28][283] * vector[28] +matrix[29][283] * vector[29] +matrix[30][283] * vector[30] +matrix[31][283] * vector[31] +matrix[32][283] * vector[32] +matrix[33][283] * vector[33] +matrix[34][283] * vector[34] +matrix[35][283] * vector[35] +matrix[36][283] * vector[36] +matrix[37][283] * vector[37] +matrix[38][283] * vector[38] +matrix[39][283] * vector[39] +matrix[40][283] * vector[40] +matrix[41][283] * vector[41] +matrix[42][283] * vector[42] +matrix[43][283] * vector[43] +matrix[44][283] * vector[44] +matrix[45][283] * vector[45] +matrix[46][283] * vector[46] +matrix[47][283] * vector[47] +matrix[48][283] * vector[48] +matrix[49][283] * vector[49] +matrix[50][283] * vector[50] +matrix[51][283] * vector[51] +matrix[52][283] * vector[52] +matrix[53][283] * vector[53] +matrix[54][283] * vector[54] +matrix[55][283] * vector[55] +matrix[56][283] * vector[56] +matrix[57][283] * vector[57] +matrix[58][283] * vector[58] +matrix[59][283] * vector[59] +matrix[60][283] * vector[60] +matrix[61][283] * vector[61] +matrix[62][283] * vector[62] +matrix[63][283] * vector[63] +matrix[64][283] * vector[64] +matrix[65][283] * vector[65] +matrix[66][283] * vector[66] +matrix[67][283] * vector[67] +matrix[68][283] * vector[68] +matrix[69][283] * vector[69] +matrix[70][283] * vector[70] +matrix[71][283] * vector[71] +matrix[72][283] * vector[72] +matrix[73][283] * vector[73] +matrix[74][283] * vector[74] +matrix[75][283] * vector[75] +matrix[76][283] * vector[76] +matrix[77][283] * vector[77] +matrix[78][283] * vector[78] +matrix[79][283] * vector[79] +matrix[80][283] * vector[80] +matrix[81][283] * vector[81] +matrix[82][283] * vector[82] +matrix[83][283] * vector[83] +matrix[84][283] * vector[84] +matrix[85][283] * vector[85] +matrix[86][283] * vector[86] +matrix[87][283] * vector[87] +matrix[88][283] * vector[88] +matrix[89][283] * vector[89] +matrix[90][283] * vector[90] +matrix[91][283] * vector[91] +matrix[92][283] * vector[92] +matrix[93][283] * vector[93] +matrix[94][283] * vector[94] +matrix[95][283] * vector[95] +matrix[96][283] * vector[96] +matrix[97][283] * vector[97] +matrix[98][283] * vector[98] +matrix[99][283] * vector[99] +b[283];
assign result[284] = matrix[0][284] * vector[0] +matrix[1][284] * vector[1] +matrix[2][284] * vector[2] +matrix[3][284] * vector[3] +matrix[4][284] * vector[4] +matrix[5][284] * vector[5] +matrix[6][284] * vector[6] +matrix[7][284] * vector[7] +matrix[8][284] * vector[8] +matrix[9][284] * vector[9] +matrix[10][284] * vector[10] +matrix[11][284] * vector[11] +matrix[12][284] * vector[12] +matrix[13][284] * vector[13] +matrix[14][284] * vector[14] +matrix[15][284] * vector[15] +matrix[16][284] * vector[16] +matrix[17][284] * vector[17] +matrix[18][284] * vector[18] +matrix[19][284] * vector[19] +matrix[20][284] * vector[20] +matrix[21][284] * vector[21] +matrix[22][284] * vector[22] +matrix[23][284] * vector[23] +matrix[24][284] * vector[24] +matrix[25][284] * vector[25] +matrix[26][284] * vector[26] +matrix[27][284] * vector[27] +matrix[28][284] * vector[28] +matrix[29][284] * vector[29] +matrix[30][284] * vector[30] +matrix[31][284] * vector[31] +matrix[32][284] * vector[32] +matrix[33][284] * vector[33] +matrix[34][284] * vector[34] +matrix[35][284] * vector[35] +matrix[36][284] * vector[36] +matrix[37][284] * vector[37] +matrix[38][284] * vector[38] +matrix[39][284] * vector[39] +matrix[40][284] * vector[40] +matrix[41][284] * vector[41] +matrix[42][284] * vector[42] +matrix[43][284] * vector[43] +matrix[44][284] * vector[44] +matrix[45][284] * vector[45] +matrix[46][284] * vector[46] +matrix[47][284] * vector[47] +matrix[48][284] * vector[48] +matrix[49][284] * vector[49] +matrix[50][284] * vector[50] +matrix[51][284] * vector[51] +matrix[52][284] * vector[52] +matrix[53][284] * vector[53] +matrix[54][284] * vector[54] +matrix[55][284] * vector[55] +matrix[56][284] * vector[56] +matrix[57][284] * vector[57] +matrix[58][284] * vector[58] +matrix[59][284] * vector[59] +matrix[60][284] * vector[60] +matrix[61][284] * vector[61] +matrix[62][284] * vector[62] +matrix[63][284] * vector[63] +matrix[64][284] * vector[64] +matrix[65][284] * vector[65] +matrix[66][284] * vector[66] +matrix[67][284] * vector[67] +matrix[68][284] * vector[68] +matrix[69][284] * vector[69] +matrix[70][284] * vector[70] +matrix[71][284] * vector[71] +matrix[72][284] * vector[72] +matrix[73][284] * vector[73] +matrix[74][284] * vector[74] +matrix[75][284] * vector[75] +matrix[76][284] * vector[76] +matrix[77][284] * vector[77] +matrix[78][284] * vector[78] +matrix[79][284] * vector[79] +matrix[80][284] * vector[80] +matrix[81][284] * vector[81] +matrix[82][284] * vector[82] +matrix[83][284] * vector[83] +matrix[84][284] * vector[84] +matrix[85][284] * vector[85] +matrix[86][284] * vector[86] +matrix[87][284] * vector[87] +matrix[88][284] * vector[88] +matrix[89][284] * vector[89] +matrix[90][284] * vector[90] +matrix[91][284] * vector[91] +matrix[92][284] * vector[92] +matrix[93][284] * vector[93] +matrix[94][284] * vector[94] +matrix[95][284] * vector[95] +matrix[96][284] * vector[96] +matrix[97][284] * vector[97] +matrix[98][284] * vector[98] +matrix[99][284] * vector[99] +b[284];
assign result[285] = matrix[0][285] * vector[0] +matrix[1][285] * vector[1] +matrix[2][285] * vector[2] +matrix[3][285] * vector[3] +matrix[4][285] * vector[4] +matrix[5][285] * vector[5] +matrix[6][285] * vector[6] +matrix[7][285] * vector[7] +matrix[8][285] * vector[8] +matrix[9][285] * vector[9] +matrix[10][285] * vector[10] +matrix[11][285] * vector[11] +matrix[12][285] * vector[12] +matrix[13][285] * vector[13] +matrix[14][285] * vector[14] +matrix[15][285] * vector[15] +matrix[16][285] * vector[16] +matrix[17][285] * vector[17] +matrix[18][285] * vector[18] +matrix[19][285] * vector[19] +matrix[20][285] * vector[20] +matrix[21][285] * vector[21] +matrix[22][285] * vector[22] +matrix[23][285] * vector[23] +matrix[24][285] * vector[24] +matrix[25][285] * vector[25] +matrix[26][285] * vector[26] +matrix[27][285] * vector[27] +matrix[28][285] * vector[28] +matrix[29][285] * vector[29] +matrix[30][285] * vector[30] +matrix[31][285] * vector[31] +matrix[32][285] * vector[32] +matrix[33][285] * vector[33] +matrix[34][285] * vector[34] +matrix[35][285] * vector[35] +matrix[36][285] * vector[36] +matrix[37][285] * vector[37] +matrix[38][285] * vector[38] +matrix[39][285] * vector[39] +matrix[40][285] * vector[40] +matrix[41][285] * vector[41] +matrix[42][285] * vector[42] +matrix[43][285] * vector[43] +matrix[44][285] * vector[44] +matrix[45][285] * vector[45] +matrix[46][285] * vector[46] +matrix[47][285] * vector[47] +matrix[48][285] * vector[48] +matrix[49][285] * vector[49] +matrix[50][285] * vector[50] +matrix[51][285] * vector[51] +matrix[52][285] * vector[52] +matrix[53][285] * vector[53] +matrix[54][285] * vector[54] +matrix[55][285] * vector[55] +matrix[56][285] * vector[56] +matrix[57][285] * vector[57] +matrix[58][285] * vector[58] +matrix[59][285] * vector[59] +matrix[60][285] * vector[60] +matrix[61][285] * vector[61] +matrix[62][285] * vector[62] +matrix[63][285] * vector[63] +matrix[64][285] * vector[64] +matrix[65][285] * vector[65] +matrix[66][285] * vector[66] +matrix[67][285] * vector[67] +matrix[68][285] * vector[68] +matrix[69][285] * vector[69] +matrix[70][285] * vector[70] +matrix[71][285] * vector[71] +matrix[72][285] * vector[72] +matrix[73][285] * vector[73] +matrix[74][285] * vector[74] +matrix[75][285] * vector[75] +matrix[76][285] * vector[76] +matrix[77][285] * vector[77] +matrix[78][285] * vector[78] +matrix[79][285] * vector[79] +matrix[80][285] * vector[80] +matrix[81][285] * vector[81] +matrix[82][285] * vector[82] +matrix[83][285] * vector[83] +matrix[84][285] * vector[84] +matrix[85][285] * vector[85] +matrix[86][285] * vector[86] +matrix[87][285] * vector[87] +matrix[88][285] * vector[88] +matrix[89][285] * vector[89] +matrix[90][285] * vector[90] +matrix[91][285] * vector[91] +matrix[92][285] * vector[92] +matrix[93][285] * vector[93] +matrix[94][285] * vector[94] +matrix[95][285] * vector[95] +matrix[96][285] * vector[96] +matrix[97][285] * vector[97] +matrix[98][285] * vector[98] +matrix[99][285] * vector[99] +b[285];
assign result[286] = matrix[0][286] * vector[0] +matrix[1][286] * vector[1] +matrix[2][286] * vector[2] +matrix[3][286] * vector[3] +matrix[4][286] * vector[4] +matrix[5][286] * vector[5] +matrix[6][286] * vector[6] +matrix[7][286] * vector[7] +matrix[8][286] * vector[8] +matrix[9][286] * vector[9] +matrix[10][286] * vector[10] +matrix[11][286] * vector[11] +matrix[12][286] * vector[12] +matrix[13][286] * vector[13] +matrix[14][286] * vector[14] +matrix[15][286] * vector[15] +matrix[16][286] * vector[16] +matrix[17][286] * vector[17] +matrix[18][286] * vector[18] +matrix[19][286] * vector[19] +matrix[20][286] * vector[20] +matrix[21][286] * vector[21] +matrix[22][286] * vector[22] +matrix[23][286] * vector[23] +matrix[24][286] * vector[24] +matrix[25][286] * vector[25] +matrix[26][286] * vector[26] +matrix[27][286] * vector[27] +matrix[28][286] * vector[28] +matrix[29][286] * vector[29] +matrix[30][286] * vector[30] +matrix[31][286] * vector[31] +matrix[32][286] * vector[32] +matrix[33][286] * vector[33] +matrix[34][286] * vector[34] +matrix[35][286] * vector[35] +matrix[36][286] * vector[36] +matrix[37][286] * vector[37] +matrix[38][286] * vector[38] +matrix[39][286] * vector[39] +matrix[40][286] * vector[40] +matrix[41][286] * vector[41] +matrix[42][286] * vector[42] +matrix[43][286] * vector[43] +matrix[44][286] * vector[44] +matrix[45][286] * vector[45] +matrix[46][286] * vector[46] +matrix[47][286] * vector[47] +matrix[48][286] * vector[48] +matrix[49][286] * vector[49] +matrix[50][286] * vector[50] +matrix[51][286] * vector[51] +matrix[52][286] * vector[52] +matrix[53][286] * vector[53] +matrix[54][286] * vector[54] +matrix[55][286] * vector[55] +matrix[56][286] * vector[56] +matrix[57][286] * vector[57] +matrix[58][286] * vector[58] +matrix[59][286] * vector[59] +matrix[60][286] * vector[60] +matrix[61][286] * vector[61] +matrix[62][286] * vector[62] +matrix[63][286] * vector[63] +matrix[64][286] * vector[64] +matrix[65][286] * vector[65] +matrix[66][286] * vector[66] +matrix[67][286] * vector[67] +matrix[68][286] * vector[68] +matrix[69][286] * vector[69] +matrix[70][286] * vector[70] +matrix[71][286] * vector[71] +matrix[72][286] * vector[72] +matrix[73][286] * vector[73] +matrix[74][286] * vector[74] +matrix[75][286] * vector[75] +matrix[76][286] * vector[76] +matrix[77][286] * vector[77] +matrix[78][286] * vector[78] +matrix[79][286] * vector[79] +matrix[80][286] * vector[80] +matrix[81][286] * vector[81] +matrix[82][286] * vector[82] +matrix[83][286] * vector[83] +matrix[84][286] * vector[84] +matrix[85][286] * vector[85] +matrix[86][286] * vector[86] +matrix[87][286] * vector[87] +matrix[88][286] * vector[88] +matrix[89][286] * vector[89] +matrix[90][286] * vector[90] +matrix[91][286] * vector[91] +matrix[92][286] * vector[92] +matrix[93][286] * vector[93] +matrix[94][286] * vector[94] +matrix[95][286] * vector[95] +matrix[96][286] * vector[96] +matrix[97][286] * vector[97] +matrix[98][286] * vector[98] +matrix[99][286] * vector[99] +b[286];
assign result[287] = matrix[0][287] * vector[0] +matrix[1][287] * vector[1] +matrix[2][287] * vector[2] +matrix[3][287] * vector[3] +matrix[4][287] * vector[4] +matrix[5][287] * vector[5] +matrix[6][287] * vector[6] +matrix[7][287] * vector[7] +matrix[8][287] * vector[8] +matrix[9][287] * vector[9] +matrix[10][287] * vector[10] +matrix[11][287] * vector[11] +matrix[12][287] * vector[12] +matrix[13][287] * vector[13] +matrix[14][287] * vector[14] +matrix[15][287] * vector[15] +matrix[16][287] * vector[16] +matrix[17][287] * vector[17] +matrix[18][287] * vector[18] +matrix[19][287] * vector[19] +matrix[20][287] * vector[20] +matrix[21][287] * vector[21] +matrix[22][287] * vector[22] +matrix[23][287] * vector[23] +matrix[24][287] * vector[24] +matrix[25][287] * vector[25] +matrix[26][287] * vector[26] +matrix[27][287] * vector[27] +matrix[28][287] * vector[28] +matrix[29][287] * vector[29] +matrix[30][287] * vector[30] +matrix[31][287] * vector[31] +matrix[32][287] * vector[32] +matrix[33][287] * vector[33] +matrix[34][287] * vector[34] +matrix[35][287] * vector[35] +matrix[36][287] * vector[36] +matrix[37][287] * vector[37] +matrix[38][287] * vector[38] +matrix[39][287] * vector[39] +matrix[40][287] * vector[40] +matrix[41][287] * vector[41] +matrix[42][287] * vector[42] +matrix[43][287] * vector[43] +matrix[44][287] * vector[44] +matrix[45][287] * vector[45] +matrix[46][287] * vector[46] +matrix[47][287] * vector[47] +matrix[48][287] * vector[48] +matrix[49][287] * vector[49] +matrix[50][287] * vector[50] +matrix[51][287] * vector[51] +matrix[52][287] * vector[52] +matrix[53][287] * vector[53] +matrix[54][287] * vector[54] +matrix[55][287] * vector[55] +matrix[56][287] * vector[56] +matrix[57][287] * vector[57] +matrix[58][287] * vector[58] +matrix[59][287] * vector[59] +matrix[60][287] * vector[60] +matrix[61][287] * vector[61] +matrix[62][287] * vector[62] +matrix[63][287] * vector[63] +matrix[64][287] * vector[64] +matrix[65][287] * vector[65] +matrix[66][287] * vector[66] +matrix[67][287] * vector[67] +matrix[68][287] * vector[68] +matrix[69][287] * vector[69] +matrix[70][287] * vector[70] +matrix[71][287] * vector[71] +matrix[72][287] * vector[72] +matrix[73][287] * vector[73] +matrix[74][287] * vector[74] +matrix[75][287] * vector[75] +matrix[76][287] * vector[76] +matrix[77][287] * vector[77] +matrix[78][287] * vector[78] +matrix[79][287] * vector[79] +matrix[80][287] * vector[80] +matrix[81][287] * vector[81] +matrix[82][287] * vector[82] +matrix[83][287] * vector[83] +matrix[84][287] * vector[84] +matrix[85][287] * vector[85] +matrix[86][287] * vector[86] +matrix[87][287] * vector[87] +matrix[88][287] * vector[88] +matrix[89][287] * vector[89] +matrix[90][287] * vector[90] +matrix[91][287] * vector[91] +matrix[92][287] * vector[92] +matrix[93][287] * vector[93] +matrix[94][287] * vector[94] +matrix[95][287] * vector[95] +matrix[96][287] * vector[96] +matrix[97][287] * vector[97] +matrix[98][287] * vector[98] +matrix[99][287] * vector[99] +b[287];
assign result[288] = matrix[0][288] * vector[0] +matrix[1][288] * vector[1] +matrix[2][288] * vector[2] +matrix[3][288] * vector[3] +matrix[4][288] * vector[4] +matrix[5][288] * vector[5] +matrix[6][288] * vector[6] +matrix[7][288] * vector[7] +matrix[8][288] * vector[8] +matrix[9][288] * vector[9] +matrix[10][288] * vector[10] +matrix[11][288] * vector[11] +matrix[12][288] * vector[12] +matrix[13][288] * vector[13] +matrix[14][288] * vector[14] +matrix[15][288] * vector[15] +matrix[16][288] * vector[16] +matrix[17][288] * vector[17] +matrix[18][288] * vector[18] +matrix[19][288] * vector[19] +matrix[20][288] * vector[20] +matrix[21][288] * vector[21] +matrix[22][288] * vector[22] +matrix[23][288] * vector[23] +matrix[24][288] * vector[24] +matrix[25][288] * vector[25] +matrix[26][288] * vector[26] +matrix[27][288] * vector[27] +matrix[28][288] * vector[28] +matrix[29][288] * vector[29] +matrix[30][288] * vector[30] +matrix[31][288] * vector[31] +matrix[32][288] * vector[32] +matrix[33][288] * vector[33] +matrix[34][288] * vector[34] +matrix[35][288] * vector[35] +matrix[36][288] * vector[36] +matrix[37][288] * vector[37] +matrix[38][288] * vector[38] +matrix[39][288] * vector[39] +matrix[40][288] * vector[40] +matrix[41][288] * vector[41] +matrix[42][288] * vector[42] +matrix[43][288] * vector[43] +matrix[44][288] * vector[44] +matrix[45][288] * vector[45] +matrix[46][288] * vector[46] +matrix[47][288] * vector[47] +matrix[48][288] * vector[48] +matrix[49][288] * vector[49] +matrix[50][288] * vector[50] +matrix[51][288] * vector[51] +matrix[52][288] * vector[52] +matrix[53][288] * vector[53] +matrix[54][288] * vector[54] +matrix[55][288] * vector[55] +matrix[56][288] * vector[56] +matrix[57][288] * vector[57] +matrix[58][288] * vector[58] +matrix[59][288] * vector[59] +matrix[60][288] * vector[60] +matrix[61][288] * vector[61] +matrix[62][288] * vector[62] +matrix[63][288] * vector[63] +matrix[64][288] * vector[64] +matrix[65][288] * vector[65] +matrix[66][288] * vector[66] +matrix[67][288] * vector[67] +matrix[68][288] * vector[68] +matrix[69][288] * vector[69] +matrix[70][288] * vector[70] +matrix[71][288] * vector[71] +matrix[72][288] * vector[72] +matrix[73][288] * vector[73] +matrix[74][288] * vector[74] +matrix[75][288] * vector[75] +matrix[76][288] * vector[76] +matrix[77][288] * vector[77] +matrix[78][288] * vector[78] +matrix[79][288] * vector[79] +matrix[80][288] * vector[80] +matrix[81][288] * vector[81] +matrix[82][288] * vector[82] +matrix[83][288] * vector[83] +matrix[84][288] * vector[84] +matrix[85][288] * vector[85] +matrix[86][288] * vector[86] +matrix[87][288] * vector[87] +matrix[88][288] * vector[88] +matrix[89][288] * vector[89] +matrix[90][288] * vector[90] +matrix[91][288] * vector[91] +matrix[92][288] * vector[92] +matrix[93][288] * vector[93] +matrix[94][288] * vector[94] +matrix[95][288] * vector[95] +matrix[96][288] * vector[96] +matrix[97][288] * vector[97] +matrix[98][288] * vector[98] +matrix[99][288] * vector[99] +b[288];
assign result[289] = matrix[0][289] * vector[0] +matrix[1][289] * vector[1] +matrix[2][289] * vector[2] +matrix[3][289] * vector[3] +matrix[4][289] * vector[4] +matrix[5][289] * vector[5] +matrix[6][289] * vector[6] +matrix[7][289] * vector[7] +matrix[8][289] * vector[8] +matrix[9][289] * vector[9] +matrix[10][289] * vector[10] +matrix[11][289] * vector[11] +matrix[12][289] * vector[12] +matrix[13][289] * vector[13] +matrix[14][289] * vector[14] +matrix[15][289] * vector[15] +matrix[16][289] * vector[16] +matrix[17][289] * vector[17] +matrix[18][289] * vector[18] +matrix[19][289] * vector[19] +matrix[20][289] * vector[20] +matrix[21][289] * vector[21] +matrix[22][289] * vector[22] +matrix[23][289] * vector[23] +matrix[24][289] * vector[24] +matrix[25][289] * vector[25] +matrix[26][289] * vector[26] +matrix[27][289] * vector[27] +matrix[28][289] * vector[28] +matrix[29][289] * vector[29] +matrix[30][289] * vector[30] +matrix[31][289] * vector[31] +matrix[32][289] * vector[32] +matrix[33][289] * vector[33] +matrix[34][289] * vector[34] +matrix[35][289] * vector[35] +matrix[36][289] * vector[36] +matrix[37][289] * vector[37] +matrix[38][289] * vector[38] +matrix[39][289] * vector[39] +matrix[40][289] * vector[40] +matrix[41][289] * vector[41] +matrix[42][289] * vector[42] +matrix[43][289] * vector[43] +matrix[44][289] * vector[44] +matrix[45][289] * vector[45] +matrix[46][289] * vector[46] +matrix[47][289] * vector[47] +matrix[48][289] * vector[48] +matrix[49][289] * vector[49] +matrix[50][289] * vector[50] +matrix[51][289] * vector[51] +matrix[52][289] * vector[52] +matrix[53][289] * vector[53] +matrix[54][289] * vector[54] +matrix[55][289] * vector[55] +matrix[56][289] * vector[56] +matrix[57][289] * vector[57] +matrix[58][289] * vector[58] +matrix[59][289] * vector[59] +matrix[60][289] * vector[60] +matrix[61][289] * vector[61] +matrix[62][289] * vector[62] +matrix[63][289] * vector[63] +matrix[64][289] * vector[64] +matrix[65][289] * vector[65] +matrix[66][289] * vector[66] +matrix[67][289] * vector[67] +matrix[68][289] * vector[68] +matrix[69][289] * vector[69] +matrix[70][289] * vector[70] +matrix[71][289] * vector[71] +matrix[72][289] * vector[72] +matrix[73][289] * vector[73] +matrix[74][289] * vector[74] +matrix[75][289] * vector[75] +matrix[76][289] * vector[76] +matrix[77][289] * vector[77] +matrix[78][289] * vector[78] +matrix[79][289] * vector[79] +matrix[80][289] * vector[80] +matrix[81][289] * vector[81] +matrix[82][289] * vector[82] +matrix[83][289] * vector[83] +matrix[84][289] * vector[84] +matrix[85][289] * vector[85] +matrix[86][289] * vector[86] +matrix[87][289] * vector[87] +matrix[88][289] * vector[88] +matrix[89][289] * vector[89] +matrix[90][289] * vector[90] +matrix[91][289] * vector[91] +matrix[92][289] * vector[92] +matrix[93][289] * vector[93] +matrix[94][289] * vector[94] +matrix[95][289] * vector[95] +matrix[96][289] * vector[96] +matrix[97][289] * vector[97] +matrix[98][289] * vector[98] +matrix[99][289] * vector[99] +b[289];
assign result[290] = matrix[0][290] * vector[0] +matrix[1][290] * vector[1] +matrix[2][290] * vector[2] +matrix[3][290] * vector[3] +matrix[4][290] * vector[4] +matrix[5][290] * vector[5] +matrix[6][290] * vector[6] +matrix[7][290] * vector[7] +matrix[8][290] * vector[8] +matrix[9][290] * vector[9] +matrix[10][290] * vector[10] +matrix[11][290] * vector[11] +matrix[12][290] * vector[12] +matrix[13][290] * vector[13] +matrix[14][290] * vector[14] +matrix[15][290] * vector[15] +matrix[16][290] * vector[16] +matrix[17][290] * vector[17] +matrix[18][290] * vector[18] +matrix[19][290] * vector[19] +matrix[20][290] * vector[20] +matrix[21][290] * vector[21] +matrix[22][290] * vector[22] +matrix[23][290] * vector[23] +matrix[24][290] * vector[24] +matrix[25][290] * vector[25] +matrix[26][290] * vector[26] +matrix[27][290] * vector[27] +matrix[28][290] * vector[28] +matrix[29][290] * vector[29] +matrix[30][290] * vector[30] +matrix[31][290] * vector[31] +matrix[32][290] * vector[32] +matrix[33][290] * vector[33] +matrix[34][290] * vector[34] +matrix[35][290] * vector[35] +matrix[36][290] * vector[36] +matrix[37][290] * vector[37] +matrix[38][290] * vector[38] +matrix[39][290] * vector[39] +matrix[40][290] * vector[40] +matrix[41][290] * vector[41] +matrix[42][290] * vector[42] +matrix[43][290] * vector[43] +matrix[44][290] * vector[44] +matrix[45][290] * vector[45] +matrix[46][290] * vector[46] +matrix[47][290] * vector[47] +matrix[48][290] * vector[48] +matrix[49][290] * vector[49] +matrix[50][290] * vector[50] +matrix[51][290] * vector[51] +matrix[52][290] * vector[52] +matrix[53][290] * vector[53] +matrix[54][290] * vector[54] +matrix[55][290] * vector[55] +matrix[56][290] * vector[56] +matrix[57][290] * vector[57] +matrix[58][290] * vector[58] +matrix[59][290] * vector[59] +matrix[60][290] * vector[60] +matrix[61][290] * vector[61] +matrix[62][290] * vector[62] +matrix[63][290] * vector[63] +matrix[64][290] * vector[64] +matrix[65][290] * vector[65] +matrix[66][290] * vector[66] +matrix[67][290] * vector[67] +matrix[68][290] * vector[68] +matrix[69][290] * vector[69] +matrix[70][290] * vector[70] +matrix[71][290] * vector[71] +matrix[72][290] * vector[72] +matrix[73][290] * vector[73] +matrix[74][290] * vector[74] +matrix[75][290] * vector[75] +matrix[76][290] * vector[76] +matrix[77][290] * vector[77] +matrix[78][290] * vector[78] +matrix[79][290] * vector[79] +matrix[80][290] * vector[80] +matrix[81][290] * vector[81] +matrix[82][290] * vector[82] +matrix[83][290] * vector[83] +matrix[84][290] * vector[84] +matrix[85][290] * vector[85] +matrix[86][290] * vector[86] +matrix[87][290] * vector[87] +matrix[88][290] * vector[88] +matrix[89][290] * vector[89] +matrix[90][290] * vector[90] +matrix[91][290] * vector[91] +matrix[92][290] * vector[92] +matrix[93][290] * vector[93] +matrix[94][290] * vector[94] +matrix[95][290] * vector[95] +matrix[96][290] * vector[96] +matrix[97][290] * vector[97] +matrix[98][290] * vector[98] +matrix[99][290] * vector[99] +b[290];
assign result[291] = matrix[0][291] * vector[0] +matrix[1][291] * vector[1] +matrix[2][291] * vector[2] +matrix[3][291] * vector[3] +matrix[4][291] * vector[4] +matrix[5][291] * vector[5] +matrix[6][291] * vector[6] +matrix[7][291] * vector[7] +matrix[8][291] * vector[8] +matrix[9][291] * vector[9] +matrix[10][291] * vector[10] +matrix[11][291] * vector[11] +matrix[12][291] * vector[12] +matrix[13][291] * vector[13] +matrix[14][291] * vector[14] +matrix[15][291] * vector[15] +matrix[16][291] * vector[16] +matrix[17][291] * vector[17] +matrix[18][291] * vector[18] +matrix[19][291] * vector[19] +matrix[20][291] * vector[20] +matrix[21][291] * vector[21] +matrix[22][291] * vector[22] +matrix[23][291] * vector[23] +matrix[24][291] * vector[24] +matrix[25][291] * vector[25] +matrix[26][291] * vector[26] +matrix[27][291] * vector[27] +matrix[28][291] * vector[28] +matrix[29][291] * vector[29] +matrix[30][291] * vector[30] +matrix[31][291] * vector[31] +matrix[32][291] * vector[32] +matrix[33][291] * vector[33] +matrix[34][291] * vector[34] +matrix[35][291] * vector[35] +matrix[36][291] * vector[36] +matrix[37][291] * vector[37] +matrix[38][291] * vector[38] +matrix[39][291] * vector[39] +matrix[40][291] * vector[40] +matrix[41][291] * vector[41] +matrix[42][291] * vector[42] +matrix[43][291] * vector[43] +matrix[44][291] * vector[44] +matrix[45][291] * vector[45] +matrix[46][291] * vector[46] +matrix[47][291] * vector[47] +matrix[48][291] * vector[48] +matrix[49][291] * vector[49] +matrix[50][291] * vector[50] +matrix[51][291] * vector[51] +matrix[52][291] * vector[52] +matrix[53][291] * vector[53] +matrix[54][291] * vector[54] +matrix[55][291] * vector[55] +matrix[56][291] * vector[56] +matrix[57][291] * vector[57] +matrix[58][291] * vector[58] +matrix[59][291] * vector[59] +matrix[60][291] * vector[60] +matrix[61][291] * vector[61] +matrix[62][291] * vector[62] +matrix[63][291] * vector[63] +matrix[64][291] * vector[64] +matrix[65][291] * vector[65] +matrix[66][291] * vector[66] +matrix[67][291] * vector[67] +matrix[68][291] * vector[68] +matrix[69][291] * vector[69] +matrix[70][291] * vector[70] +matrix[71][291] * vector[71] +matrix[72][291] * vector[72] +matrix[73][291] * vector[73] +matrix[74][291] * vector[74] +matrix[75][291] * vector[75] +matrix[76][291] * vector[76] +matrix[77][291] * vector[77] +matrix[78][291] * vector[78] +matrix[79][291] * vector[79] +matrix[80][291] * vector[80] +matrix[81][291] * vector[81] +matrix[82][291] * vector[82] +matrix[83][291] * vector[83] +matrix[84][291] * vector[84] +matrix[85][291] * vector[85] +matrix[86][291] * vector[86] +matrix[87][291] * vector[87] +matrix[88][291] * vector[88] +matrix[89][291] * vector[89] +matrix[90][291] * vector[90] +matrix[91][291] * vector[91] +matrix[92][291] * vector[92] +matrix[93][291] * vector[93] +matrix[94][291] * vector[94] +matrix[95][291] * vector[95] +matrix[96][291] * vector[96] +matrix[97][291] * vector[97] +matrix[98][291] * vector[98] +matrix[99][291] * vector[99] +b[291];
assign result[292] = matrix[0][292] * vector[0] +matrix[1][292] * vector[1] +matrix[2][292] * vector[2] +matrix[3][292] * vector[3] +matrix[4][292] * vector[4] +matrix[5][292] * vector[5] +matrix[6][292] * vector[6] +matrix[7][292] * vector[7] +matrix[8][292] * vector[8] +matrix[9][292] * vector[9] +matrix[10][292] * vector[10] +matrix[11][292] * vector[11] +matrix[12][292] * vector[12] +matrix[13][292] * vector[13] +matrix[14][292] * vector[14] +matrix[15][292] * vector[15] +matrix[16][292] * vector[16] +matrix[17][292] * vector[17] +matrix[18][292] * vector[18] +matrix[19][292] * vector[19] +matrix[20][292] * vector[20] +matrix[21][292] * vector[21] +matrix[22][292] * vector[22] +matrix[23][292] * vector[23] +matrix[24][292] * vector[24] +matrix[25][292] * vector[25] +matrix[26][292] * vector[26] +matrix[27][292] * vector[27] +matrix[28][292] * vector[28] +matrix[29][292] * vector[29] +matrix[30][292] * vector[30] +matrix[31][292] * vector[31] +matrix[32][292] * vector[32] +matrix[33][292] * vector[33] +matrix[34][292] * vector[34] +matrix[35][292] * vector[35] +matrix[36][292] * vector[36] +matrix[37][292] * vector[37] +matrix[38][292] * vector[38] +matrix[39][292] * vector[39] +matrix[40][292] * vector[40] +matrix[41][292] * vector[41] +matrix[42][292] * vector[42] +matrix[43][292] * vector[43] +matrix[44][292] * vector[44] +matrix[45][292] * vector[45] +matrix[46][292] * vector[46] +matrix[47][292] * vector[47] +matrix[48][292] * vector[48] +matrix[49][292] * vector[49] +matrix[50][292] * vector[50] +matrix[51][292] * vector[51] +matrix[52][292] * vector[52] +matrix[53][292] * vector[53] +matrix[54][292] * vector[54] +matrix[55][292] * vector[55] +matrix[56][292] * vector[56] +matrix[57][292] * vector[57] +matrix[58][292] * vector[58] +matrix[59][292] * vector[59] +matrix[60][292] * vector[60] +matrix[61][292] * vector[61] +matrix[62][292] * vector[62] +matrix[63][292] * vector[63] +matrix[64][292] * vector[64] +matrix[65][292] * vector[65] +matrix[66][292] * vector[66] +matrix[67][292] * vector[67] +matrix[68][292] * vector[68] +matrix[69][292] * vector[69] +matrix[70][292] * vector[70] +matrix[71][292] * vector[71] +matrix[72][292] * vector[72] +matrix[73][292] * vector[73] +matrix[74][292] * vector[74] +matrix[75][292] * vector[75] +matrix[76][292] * vector[76] +matrix[77][292] * vector[77] +matrix[78][292] * vector[78] +matrix[79][292] * vector[79] +matrix[80][292] * vector[80] +matrix[81][292] * vector[81] +matrix[82][292] * vector[82] +matrix[83][292] * vector[83] +matrix[84][292] * vector[84] +matrix[85][292] * vector[85] +matrix[86][292] * vector[86] +matrix[87][292] * vector[87] +matrix[88][292] * vector[88] +matrix[89][292] * vector[89] +matrix[90][292] * vector[90] +matrix[91][292] * vector[91] +matrix[92][292] * vector[92] +matrix[93][292] * vector[93] +matrix[94][292] * vector[94] +matrix[95][292] * vector[95] +matrix[96][292] * vector[96] +matrix[97][292] * vector[97] +matrix[98][292] * vector[98] +matrix[99][292] * vector[99] +b[292];
assign result[293] = matrix[0][293] * vector[0] +matrix[1][293] * vector[1] +matrix[2][293] * vector[2] +matrix[3][293] * vector[3] +matrix[4][293] * vector[4] +matrix[5][293] * vector[5] +matrix[6][293] * vector[6] +matrix[7][293] * vector[7] +matrix[8][293] * vector[8] +matrix[9][293] * vector[9] +matrix[10][293] * vector[10] +matrix[11][293] * vector[11] +matrix[12][293] * vector[12] +matrix[13][293] * vector[13] +matrix[14][293] * vector[14] +matrix[15][293] * vector[15] +matrix[16][293] * vector[16] +matrix[17][293] * vector[17] +matrix[18][293] * vector[18] +matrix[19][293] * vector[19] +matrix[20][293] * vector[20] +matrix[21][293] * vector[21] +matrix[22][293] * vector[22] +matrix[23][293] * vector[23] +matrix[24][293] * vector[24] +matrix[25][293] * vector[25] +matrix[26][293] * vector[26] +matrix[27][293] * vector[27] +matrix[28][293] * vector[28] +matrix[29][293] * vector[29] +matrix[30][293] * vector[30] +matrix[31][293] * vector[31] +matrix[32][293] * vector[32] +matrix[33][293] * vector[33] +matrix[34][293] * vector[34] +matrix[35][293] * vector[35] +matrix[36][293] * vector[36] +matrix[37][293] * vector[37] +matrix[38][293] * vector[38] +matrix[39][293] * vector[39] +matrix[40][293] * vector[40] +matrix[41][293] * vector[41] +matrix[42][293] * vector[42] +matrix[43][293] * vector[43] +matrix[44][293] * vector[44] +matrix[45][293] * vector[45] +matrix[46][293] * vector[46] +matrix[47][293] * vector[47] +matrix[48][293] * vector[48] +matrix[49][293] * vector[49] +matrix[50][293] * vector[50] +matrix[51][293] * vector[51] +matrix[52][293] * vector[52] +matrix[53][293] * vector[53] +matrix[54][293] * vector[54] +matrix[55][293] * vector[55] +matrix[56][293] * vector[56] +matrix[57][293] * vector[57] +matrix[58][293] * vector[58] +matrix[59][293] * vector[59] +matrix[60][293] * vector[60] +matrix[61][293] * vector[61] +matrix[62][293] * vector[62] +matrix[63][293] * vector[63] +matrix[64][293] * vector[64] +matrix[65][293] * vector[65] +matrix[66][293] * vector[66] +matrix[67][293] * vector[67] +matrix[68][293] * vector[68] +matrix[69][293] * vector[69] +matrix[70][293] * vector[70] +matrix[71][293] * vector[71] +matrix[72][293] * vector[72] +matrix[73][293] * vector[73] +matrix[74][293] * vector[74] +matrix[75][293] * vector[75] +matrix[76][293] * vector[76] +matrix[77][293] * vector[77] +matrix[78][293] * vector[78] +matrix[79][293] * vector[79] +matrix[80][293] * vector[80] +matrix[81][293] * vector[81] +matrix[82][293] * vector[82] +matrix[83][293] * vector[83] +matrix[84][293] * vector[84] +matrix[85][293] * vector[85] +matrix[86][293] * vector[86] +matrix[87][293] * vector[87] +matrix[88][293] * vector[88] +matrix[89][293] * vector[89] +matrix[90][293] * vector[90] +matrix[91][293] * vector[91] +matrix[92][293] * vector[92] +matrix[93][293] * vector[93] +matrix[94][293] * vector[94] +matrix[95][293] * vector[95] +matrix[96][293] * vector[96] +matrix[97][293] * vector[97] +matrix[98][293] * vector[98] +matrix[99][293] * vector[99] +b[293];
assign result[294] = matrix[0][294] * vector[0] +matrix[1][294] * vector[1] +matrix[2][294] * vector[2] +matrix[3][294] * vector[3] +matrix[4][294] * vector[4] +matrix[5][294] * vector[5] +matrix[6][294] * vector[6] +matrix[7][294] * vector[7] +matrix[8][294] * vector[8] +matrix[9][294] * vector[9] +matrix[10][294] * vector[10] +matrix[11][294] * vector[11] +matrix[12][294] * vector[12] +matrix[13][294] * vector[13] +matrix[14][294] * vector[14] +matrix[15][294] * vector[15] +matrix[16][294] * vector[16] +matrix[17][294] * vector[17] +matrix[18][294] * vector[18] +matrix[19][294] * vector[19] +matrix[20][294] * vector[20] +matrix[21][294] * vector[21] +matrix[22][294] * vector[22] +matrix[23][294] * vector[23] +matrix[24][294] * vector[24] +matrix[25][294] * vector[25] +matrix[26][294] * vector[26] +matrix[27][294] * vector[27] +matrix[28][294] * vector[28] +matrix[29][294] * vector[29] +matrix[30][294] * vector[30] +matrix[31][294] * vector[31] +matrix[32][294] * vector[32] +matrix[33][294] * vector[33] +matrix[34][294] * vector[34] +matrix[35][294] * vector[35] +matrix[36][294] * vector[36] +matrix[37][294] * vector[37] +matrix[38][294] * vector[38] +matrix[39][294] * vector[39] +matrix[40][294] * vector[40] +matrix[41][294] * vector[41] +matrix[42][294] * vector[42] +matrix[43][294] * vector[43] +matrix[44][294] * vector[44] +matrix[45][294] * vector[45] +matrix[46][294] * vector[46] +matrix[47][294] * vector[47] +matrix[48][294] * vector[48] +matrix[49][294] * vector[49] +matrix[50][294] * vector[50] +matrix[51][294] * vector[51] +matrix[52][294] * vector[52] +matrix[53][294] * vector[53] +matrix[54][294] * vector[54] +matrix[55][294] * vector[55] +matrix[56][294] * vector[56] +matrix[57][294] * vector[57] +matrix[58][294] * vector[58] +matrix[59][294] * vector[59] +matrix[60][294] * vector[60] +matrix[61][294] * vector[61] +matrix[62][294] * vector[62] +matrix[63][294] * vector[63] +matrix[64][294] * vector[64] +matrix[65][294] * vector[65] +matrix[66][294] * vector[66] +matrix[67][294] * vector[67] +matrix[68][294] * vector[68] +matrix[69][294] * vector[69] +matrix[70][294] * vector[70] +matrix[71][294] * vector[71] +matrix[72][294] * vector[72] +matrix[73][294] * vector[73] +matrix[74][294] * vector[74] +matrix[75][294] * vector[75] +matrix[76][294] * vector[76] +matrix[77][294] * vector[77] +matrix[78][294] * vector[78] +matrix[79][294] * vector[79] +matrix[80][294] * vector[80] +matrix[81][294] * vector[81] +matrix[82][294] * vector[82] +matrix[83][294] * vector[83] +matrix[84][294] * vector[84] +matrix[85][294] * vector[85] +matrix[86][294] * vector[86] +matrix[87][294] * vector[87] +matrix[88][294] * vector[88] +matrix[89][294] * vector[89] +matrix[90][294] * vector[90] +matrix[91][294] * vector[91] +matrix[92][294] * vector[92] +matrix[93][294] * vector[93] +matrix[94][294] * vector[94] +matrix[95][294] * vector[95] +matrix[96][294] * vector[96] +matrix[97][294] * vector[97] +matrix[98][294] * vector[98] +matrix[99][294] * vector[99] +b[294];
assign result[295] = matrix[0][295] * vector[0] +matrix[1][295] * vector[1] +matrix[2][295] * vector[2] +matrix[3][295] * vector[3] +matrix[4][295] * vector[4] +matrix[5][295] * vector[5] +matrix[6][295] * vector[6] +matrix[7][295] * vector[7] +matrix[8][295] * vector[8] +matrix[9][295] * vector[9] +matrix[10][295] * vector[10] +matrix[11][295] * vector[11] +matrix[12][295] * vector[12] +matrix[13][295] * vector[13] +matrix[14][295] * vector[14] +matrix[15][295] * vector[15] +matrix[16][295] * vector[16] +matrix[17][295] * vector[17] +matrix[18][295] * vector[18] +matrix[19][295] * vector[19] +matrix[20][295] * vector[20] +matrix[21][295] * vector[21] +matrix[22][295] * vector[22] +matrix[23][295] * vector[23] +matrix[24][295] * vector[24] +matrix[25][295] * vector[25] +matrix[26][295] * vector[26] +matrix[27][295] * vector[27] +matrix[28][295] * vector[28] +matrix[29][295] * vector[29] +matrix[30][295] * vector[30] +matrix[31][295] * vector[31] +matrix[32][295] * vector[32] +matrix[33][295] * vector[33] +matrix[34][295] * vector[34] +matrix[35][295] * vector[35] +matrix[36][295] * vector[36] +matrix[37][295] * vector[37] +matrix[38][295] * vector[38] +matrix[39][295] * vector[39] +matrix[40][295] * vector[40] +matrix[41][295] * vector[41] +matrix[42][295] * vector[42] +matrix[43][295] * vector[43] +matrix[44][295] * vector[44] +matrix[45][295] * vector[45] +matrix[46][295] * vector[46] +matrix[47][295] * vector[47] +matrix[48][295] * vector[48] +matrix[49][295] * vector[49] +matrix[50][295] * vector[50] +matrix[51][295] * vector[51] +matrix[52][295] * vector[52] +matrix[53][295] * vector[53] +matrix[54][295] * vector[54] +matrix[55][295] * vector[55] +matrix[56][295] * vector[56] +matrix[57][295] * vector[57] +matrix[58][295] * vector[58] +matrix[59][295] * vector[59] +matrix[60][295] * vector[60] +matrix[61][295] * vector[61] +matrix[62][295] * vector[62] +matrix[63][295] * vector[63] +matrix[64][295] * vector[64] +matrix[65][295] * vector[65] +matrix[66][295] * vector[66] +matrix[67][295] * vector[67] +matrix[68][295] * vector[68] +matrix[69][295] * vector[69] +matrix[70][295] * vector[70] +matrix[71][295] * vector[71] +matrix[72][295] * vector[72] +matrix[73][295] * vector[73] +matrix[74][295] * vector[74] +matrix[75][295] * vector[75] +matrix[76][295] * vector[76] +matrix[77][295] * vector[77] +matrix[78][295] * vector[78] +matrix[79][295] * vector[79] +matrix[80][295] * vector[80] +matrix[81][295] * vector[81] +matrix[82][295] * vector[82] +matrix[83][295] * vector[83] +matrix[84][295] * vector[84] +matrix[85][295] * vector[85] +matrix[86][295] * vector[86] +matrix[87][295] * vector[87] +matrix[88][295] * vector[88] +matrix[89][295] * vector[89] +matrix[90][295] * vector[90] +matrix[91][295] * vector[91] +matrix[92][295] * vector[92] +matrix[93][295] * vector[93] +matrix[94][295] * vector[94] +matrix[95][295] * vector[95] +matrix[96][295] * vector[96] +matrix[97][295] * vector[97] +matrix[98][295] * vector[98] +matrix[99][295] * vector[99] +b[295];
assign result[296] = matrix[0][296] * vector[0] +matrix[1][296] * vector[1] +matrix[2][296] * vector[2] +matrix[3][296] * vector[3] +matrix[4][296] * vector[4] +matrix[5][296] * vector[5] +matrix[6][296] * vector[6] +matrix[7][296] * vector[7] +matrix[8][296] * vector[8] +matrix[9][296] * vector[9] +matrix[10][296] * vector[10] +matrix[11][296] * vector[11] +matrix[12][296] * vector[12] +matrix[13][296] * vector[13] +matrix[14][296] * vector[14] +matrix[15][296] * vector[15] +matrix[16][296] * vector[16] +matrix[17][296] * vector[17] +matrix[18][296] * vector[18] +matrix[19][296] * vector[19] +matrix[20][296] * vector[20] +matrix[21][296] * vector[21] +matrix[22][296] * vector[22] +matrix[23][296] * vector[23] +matrix[24][296] * vector[24] +matrix[25][296] * vector[25] +matrix[26][296] * vector[26] +matrix[27][296] * vector[27] +matrix[28][296] * vector[28] +matrix[29][296] * vector[29] +matrix[30][296] * vector[30] +matrix[31][296] * vector[31] +matrix[32][296] * vector[32] +matrix[33][296] * vector[33] +matrix[34][296] * vector[34] +matrix[35][296] * vector[35] +matrix[36][296] * vector[36] +matrix[37][296] * vector[37] +matrix[38][296] * vector[38] +matrix[39][296] * vector[39] +matrix[40][296] * vector[40] +matrix[41][296] * vector[41] +matrix[42][296] * vector[42] +matrix[43][296] * vector[43] +matrix[44][296] * vector[44] +matrix[45][296] * vector[45] +matrix[46][296] * vector[46] +matrix[47][296] * vector[47] +matrix[48][296] * vector[48] +matrix[49][296] * vector[49] +matrix[50][296] * vector[50] +matrix[51][296] * vector[51] +matrix[52][296] * vector[52] +matrix[53][296] * vector[53] +matrix[54][296] * vector[54] +matrix[55][296] * vector[55] +matrix[56][296] * vector[56] +matrix[57][296] * vector[57] +matrix[58][296] * vector[58] +matrix[59][296] * vector[59] +matrix[60][296] * vector[60] +matrix[61][296] * vector[61] +matrix[62][296] * vector[62] +matrix[63][296] * vector[63] +matrix[64][296] * vector[64] +matrix[65][296] * vector[65] +matrix[66][296] * vector[66] +matrix[67][296] * vector[67] +matrix[68][296] * vector[68] +matrix[69][296] * vector[69] +matrix[70][296] * vector[70] +matrix[71][296] * vector[71] +matrix[72][296] * vector[72] +matrix[73][296] * vector[73] +matrix[74][296] * vector[74] +matrix[75][296] * vector[75] +matrix[76][296] * vector[76] +matrix[77][296] * vector[77] +matrix[78][296] * vector[78] +matrix[79][296] * vector[79] +matrix[80][296] * vector[80] +matrix[81][296] * vector[81] +matrix[82][296] * vector[82] +matrix[83][296] * vector[83] +matrix[84][296] * vector[84] +matrix[85][296] * vector[85] +matrix[86][296] * vector[86] +matrix[87][296] * vector[87] +matrix[88][296] * vector[88] +matrix[89][296] * vector[89] +matrix[90][296] * vector[90] +matrix[91][296] * vector[91] +matrix[92][296] * vector[92] +matrix[93][296] * vector[93] +matrix[94][296] * vector[94] +matrix[95][296] * vector[95] +matrix[96][296] * vector[96] +matrix[97][296] * vector[97] +matrix[98][296] * vector[98] +matrix[99][296] * vector[99] +b[296];
assign result[297] = matrix[0][297] * vector[0] +matrix[1][297] * vector[1] +matrix[2][297] * vector[2] +matrix[3][297] * vector[3] +matrix[4][297] * vector[4] +matrix[5][297] * vector[5] +matrix[6][297] * vector[6] +matrix[7][297] * vector[7] +matrix[8][297] * vector[8] +matrix[9][297] * vector[9] +matrix[10][297] * vector[10] +matrix[11][297] * vector[11] +matrix[12][297] * vector[12] +matrix[13][297] * vector[13] +matrix[14][297] * vector[14] +matrix[15][297] * vector[15] +matrix[16][297] * vector[16] +matrix[17][297] * vector[17] +matrix[18][297] * vector[18] +matrix[19][297] * vector[19] +matrix[20][297] * vector[20] +matrix[21][297] * vector[21] +matrix[22][297] * vector[22] +matrix[23][297] * vector[23] +matrix[24][297] * vector[24] +matrix[25][297] * vector[25] +matrix[26][297] * vector[26] +matrix[27][297] * vector[27] +matrix[28][297] * vector[28] +matrix[29][297] * vector[29] +matrix[30][297] * vector[30] +matrix[31][297] * vector[31] +matrix[32][297] * vector[32] +matrix[33][297] * vector[33] +matrix[34][297] * vector[34] +matrix[35][297] * vector[35] +matrix[36][297] * vector[36] +matrix[37][297] * vector[37] +matrix[38][297] * vector[38] +matrix[39][297] * vector[39] +matrix[40][297] * vector[40] +matrix[41][297] * vector[41] +matrix[42][297] * vector[42] +matrix[43][297] * vector[43] +matrix[44][297] * vector[44] +matrix[45][297] * vector[45] +matrix[46][297] * vector[46] +matrix[47][297] * vector[47] +matrix[48][297] * vector[48] +matrix[49][297] * vector[49] +matrix[50][297] * vector[50] +matrix[51][297] * vector[51] +matrix[52][297] * vector[52] +matrix[53][297] * vector[53] +matrix[54][297] * vector[54] +matrix[55][297] * vector[55] +matrix[56][297] * vector[56] +matrix[57][297] * vector[57] +matrix[58][297] * vector[58] +matrix[59][297] * vector[59] +matrix[60][297] * vector[60] +matrix[61][297] * vector[61] +matrix[62][297] * vector[62] +matrix[63][297] * vector[63] +matrix[64][297] * vector[64] +matrix[65][297] * vector[65] +matrix[66][297] * vector[66] +matrix[67][297] * vector[67] +matrix[68][297] * vector[68] +matrix[69][297] * vector[69] +matrix[70][297] * vector[70] +matrix[71][297] * vector[71] +matrix[72][297] * vector[72] +matrix[73][297] * vector[73] +matrix[74][297] * vector[74] +matrix[75][297] * vector[75] +matrix[76][297] * vector[76] +matrix[77][297] * vector[77] +matrix[78][297] * vector[78] +matrix[79][297] * vector[79] +matrix[80][297] * vector[80] +matrix[81][297] * vector[81] +matrix[82][297] * vector[82] +matrix[83][297] * vector[83] +matrix[84][297] * vector[84] +matrix[85][297] * vector[85] +matrix[86][297] * vector[86] +matrix[87][297] * vector[87] +matrix[88][297] * vector[88] +matrix[89][297] * vector[89] +matrix[90][297] * vector[90] +matrix[91][297] * vector[91] +matrix[92][297] * vector[92] +matrix[93][297] * vector[93] +matrix[94][297] * vector[94] +matrix[95][297] * vector[95] +matrix[96][297] * vector[96] +matrix[97][297] * vector[97] +matrix[98][297] * vector[98] +matrix[99][297] * vector[99] +b[297];
assign result[298] = matrix[0][298] * vector[0] +matrix[1][298] * vector[1] +matrix[2][298] * vector[2] +matrix[3][298] * vector[3] +matrix[4][298] * vector[4] +matrix[5][298] * vector[5] +matrix[6][298] * vector[6] +matrix[7][298] * vector[7] +matrix[8][298] * vector[8] +matrix[9][298] * vector[9] +matrix[10][298] * vector[10] +matrix[11][298] * vector[11] +matrix[12][298] * vector[12] +matrix[13][298] * vector[13] +matrix[14][298] * vector[14] +matrix[15][298] * vector[15] +matrix[16][298] * vector[16] +matrix[17][298] * vector[17] +matrix[18][298] * vector[18] +matrix[19][298] * vector[19] +matrix[20][298] * vector[20] +matrix[21][298] * vector[21] +matrix[22][298] * vector[22] +matrix[23][298] * vector[23] +matrix[24][298] * vector[24] +matrix[25][298] * vector[25] +matrix[26][298] * vector[26] +matrix[27][298] * vector[27] +matrix[28][298] * vector[28] +matrix[29][298] * vector[29] +matrix[30][298] * vector[30] +matrix[31][298] * vector[31] +matrix[32][298] * vector[32] +matrix[33][298] * vector[33] +matrix[34][298] * vector[34] +matrix[35][298] * vector[35] +matrix[36][298] * vector[36] +matrix[37][298] * vector[37] +matrix[38][298] * vector[38] +matrix[39][298] * vector[39] +matrix[40][298] * vector[40] +matrix[41][298] * vector[41] +matrix[42][298] * vector[42] +matrix[43][298] * vector[43] +matrix[44][298] * vector[44] +matrix[45][298] * vector[45] +matrix[46][298] * vector[46] +matrix[47][298] * vector[47] +matrix[48][298] * vector[48] +matrix[49][298] * vector[49] +matrix[50][298] * vector[50] +matrix[51][298] * vector[51] +matrix[52][298] * vector[52] +matrix[53][298] * vector[53] +matrix[54][298] * vector[54] +matrix[55][298] * vector[55] +matrix[56][298] * vector[56] +matrix[57][298] * vector[57] +matrix[58][298] * vector[58] +matrix[59][298] * vector[59] +matrix[60][298] * vector[60] +matrix[61][298] * vector[61] +matrix[62][298] * vector[62] +matrix[63][298] * vector[63] +matrix[64][298] * vector[64] +matrix[65][298] * vector[65] +matrix[66][298] * vector[66] +matrix[67][298] * vector[67] +matrix[68][298] * vector[68] +matrix[69][298] * vector[69] +matrix[70][298] * vector[70] +matrix[71][298] * vector[71] +matrix[72][298] * vector[72] +matrix[73][298] * vector[73] +matrix[74][298] * vector[74] +matrix[75][298] * vector[75] +matrix[76][298] * vector[76] +matrix[77][298] * vector[77] +matrix[78][298] * vector[78] +matrix[79][298] * vector[79] +matrix[80][298] * vector[80] +matrix[81][298] * vector[81] +matrix[82][298] * vector[82] +matrix[83][298] * vector[83] +matrix[84][298] * vector[84] +matrix[85][298] * vector[85] +matrix[86][298] * vector[86] +matrix[87][298] * vector[87] +matrix[88][298] * vector[88] +matrix[89][298] * vector[89] +matrix[90][298] * vector[90] +matrix[91][298] * vector[91] +matrix[92][298] * vector[92] +matrix[93][298] * vector[93] +matrix[94][298] * vector[94] +matrix[95][298] * vector[95] +matrix[96][298] * vector[96] +matrix[97][298] * vector[97] +matrix[98][298] * vector[98] +matrix[99][298] * vector[99] +b[298];
assign result[299] = matrix[0][299] * vector[0] +matrix[1][299] * vector[1] +matrix[2][299] * vector[2] +matrix[3][299] * vector[3] +matrix[4][299] * vector[4] +matrix[5][299] * vector[5] +matrix[6][299] * vector[6] +matrix[7][299] * vector[7] +matrix[8][299] * vector[8] +matrix[9][299] * vector[9] +matrix[10][299] * vector[10] +matrix[11][299] * vector[11] +matrix[12][299] * vector[12] +matrix[13][299] * vector[13] +matrix[14][299] * vector[14] +matrix[15][299] * vector[15] +matrix[16][299] * vector[16] +matrix[17][299] * vector[17] +matrix[18][299] * vector[18] +matrix[19][299] * vector[19] +matrix[20][299] * vector[20] +matrix[21][299] * vector[21] +matrix[22][299] * vector[22] +matrix[23][299] * vector[23] +matrix[24][299] * vector[24] +matrix[25][299] * vector[25] +matrix[26][299] * vector[26] +matrix[27][299] * vector[27] +matrix[28][299] * vector[28] +matrix[29][299] * vector[29] +matrix[30][299] * vector[30] +matrix[31][299] * vector[31] +matrix[32][299] * vector[32] +matrix[33][299] * vector[33] +matrix[34][299] * vector[34] +matrix[35][299] * vector[35] +matrix[36][299] * vector[36] +matrix[37][299] * vector[37] +matrix[38][299] * vector[38] +matrix[39][299] * vector[39] +matrix[40][299] * vector[40] +matrix[41][299] * vector[41] +matrix[42][299] * vector[42] +matrix[43][299] * vector[43] +matrix[44][299] * vector[44] +matrix[45][299] * vector[45] +matrix[46][299] * vector[46] +matrix[47][299] * vector[47] +matrix[48][299] * vector[48] +matrix[49][299] * vector[49] +matrix[50][299] * vector[50] +matrix[51][299] * vector[51] +matrix[52][299] * vector[52] +matrix[53][299] * vector[53] +matrix[54][299] * vector[54] +matrix[55][299] * vector[55] +matrix[56][299] * vector[56] +matrix[57][299] * vector[57] +matrix[58][299] * vector[58] +matrix[59][299] * vector[59] +matrix[60][299] * vector[60] +matrix[61][299] * vector[61] +matrix[62][299] * vector[62] +matrix[63][299] * vector[63] +matrix[64][299] * vector[64] +matrix[65][299] * vector[65] +matrix[66][299] * vector[66] +matrix[67][299] * vector[67] +matrix[68][299] * vector[68] +matrix[69][299] * vector[69] +matrix[70][299] * vector[70] +matrix[71][299] * vector[71] +matrix[72][299] * vector[72] +matrix[73][299] * vector[73] +matrix[74][299] * vector[74] +matrix[75][299] * vector[75] +matrix[76][299] * vector[76] +matrix[77][299] * vector[77] +matrix[78][299] * vector[78] +matrix[79][299] * vector[79] +matrix[80][299] * vector[80] +matrix[81][299] * vector[81] +matrix[82][299] * vector[82] +matrix[83][299] * vector[83] +matrix[84][299] * vector[84] +matrix[85][299] * vector[85] +matrix[86][299] * vector[86] +matrix[87][299] * vector[87] +matrix[88][299] * vector[88] +matrix[89][299] * vector[89] +matrix[90][299] * vector[90] +matrix[91][299] * vector[91] +matrix[92][299] * vector[92] +matrix[93][299] * vector[93] +matrix[94][299] * vector[94] +matrix[95][299] * vector[95] +matrix[96][299] * vector[96] +matrix[97][299] * vector[97] +matrix[98][299] * vector[98] +matrix[99][299] * vector[99] +b[299];
assign result[300] = matrix[0][300] * vector[0] +matrix[1][300] * vector[1] +matrix[2][300] * vector[2] +matrix[3][300] * vector[3] +matrix[4][300] * vector[4] +matrix[5][300] * vector[5] +matrix[6][300] * vector[6] +matrix[7][300] * vector[7] +matrix[8][300] * vector[8] +matrix[9][300] * vector[9] +matrix[10][300] * vector[10] +matrix[11][300] * vector[11] +matrix[12][300] * vector[12] +matrix[13][300] * vector[13] +matrix[14][300] * vector[14] +matrix[15][300] * vector[15] +matrix[16][300] * vector[16] +matrix[17][300] * vector[17] +matrix[18][300] * vector[18] +matrix[19][300] * vector[19] +matrix[20][300] * vector[20] +matrix[21][300] * vector[21] +matrix[22][300] * vector[22] +matrix[23][300] * vector[23] +matrix[24][300] * vector[24] +matrix[25][300] * vector[25] +matrix[26][300] * vector[26] +matrix[27][300] * vector[27] +matrix[28][300] * vector[28] +matrix[29][300] * vector[29] +matrix[30][300] * vector[30] +matrix[31][300] * vector[31] +matrix[32][300] * vector[32] +matrix[33][300] * vector[33] +matrix[34][300] * vector[34] +matrix[35][300] * vector[35] +matrix[36][300] * vector[36] +matrix[37][300] * vector[37] +matrix[38][300] * vector[38] +matrix[39][300] * vector[39] +matrix[40][300] * vector[40] +matrix[41][300] * vector[41] +matrix[42][300] * vector[42] +matrix[43][300] * vector[43] +matrix[44][300] * vector[44] +matrix[45][300] * vector[45] +matrix[46][300] * vector[46] +matrix[47][300] * vector[47] +matrix[48][300] * vector[48] +matrix[49][300] * vector[49] +matrix[50][300] * vector[50] +matrix[51][300] * vector[51] +matrix[52][300] * vector[52] +matrix[53][300] * vector[53] +matrix[54][300] * vector[54] +matrix[55][300] * vector[55] +matrix[56][300] * vector[56] +matrix[57][300] * vector[57] +matrix[58][300] * vector[58] +matrix[59][300] * vector[59] +matrix[60][300] * vector[60] +matrix[61][300] * vector[61] +matrix[62][300] * vector[62] +matrix[63][300] * vector[63] +matrix[64][300] * vector[64] +matrix[65][300] * vector[65] +matrix[66][300] * vector[66] +matrix[67][300] * vector[67] +matrix[68][300] * vector[68] +matrix[69][300] * vector[69] +matrix[70][300] * vector[70] +matrix[71][300] * vector[71] +matrix[72][300] * vector[72] +matrix[73][300] * vector[73] +matrix[74][300] * vector[74] +matrix[75][300] * vector[75] +matrix[76][300] * vector[76] +matrix[77][300] * vector[77] +matrix[78][300] * vector[78] +matrix[79][300] * vector[79] +matrix[80][300] * vector[80] +matrix[81][300] * vector[81] +matrix[82][300] * vector[82] +matrix[83][300] * vector[83] +matrix[84][300] * vector[84] +matrix[85][300] * vector[85] +matrix[86][300] * vector[86] +matrix[87][300] * vector[87] +matrix[88][300] * vector[88] +matrix[89][300] * vector[89] +matrix[90][300] * vector[90] +matrix[91][300] * vector[91] +matrix[92][300] * vector[92] +matrix[93][300] * vector[93] +matrix[94][300] * vector[94] +matrix[95][300] * vector[95] +matrix[96][300] * vector[96] +matrix[97][300] * vector[97] +matrix[98][300] * vector[98] +matrix[99][300] * vector[99] +b[300];
assign result[301] = matrix[0][301] * vector[0] +matrix[1][301] * vector[1] +matrix[2][301] * vector[2] +matrix[3][301] * vector[3] +matrix[4][301] * vector[4] +matrix[5][301] * vector[5] +matrix[6][301] * vector[6] +matrix[7][301] * vector[7] +matrix[8][301] * vector[8] +matrix[9][301] * vector[9] +matrix[10][301] * vector[10] +matrix[11][301] * vector[11] +matrix[12][301] * vector[12] +matrix[13][301] * vector[13] +matrix[14][301] * vector[14] +matrix[15][301] * vector[15] +matrix[16][301] * vector[16] +matrix[17][301] * vector[17] +matrix[18][301] * vector[18] +matrix[19][301] * vector[19] +matrix[20][301] * vector[20] +matrix[21][301] * vector[21] +matrix[22][301] * vector[22] +matrix[23][301] * vector[23] +matrix[24][301] * vector[24] +matrix[25][301] * vector[25] +matrix[26][301] * vector[26] +matrix[27][301] * vector[27] +matrix[28][301] * vector[28] +matrix[29][301] * vector[29] +matrix[30][301] * vector[30] +matrix[31][301] * vector[31] +matrix[32][301] * vector[32] +matrix[33][301] * vector[33] +matrix[34][301] * vector[34] +matrix[35][301] * vector[35] +matrix[36][301] * vector[36] +matrix[37][301] * vector[37] +matrix[38][301] * vector[38] +matrix[39][301] * vector[39] +matrix[40][301] * vector[40] +matrix[41][301] * vector[41] +matrix[42][301] * vector[42] +matrix[43][301] * vector[43] +matrix[44][301] * vector[44] +matrix[45][301] * vector[45] +matrix[46][301] * vector[46] +matrix[47][301] * vector[47] +matrix[48][301] * vector[48] +matrix[49][301] * vector[49] +matrix[50][301] * vector[50] +matrix[51][301] * vector[51] +matrix[52][301] * vector[52] +matrix[53][301] * vector[53] +matrix[54][301] * vector[54] +matrix[55][301] * vector[55] +matrix[56][301] * vector[56] +matrix[57][301] * vector[57] +matrix[58][301] * vector[58] +matrix[59][301] * vector[59] +matrix[60][301] * vector[60] +matrix[61][301] * vector[61] +matrix[62][301] * vector[62] +matrix[63][301] * vector[63] +matrix[64][301] * vector[64] +matrix[65][301] * vector[65] +matrix[66][301] * vector[66] +matrix[67][301] * vector[67] +matrix[68][301] * vector[68] +matrix[69][301] * vector[69] +matrix[70][301] * vector[70] +matrix[71][301] * vector[71] +matrix[72][301] * vector[72] +matrix[73][301] * vector[73] +matrix[74][301] * vector[74] +matrix[75][301] * vector[75] +matrix[76][301] * vector[76] +matrix[77][301] * vector[77] +matrix[78][301] * vector[78] +matrix[79][301] * vector[79] +matrix[80][301] * vector[80] +matrix[81][301] * vector[81] +matrix[82][301] * vector[82] +matrix[83][301] * vector[83] +matrix[84][301] * vector[84] +matrix[85][301] * vector[85] +matrix[86][301] * vector[86] +matrix[87][301] * vector[87] +matrix[88][301] * vector[88] +matrix[89][301] * vector[89] +matrix[90][301] * vector[90] +matrix[91][301] * vector[91] +matrix[92][301] * vector[92] +matrix[93][301] * vector[93] +matrix[94][301] * vector[94] +matrix[95][301] * vector[95] +matrix[96][301] * vector[96] +matrix[97][301] * vector[97] +matrix[98][301] * vector[98] +matrix[99][301] * vector[99] +b[301];
assign result[302] = matrix[0][302] * vector[0] +matrix[1][302] * vector[1] +matrix[2][302] * vector[2] +matrix[3][302] * vector[3] +matrix[4][302] * vector[4] +matrix[5][302] * vector[5] +matrix[6][302] * vector[6] +matrix[7][302] * vector[7] +matrix[8][302] * vector[8] +matrix[9][302] * vector[9] +matrix[10][302] * vector[10] +matrix[11][302] * vector[11] +matrix[12][302] * vector[12] +matrix[13][302] * vector[13] +matrix[14][302] * vector[14] +matrix[15][302] * vector[15] +matrix[16][302] * vector[16] +matrix[17][302] * vector[17] +matrix[18][302] * vector[18] +matrix[19][302] * vector[19] +matrix[20][302] * vector[20] +matrix[21][302] * vector[21] +matrix[22][302] * vector[22] +matrix[23][302] * vector[23] +matrix[24][302] * vector[24] +matrix[25][302] * vector[25] +matrix[26][302] * vector[26] +matrix[27][302] * vector[27] +matrix[28][302] * vector[28] +matrix[29][302] * vector[29] +matrix[30][302] * vector[30] +matrix[31][302] * vector[31] +matrix[32][302] * vector[32] +matrix[33][302] * vector[33] +matrix[34][302] * vector[34] +matrix[35][302] * vector[35] +matrix[36][302] * vector[36] +matrix[37][302] * vector[37] +matrix[38][302] * vector[38] +matrix[39][302] * vector[39] +matrix[40][302] * vector[40] +matrix[41][302] * vector[41] +matrix[42][302] * vector[42] +matrix[43][302] * vector[43] +matrix[44][302] * vector[44] +matrix[45][302] * vector[45] +matrix[46][302] * vector[46] +matrix[47][302] * vector[47] +matrix[48][302] * vector[48] +matrix[49][302] * vector[49] +matrix[50][302] * vector[50] +matrix[51][302] * vector[51] +matrix[52][302] * vector[52] +matrix[53][302] * vector[53] +matrix[54][302] * vector[54] +matrix[55][302] * vector[55] +matrix[56][302] * vector[56] +matrix[57][302] * vector[57] +matrix[58][302] * vector[58] +matrix[59][302] * vector[59] +matrix[60][302] * vector[60] +matrix[61][302] * vector[61] +matrix[62][302] * vector[62] +matrix[63][302] * vector[63] +matrix[64][302] * vector[64] +matrix[65][302] * vector[65] +matrix[66][302] * vector[66] +matrix[67][302] * vector[67] +matrix[68][302] * vector[68] +matrix[69][302] * vector[69] +matrix[70][302] * vector[70] +matrix[71][302] * vector[71] +matrix[72][302] * vector[72] +matrix[73][302] * vector[73] +matrix[74][302] * vector[74] +matrix[75][302] * vector[75] +matrix[76][302] * vector[76] +matrix[77][302] * vector[77] +matrix[78][302] * vector[78] +matrix[79][302] * vector[79] +matrix[80][302] * vector[80] +matrix[81][302] * vector[81] +matrix[82][302] * vector[82] +matrix[83][302] * vector[83] +matrix[84][302] * vector[84] +matrix[85][302] * vector[85] +matrix[86][302] * vector[86] +matrix[87][302] * vector[87] +matrix[88][302] * vector[88] +matrix[89][302] * vector[89] +matrix[90][302] * vector[90] +matrix[91][302] * vector[91] +matrix[92][302] * vector[92] +matrix[93][302] * vector[93] +matrix[94][302] * vector[94] +matrix[95][302] * vector[95] +matrix[96][302] * vector[96] +matrix[97][302] * vector[97] +matrix[98][302] * vector[98] +matrix[99][302] * vector[99] +b[302];
assign result[303] = matrix[0][303] * vector[0] +matrix[1][303] * vector[1] +matrix[2][303] * vector[2] +matrix[3][303] * vector[3] +matrix[4][303] * vector[4] +matrix[5][303] * vector[5] +matrix[6][303] * vector[6] +matrix[7][303] * vector[7] +matrix[8][303] * vector[8] +matrix[9][303] * vector[9] +matrix[10][303] * vector[10] +matrix[11][303] * vector[11] +matrix[12][303] * vector[12] +matrix[13][303] * vector[13] +matrix[14][303] * vector[14] +matrix[15][303] * vector[15] +matrix[16][303] * vector[16] +matrix[17][303] * vector[17] +matrix[18][303] * vector[18] +matrix[19][303] * vector[19] +matrix[20][303] * vector[20] +matrix[21][303] * vector[21] +matrix[22][303] * vector[22] +matrix[23][303] * vector[23] +matrix[24][303] * vector[24] +matrix[25][303] * vector[25] +matrix[26][303] * vector[26] +matrix[27][303] * vector[27] +matrix[28][303] * vector[28] +matrix[29][303] * vector[29] +matrix[30][303] * vector[30] +matrix[31][303] * vector[31] +matrix[32][303] * vector[32] +matrix[33][303] * vector[33] +matrix[34][303] * vector[34] +matrix[35][303] * vector[35] +matrix[36][303] * vector[36] +matrix[37][303] * vector[37] +matrix[38][303] * vector[38] +matrix[39][303] * vector[39] +matrix[40][303] * vector[40] +matrix[41][303] * vector[41] +matrix[42][303] * vector[42] +matrix[43][303] * vector[43] +matrix[44][303] * vector[44] +matrix[45][303] * vector[45] +matrix[46][303] * vector[46] +matrix[47][303] * vector[47] +matrix[48][303] * vector[48] +matrix[49][303] * vector[49] +matrix[50][303] * vector[50] +matrix[51][303] * vector[51] +matrix[52][303] * vector[52] +matrix[53][303] * vector[53] +matrix[54][303] * vector[54] +matrix[55][303] * vector[55] +matrix[56][303] * vector[56] +matrix[57][303] * vector[57] +matrix[58][303] * vector[58] +matrix[59][303] * vector[59] +matrix[60][303] * vector[60] +matrix[61][303] * vector[61] +matrix[62][303] * vector[62] +matrix[63][303] * vector[63] +matrix[64][303] * vector[64] +matrix[65][303] * vector[65] +matrix[66][303] * vector[66] +matrix[67][303] * vector[67] +matrix[68][303] * vector[68] +matrix[69][303] * vector[69] +matrix[70][303] * vector[70] +matrix[71][303] * vector[71] +matrix[72][303] * vector[72] +matrix[73][303] * vector[73] +matrix[74][303] * vector[74] +matrix[75][303] * vector[75] +matrix[76][303] * vector[76] +matrix[77][303] * vector[77] +matrix[78][303] * vector[78] +matrix[79][303] * vector[79] +matrix[80][303] * vector[80] +matrix[81][303] * vector[81] +matrix[82][303] * vector[82] +matrix[83][303] * vector[83] +matrix[84][303] * vector[84] +matrix[85][303] * vector[85] +matrix[86][303] * vector[86] +matrix[87][303] * vector[87] +matrix[88][303] * vector[88] +matrix[89][303] * vector[89] +matrix[90][303] * vector[90] +matrix[91][303] * vector[91] +matrix[92][303] * vector[92] +matrix[93][303] * vector[93] +matrix[94][303] * vector[94] +matrix[95][303] * vector[95] +matrix[96][303] * vector[96] +matrix[97][303] * vector[97] +matrix[98][303] * vector[98] +matrix[99][303] * vector[99] +b[303];
assign result[304] = matrix[0][304] * vector[0] +matrix[1][304] * vector[1] +matrix[2][304] * vector[2] +matrix[3][304] * vector[3] +matrix[4][304] * vector[4] +matrix[5][304] * vector[5] +matrix[6][304] * vector[6] +matrix[7][304] * vector[7] +matrix[8][304] * vector[8] +matrix[9][304] * vector[9] +matrix[10][304] * vector[10] +matrix[11][304] * vector[11] +matrix[12][304] * vector[12] +matrix[13][304] * vector[13] +matrix[14][304] * vector[14] +matrix[15][304] * vector[15] +matrix[16][304] * vector[16] +matrix[17][304] * vector[17] +matrix[18][304] * vector[18] +matrix[19][304] * vector[19] +matrix[20][304] * vector[20] +matrix[21][304] * vector[21] +matrix[22][304] * vector[22] +matrix[23][304] * vector[23] +matrix[24][304] * vector[24] +matrix[25][304] * vector[25] +matrix[26][304] * vector[26] +matrix[27][304] * vector[27] +matrix[28][304] * vector[28] +matrix[29][304] * vector[29] +matrix[30][304] * vector[30] +matrix[31][304] * vector[31] +matrix[32][304] * vector[32] +matrix[33][304] * vector[33] +matrix[34][304] * vector[34] +matrix[35][304] * vector[35] +matrix[36][304] * vector[36] +matrix[37][304] * vector[37] +matrix[38][304] * vector[38] +matrix[39][304] * vector[39] +matrix[40][304] * vector[40] +matrix[41][304] * vector[41] +matrix[42][304] * vector[42] +matrix[43][304] * vector[43] +matrix[44][304] * vector[44] +matrix[45][304] * vector[45] +matrix[46][304] * vector[46] +matrix[47][304] * vector[47] +matrix[48][304] * vector[48] +matrix[49][304] * vector[49] +matrix[50][304] * vector[50] +matrix[51][304] * vector[51] +matrix[52][304] * vector[52] +matrix[53][304] * vector[53] +matrix[54][304] * vector[54] +matrix[55][304] * vector[55] +matrix[56][304] * vector[56] +matrix[57][304] * vector[57] +matrix[58][304] * vector[58] +matrix[59][304] * vector[59] +matrix[60][304] * vector[60] +matrix[61][304] * vector[61] +matrix[62][304] * vector[62] +matrix[63][304] * vector[63] +matrix[64][304] * vector[64] +matrix[65][304] * vector[65] +matrix[66][304] * vector[66] +matrix[67][304] * vector[67] +matrix[68][304] * vector[68] +matrix[69][304] * vector[69] +matrix[70][304] * vector[70] +matrix[71][304] * vector[71] +matrix[72][304] * vector[72] +matrix[73][304] * vector[73] +matrix[74][304] * vector[74] +matrix[75][304] * vector[75] +matrix[76][304] * vector[76] +matrix[77][304] * vector[77] +matrix[78][304] * vector[78] +matrix[79][304] * vector[79] +matrix[80][304] * vector[80] +matrix[81][304] * vector[81] +matrix[82][304] * vector[82] +matrix[83][304] * vector[83] +matrix[84][304] * vector[84] +matrix[85][304] * vector[85] +matrix[86][304] * vector[86] +matrix[87][304] * vector[87] +matrix[88][304] * vector[88] +matrix[89][304] * vector[89] +matrix[90][304] * vector[90] +matrix[91][304] * vector[91] +matrix[92][304] * vector[92] +matrix[93][304] * vector[93] +matrix[94][304] * vector[94] +matrix[95][304] * vector[95] +matrix[96][304] * vector[96] +matrix[97][304] * vector[97] +matrix[98][304] * vector[98] +matrix[99][304] * vector[99] +b[304];
assign result[305] = matrix[0][305] * vector[0] +matrix[1][305] * vector[1] +matrix[2][305] * vector[2] +matrix[3][305] * vector[3] +matrix[4][305] * vector[4] +matrix[5][305] * vector[5] +matrix[6][305] * vector[6] +matrix[7][305] * vector[7] +matrix[8][305] * vector[8] +matrix[9][305] * vector[9] +matrix[10][305] * vector[10] +matrix[11][305] * vector[11] +matrix[12][305] * vector[12] +matrix[13][305] * vector[13] +matrix[14][305] * vector[14] +matrix[15][305] * vector[15] +matrix[16][305] * vector[16] +matrix[17][305] * vector[17] +matrix[18][305] * vector[18] +matrix[19][305] * vector[19] +matrix[20][305] * vector[20] +matrix[21][305] * vector[21] +matrix[22][305] * vector[22] +matrix[23][305] * vector[23] +matrix[24][305] * vector[24] +matrix[25][305] * vector[25] +matrix[26][305] * vector[26] +matrix[27][305] * vector[27] +matrix[28][305] * vector[28] +matrix[29][305] * vector[29] +matrix[30][305] * vector[30] +matrix[31][305] * vector[31] +matrix[32][305] * vector[32] +matrix[33][305] * vector[33] +matrix[34][305] * vector[34] +matrix[35][305] * vector[35] +matrix[36][305] * vector[36] +matrix[37][305] * vector[37] +matrix[38][305] * vector[38] +matrix[39][305] * vector[39] +matrix[40][305] * vector[40] +matrix[41][305] * vector[41] +matrix[42][305] * vector[42] +matrix[43][305] * vector[43] +matrix[44][305] * vector[44] +matrix[45][305] * vector[45] +matrix[46][305] * vector[46] +matrix[47][305] * vector[47] +matrix[48][305] * vector[48] +matrix[49][305] * vector[49] +matrix[50][305] * vector[50] +matrix[51][305] * vector[51] +matrix[52][305] * vector[52] +matrix[53][305] * vector[53] +matrix[54][305] * vector[54] +matrix[55][305] * vector[55] +matrix[56][305] * vector[56] +matrix[57][305] * vector[57] +matrix[58][305] * vector[58] +matrix[59][305] * vector[59] +matrix[60][305] * vector[60] +matrix[61][305] * vector[61] +matrix[62][305] * vector[62] +matrix[63][305] * vector[63] +matrix[64][305] * vector[64] +matrix[65][305] * vector[65] +matrix[66][305] * vector[66] +matrix[67][305] * vector[67] +matrix[68][305] * vector[68] +matrix[69][305] * vector[69] +matrix[70][305] * vector[70] +matrix[71][305] * vector[71] +matrix[72][305] * vector[72] +matrix[73][305] * vector[73] +matrix[74][305] * vector[74] +matrix[75][305] * vector[75] +matrix[76][305] * vector[76] +matrix[77][305] * vector[77] +matrix[78][305] * vector[78] +matrix[79][305] * vector[79] +matrix[80][305] * vector[80] +matrix[81][305] * vector[81] +matrix[82][305] * vector[82] +matrix[83][305] * vector[83] +matrix[84][305] * vector[84] +matrix[85][305] * vector[85] +matrix[86][305] * vector[86] +matrix[87][305] * vector[87] +matrix[88][305] * vector[88] +matrix[89][305] * vector[89] +matrix[90][305] * vector[90] +matrix[91][305] * vector[91] +matrix[92][305] * vector[92] +matrix[93][305] * vector[93] +matrix[94][305] * vector[94] +matrix[95][305] * vector[95] +matrix[96][305] * vector[96] +matrix[97][305] * vector[97] +matrix[98][305] * vector[98] +matrix[99][305] * vector[99] +b[305];
assign result[306] = matrix[0][306] * vector[0] +matrix[1][306] * vector[1] +matrix[2][306] * vector[2] +matrix[3][306] * vector[3] +matrix[4][306] * vector[4] +matrix[5][306] * vector[5] +matrix[6][306] * vector[6] +matrix[7][306] * vector[7] +matrix[8][306] * vector[8] +matrix[9][306] * vector[9] +matrix[10][306] * vector[10] +matrix[11][306] * vector[11] +matrix[12][306] * vector[12] +matrix[13][306] * vector[13] +matrix[14][306] * vector[14] +matrix[15][306] * vector[15] +matrix[16][306] * vector[16] +matrix[17][306] * vector[17] +matrix[18][306] * vector[18] +matrix[19][306] * vector[19] +matrix[20][306] * vector[20] +matrix[21][306] * vector[21] +matrix[22][306] * vector[22] +matrix[23][306] * vector[23] +matrix[24][306] * vector[24] +matrix[25][306] * vector[25] +matrix[26][306] * vector[26] +matrix[27][306] * vector[27] +matrix[28][306] * vector[28] +matrix[29][306] * vector[29] +matrix[30][306] * vector[30] +matrix[31][306] * vector[31] +matrix[32][306] * vector[32] +matrix[33][306] * vector[33] +matrix[34][306] * vector[34] +matrix[35][306] * vector[35] +matrix[36][306] * vector[36] +matrix[37][306] * vector[37] +matrix[38][306] * vector[38] +matrix[39][306] * vector[39] +matrix[40][306] * vector[40] +matrix[41][306] * vector[41] +matrix[42][306] * vector[42] +matrix[43][306] * vector[43] +matrix[44][306] * vector[44] +matrix[45][306] * vector[45] +matrix[46][306] * vector[46] +matrix[47][306] * vector[47] +matrix[48][306] * vector[48] +matrix[49][306] * vector[49] +matrix[50][306] * vector[50] +matrix[51][306] * vector[51] +matrix[52][306] * vector[52] +matrix[53][306] * vector[53] +matrix[54][306] * vector[54] +matrix[55][306] * vector[55] +matrix[56][306] * vector[56] +matrix[57][306] * vector[57] +matrix[58][306] * vector[58] +matrix[59][306] * vector[59] +matrix[60][306] * vector[60] +matrix[61][306] * vector[61] +matrix[62][306] * vector[62] +matrix[63][306] * vector[63] +matrix[64][306] * vector[64] +matrix[65][306] * vector[65] +matrix[66][306] * vector[66] +matrix[67][306] * vector[67] +matrix[68][306] * vector[68] +matrix[69][306] * vector[69] +matrix[70][306] * vector[70] +matrix[71][306] * vector[71] +matrix[72][306] * vector[72] +matrix[73][306] * vector[73] +matrix[74][306] * vector[74] +matrix[75][306] * vector[75] +matrix[76][306] * vector[76] +matrix[77][306] * vector[77] +matrix[78][306] * vector[78] +matrix[79][306] * vector[79] +matrix[80][306] * vector[80] +matrix[81][306] * vector[81] +matrix[82][306] * vector[82] +matrix[83][306] * vector[83] +matrix[84][306] * vector[84] +matrix[85][306] * vector[85] +matrix[86][306] * vector[86] +matrix[87][306] * vector[87] +matrix[88][306] * vector[88] +matrix[89][306] * vector[89] +matrix[90][306] * vector[90] +matrix[91][306] * vector[91] +matrix[92][306] * vector[92] +matrix[93][306] * vector[93] +matrix[94][306] * vector[94] +matrix[95][306] * vector[95] +matrix[96][306] * vector[96] +matrix[97][306] * vector[97] +matrix[98][306] * vector[98] +matrix[99][306] * vector[99] +b[306];
assign result[307] = matrix[0][307] * vector[0] +matrix[1][307] * vector[1] +matrix[2][307] * vector[2] +matrix[3][307] * vector[3] +matrix[4][307] * vector[4] +matrix[5][307] * vector[5] +matrix[6][307] * vector[6] +matrix[7][307] * vector[7] +matrix[8][307] * vector[8] +matrix[9][307] * vector[9] +matrix[10][307] * vector[10] +matrix[11][307] * vector[11] +matrix[12][307] * vector[12] +matrix[13][307] * vector[13] +matrix[14][307] * vector[14] +matrix[15][307] * vector[15] +matrix[16][307] * vector[16] +matrix[17][307] * vector[17] +matrix[18][307] * vector[18] +matrix[19][307] * vector[19] +matrix[20][307] * vector[20] +matrix[21][307] * vector[21] +matrix[22][307] * vector[22] +matrix[23][307] * vector[23] +matrix[24][307] * vector[24] +matrix[25][307] * vector[25] +matrix[26][307] * vector[26] +matrix[27][307] * vector[27] +matrix[28][307] * vector[28] +matrix[29][307] * vector[29] +matrix[30][307] * vector[30] +matrix[31][307] * vector[31] +matrix[32][307] * vector[32] +matrix[33][307] * vector[33] +matrix[34][307] * vector[34] +matrix[35][307] * vector[35] +matrix[36][307] * vector[36] +matrix[37][307] * vector[37] +matrix[38][307] * vector[38] +matrix[39][307] * vector[39] +matrix[40][307] * vector[40] +matrix[41][307] * vector[41] +matrix[42][307] * vector[42] +matrix[43][307] * vector[43] +matrix[44][307] * vector[44] +matrix[45][307] * vector[45] +matrix[46][307] * vector[46] +matrix[47][307] * vector[47] +matrix[48][307] * vector[48] +matrix[49][307] * vector[49] +matrix[50][307] * vector[50] +matrix[51][307] * vector[51] +matrix[52][307] * vector[52] +matrix[53][307] * vector[53] +matrix[54][307] * vector[54] +matrix[55][307] * vector[55] +matrix[56][307] * vector[56] +matrix[57][307] * vector[57] +matrix[58][307] * vector[58] +matrix[59][307] * vector[59] +matrix[60][307] * vector[60] +matrix[61][307] * vector[61] +matrix[62][307] * vector[62] +matrix[63][307] * vector[63] +matrix[64][307] * vector[64] +matrix[65][307] * vector[65] +matrix[66][307] * vector[66] +matrix[67][307] * vector[67] +matrix[68][307] * vector[68] +matrix[69][307] * vector[69] +matrix[70][307] * vector[70] +matrix[71][307] * vector[71] +matrix[72][307] * vector[72] +matrix[73][307] * vector[73] +matrix[74][307] * vector[74] +matrix[75][307] * vector[75] +matrix[76][307] * vector[76] +matrix[77][307] * vector[77] +matrix[78][307] * vector[78] +matrix[79][307] * vector[79] +matrix[80][307] * vector[80] +matrix[81][307] * vector[81] +matrix[82][307] * vector[82] +matrix[83][307] * vector[83] +matrix[84][307] * vector[84] +matrix[85][307] * vector[85] +matrix[86][307] * vector[86] +matrix[87][307] * vector[87] +matrix[88][307] * vector[88] +matrix[89][307] * vector[89] +matrix[90][307] * vector[90] +matrix[91][307] * vector[91] +matrix[92][307] * vector[92] +matrix[93][307] * vector[93] +matrix[94][307] * vector[94] +matrix[95][307] * vector[95] +matrix[96][307] * vector[96] +matrix[97][307] * vector[97] +matrix[98][307] * vector[98] +matrix[99][307] * vector[99] +b[307];
assign result[308] = matrix[0][308] * vector[0] +matrix[1][308] * vector[1] +matrix[2][308] * vector[2] +matrix[3][308] * vector[3] +matrix[4][308] * vector[4] +matrix[5][308] * vector[5] +matrix[6][308] * vector[6] +matrix[7][308] * vector[7] +matrix[8][308] * vector[8] +matrix[9][308] * vector[9] +matrix[10][308] * vector[10] +matrix[11][308] * vector[11] +matrix[12][308] * vector[12] +matrix[13][308] * vector[13] +matrix[14][308] * vector[14] +matrix[15][308] * vector[15] +matrix[16][308] * vector[16] +matrix[17][308] * vector[17] +matrix[18][308] * vector[18] +matrix[19][308] * vector[19] +matrix[20][308] * vector[20] +matrix[21][308] * vector[21] +matrix[22][308] * vector[22] +matrix[23][308] * vector[23] +matrix[24][308] * vector[24] +matrix[25][308] * vector[25] +matrix[26][308] * vector[26] +matrix[27][308] * vector[27] +matrix[28][308] * vector[28] +matrix[29][308] * vector[29] +matrix[30][308] * vector[30] +matrix[31][308] * vector[31] +matrix[32][308] * vector[32] +matrix[33][308] * vector[33] +matrix[34][308] * vector[34] +matrix[35][308] * vector[35] +matrix[36][308] * vector[36] +matrix[37][308] * vector[37] +matrix[38][308] * vector[38] +matrix[39][308] * vector[39] +matrix[40][308] * vector[40] +matrix[41][308] * vector[41] +matrix[42][308] * vector[42] +matrix[43][308] * vector[43] +matrix[44][308] * vector[44] +matrix[45][308] * vector[45] +matrix[46][308] * vector[46] +matrix[47][308] * vector[47] +matrix[48][308] * vector[48] +matrix[49][308] * vector[49] +matrix[50][308] * vector[50] +matrix[51][308] * vector[51] +matrix[52][308] * vector[52] +matrix[53][308] * vector[53] +matrix[54][308] * vector[54] +matrix[55][308] * vector[55] +matrix[56][308] * vector[56] +matrix[57][308] * vector[57] +matrix[58][308] * vector[58] +matrix[59][308] * vector[59] +matrix[60][308] * vector[60] +matrix[61][308] * vector[61] +matrix[62][308] * vector[62] +matrix[63][308] * vector[63] +matrix[64][308] * vector[64] +matrix[65][308] * vector[65] +matrix[66][308] * vector[66] +matrix[67][308] * vector[67] +matrix[68][308] * vector[68] +matrix[69][308] * vector[69] +matrix[70][308] * vector[70] +matrix[71][308] * vector[71] +matrix[72][308] * vector[72] +matrix[73][308] * vector[73] +matrix[74][308] * vector[74] +matrix[75][308] * vector[75] +matrix[76][308] * vector[76] +matrix[77][308] * vector[77] +matrix[78][308] * vector[78] +matrix[79][308] * vector[79] +matrix[80][308] * vector[80] +matrix[81][308] * vector[81] +matrix[82][308] * vector[82] +matrix[83][308] * vector[83] +matrix[84][308] * vector[84] +matrix[85][308] * vector[85] +matrix[86][308] * vector[86] +matrix[87][308] * vector[87] +matrix[88][308] * vector[88] +matrix[89][308] * vector[89] +matrix[90][308] * vector[90] +matrix[91][308] * vector[91] +matrix[92][308] * vector[92] +matrix[93][308] * vector[93] +matrix[94][308] * vector[94] +matrix[95][308] * vector[95] +matrix[96][308] * vector[96] +matrix[97][308] * vector[97] +matrix[98][308] * vector[98] +matrix[99][308] * vector[99] +b[308];
assign result[309] = matrix[0][309] * vector[0] +matrix[1][309] * vector[1] +matrix[2][309] * vector[2] +matrix[3][309] * vector[3] +matrix[4][309] * vector[4] +matrix[5][309] * vector[5] +matrix[6][309] * vector[6] +matrix[7][309] * vector[7] +matrix[8][309] * vector[8] +matrix[9][309] * vector[9] +matrix[10][309] * vector[10] +matrix[11][309] * vector[11] +matrix[12][309] * vector[12] +matrix[13][309] * vector[13] +matrix[14][309] * vector[14] +matrix[15][309] * vector[15] +matrix[16][309] * vector[16] +matrix[17][309] * vector[17] +matrix[18][309] * vector[18] +matrix[19][309] * vector[19] +matrix[20][309] * vector[20] +matrix[21][309] * vector[21] +matrix[22][309] * vector[22] +matrix[23][309] * vector[23] +matrix[24][309] * vector[24] +matrix[25][309] * vector[25] +matrix[26][309] * vector[26] +matrix[27][309] * vector[27] +matrix[28][309] * vector[28] +matrix[29][309] * vector[29] +matrix[30][309] * vector[30] +matrix[31][309] * vector[31] +matrix[32][309] * vector[32] +matrix[33][309] * vector[33] +matrix[34][309] * vector[34] +matrix[35][309] * vector[35] +matrix[36][309] * vector[36] +matrix[37][309] * vector[37] +matrix[38][309] * vector[38] +matrix[39][309] * vector[39] +matrix[40][309] * vector[40] +matrix[41][309] * vector[41] +matrix[42][309] * vector[42] +matrix[43][309] * vector[43] +matrix[44][309] * vector[44] +matrix[45][309] * vector[45] +matrix[46][309] * vector[46] +matrix[47][309] * vector[47] +matrix[48][309] * vector[48] +matrix[49][309] * vector[49] +matrix[50][309] * vector[50] +matrix[51][309] * vector[51] +matrix[52][309] * vector[52] +matrix[53][309] * vector[53] +matrix[54][309] * vector[54] +matrix[55][309] * vector[55] +matrix[56][309] * vector[56] +matrix[57][309] * vector[57] +matrix[58][309] * vector[58] +matrix[59][309] * vector[59] +matrix[60][309] * vector[60] +matrix[61][309] * vector[61] +matrix[62][309] * vector[62] +matrix[63][309] * vector[63] +matrix[64][309] * vector[64] +matrix[65][309] * vector[65] +matrix[66][309] * vector[66] +matrix[67][309] * vector[67] +matrix[68][309] * vector[68] +matrix[69][309] * vector[69] +matrix[70][309] * vector[70] +matrix[71][309] * vector[71] +matrix[72][309] * vector[72] +matrix[73][309] * vector[73] +matrix[74][309] * vector[74] +matrix[75][309] * vector[75] +matrix[76][309] * vector[76] +matrix[77][309] * vector[77] +matrix[78][309] * vector[78] +matrix[79][309] * vector[79] +matrix[80][309] * vector[80] +matrix[81][309] * vector[81] +matrix[82][309] * vector[82] +matrix[83][309] * vector[83] +matrix[84][309] * vector[84] +matrix[85][309] * vector[85] +matrix[86][309] * vector[86] +matrix[87][309] * vector[87] +matrix[88][309] * vector[88] +matrix[89][309] * vector[89] +matrix[90][309] * vector[90] +matrix[91][309] * vector[91] +matrix[92][309] * vector[92] +matrix[93][309] * vector[93] +matrix[94][309] * vector[94] +matrix[95][309] * vector[95] +matrix[96][309] * vector[96] +matrix[97][309] * vector[97] +matrix[98][309] * vector[98] +matrix[99][309] * vector[99] +b[309];
assign result[310] = matrix[0][310] * vector[0] +matrix[1][310] * vector[1] +matrix[2][310] * vector[2] +matrix[3][310] * vector[3] +matrix[4][310] * vector[4] +matrix[5][310] * vector[5] +matrix[6][310] * vector[6] +matrix[7][310] * vector[7] +matrix[8][310] * vector[8] +matrix[9][310] * vector[9] +matrix[10][310] * vector[10] +matrix[11][310] * vector[11] +matrix[12][310] * vector[12] +matrix[13][310] * vector[13] +matrix[14][310] * vector[14] +matrix[15][310] * vector[15] +matrix[16][310] * vector[16] +matrix[17][310] * vector[17] +matrix[18][310] * vector[18] +matrix[19][310] * vector[19] +matrix[20][310] * vector[20] +matrix[21][310] * vector[21] +matrix[22][310] * vector[22] +matrix[23][310] * vector[23] +matrix[24][310] * vector[24] +matrix[25][310] * vector[25] +matrix[26][310] * vector[26] +matrix[27][310] * vector[27] +matrix[28][310] * vector[28] +matrix[29][310] * vector[29] +matrix[30][310] * vector[30] +matrix[31][310] * vector[31] +matrix[32][310] * vector[32] +matrix[33][310] * vector[33] +matrix[34][310] * vector[34] +matrix[35][310] * vector[35] +matrix[36][310] * vector[36] +matrix[37][310] * vector[37] +matrix[38][310] * vector[38] +matrix[39][310] * vector[39] +matrix[40][310] * vector[40] +matrix[41][310] * vector[41] +matrix[42][310] * vector[42] +matrix[43][310] * vector[43] +matrix[44][310] * vector[44] +matrix[45][310] * vector[45] +matrix[46][310] * vector[46] +matrix[47][310] * vector[47] +matrix[48][310] * vector[48] +matrix[49][310] * vector[49] +matrix[50][310] * vector[50] +matrix[51][310] * vector[51] +matrix[52][310] * vector[52] +matrix[53][310] * vector[53] +matrix[54][310] * vector[54] +matrix[55][310] * vector[55] +matrix[56][310] * vector[56] +matrix[57][310] * vector[57] +matrix[58][310] * vector[58] +matrix[59][310] * vector[59] +matrix[60][310] * vector[60] +matrix[61][310] * vector[61] +matrix[62][310] * vector[62] +matrix[63][310] * vector[63] +matrix[64][310] * vector[64] +matrix[65][310] * vector[65] +matrix[66][310] * vector[66] +matrix[67][310] * vector[67] +matrix[68][310] * vector[68] +matrix[69][310] * vector[69] +matrix[70][310] * vector[70] +matrix[71][310] * vector[71] +matrix[72][310] * vector[72] +matrix[73][310] * vector[73] +matrix[74][310] * vector[74] +matrix[75][310] * vector[75] +matrix[76][310] * vector[76] +matrix[77][310] * vector[77] +matrix[78][310] * vector[78] +matrix[79][310] * vector[79] +matrix[80][310] * vector[80] +matrix[81][310] * vector[81] +matrix[82][310] * vector[82] +matrix[83][310] * vector[83] +matrix[84][310] * vector[84] +matrix[85][310] * vector[85] +matrix[86][310] * vector[86] +matrix[87][310] * vector[87] +matrix[88][310] * vector[88] +matrix[89][310] * vector[89] +matrix[90][310] * vector[90] +matrix[91][310] * vector[91] +matrix[92][310] * vector[92] +matrix[93][310] * vector[93] +matrix[94][310] * vector[94] +matrix[95][310] * vector[95] +matrix[96][310] * vector[96] +matrix[97][310] * vector[97] +matrix[98][310] * vector[98] +matrix[99][310] * vector[99] +b[310];
assign result[311] = matrix[0][311] * vector[0] +matrix[1][311] * vector[1] +matrix[2][311] * vector[2] +matrix[3][311] * vector[3] +matrix[4][311] * vector[4] +matrix[5][311] * vector[5] +matrix[6][311] * vector[6] +matrix[7][311] * vector[7] +matrix[8][311] * vector[8] +matrix[9][311] * vector[9] +matrix[10][311] * vector[10] +matrix[11][311] * vector[11] +matrix[12][311] * vector[12] +matrix[13][311] * vector[13] +matrix[14][311] * vector[14] +matrix[15][311] * vector[15] +matrix[16][311] * vector[16] +matrix[17][311] * vector[17] +matrix[18][311] * vector[18] +matrix[19][311] * vector[19] +matrix[20][311] * vector[20] +matrix[21][311] * vector[21] +matrix[22][311] * vector[22] +matrix[23][311] * vector[23] +matrix[24][311] * vector[24] +matrix[25][311] * vector[25] +matrix[26][311] * vector[26] +matrix[27][311] * vector[27] +matrix[28][311] * vector[28] +matrix[29][311] * vector[29] +matrix[30][311] * vector[30] +matrix[31][311] * vector[31] +matrix[32][311] * vector[32] +matrix[33][311] * vector[33] +matrix[34][311] * vector[34] +matrix[35][311] * vector[35] +matrix[36][311] * vector[36] +matrix[37][311] * vector[37] +matrix[38][311] * vector[38] +matrix[39][311] * vector[39] +matrix[40][311] * vector[40] +matrix[41][311] * vector[41] +matrix[42][311] * vector[42] +matrix[43][311] * vector[43] +matrix[44][311] * vector[44] +matrix[45][311] * vector[45] +matrix[46][311] * vector[46] +matrix[47][311] * vector[47] +matrix[48][311] * vector[48] +matrix[49][311] * vector[49] +matrix[50][311] * vector[50] +matrix[51][311] * vector[51] +matrix[52][311] * vector[52] +matrix[53][311] * vector[53] +matrix[54][311] * vector[54] +matrix[55][311] * vector[55] +matrix[56][311] * vector[56] +matrix[57][311] * vector[57] +matrix[58][311] * vector[58] +matrix[59][311] * vector[59] +matrix[60][311] * vector[60] +matrix[61][311] * vector[61] +matrix[62][311] * vector[62] +matrix[63][311] * vector[63] +matrix[64][311] * vector[64] +matrix[65][311] * vector[65] +matrix[66][311] * vector[66] +matrix[67][311] * vector[67] +matrix[68][311] * vector[68] +matrix[69][311] * vector[69] +matrix[70][311] * vector[70] +matrix[71][311] * vector[71] +matrix[72][311] * vector[72] +matrix[73][311] * vector[73] +matrix[74][311] * vector[74] +matrix[75][311] * vector[75] +matrix[76][311] * vector[76] +matrix[77][311] * vector[77] +matrix[78][311] * vector[78] +matrix[79][311] * vector[79] +matrix[80][311] * vector[80] +matrix[81][311] * vector[81] +matrix[82][311] * vector[82] +matrix[83][311] * vector[83] +matrix[84][311] * vector[84] +matrix[85][311] * vector[85] +matrix[86][311] * vector[86] +matrix[87][311] * vector[87] +matrix[88][311] * vector[88] +matrix[89][311] * vector[89] +matrix[90][311] * vector[90] +matrix[91][311] * vector[91] +matrix[92][311] * vector[92] +matrix[93][311] * vector[93] +matrix[94][311] * vector[94] +matrix[95][311] * vector[95] +matrix[96][311] * vector[96] +matrix[97][311] * vector[97] +matrix[98][311] * vector[98] +matrix[99][311] * vector[99] +b[311];
assign result[312] = matrix[0][312] * vector[0] +matrix[1][312] * vector[1] +matrix[2][312] * vector[2] +matrix[3][312] * vector[3] +matrix[4][312] * vector[4] +matrix[5][312] * vector[5] +matrix[6][312] * vector[6] +matrix[7][312] * vector[7] +matrix[8][312] * vector[8] +matrix[9][312] * vector[9] +matrix[10][312] * vector[10] +matrix[11][312] * vector[11] +matrix[12][312] * vector[12] +matrix[13][312] * vector[13] +matrix[14][312] * vector[14] +matrix[15][312] * vector[15] +matrix[16][312] * vector[16] +matrix[17][312] * vector[17] +matrix[18][312] * vector[18] +matrix[19][312] * vector[19] +matrix[20][312] * vector[20] +matrix[21][312] * vector[21] +matrix[22][312] * vector[22] +matrix[23][312] * vector[23] +matrix[24][312] * vector[24] +matrix[25][312] * vector[25] +matrix[26][312] * vector[26] +matrix[27][312] * vector[27] +matrix[28][312] * vector[28] +matrix[29][312] * vector[29] +matrix[30][312] * vector[30] +matrix[31][312] * vector[31] +matrix[32][312] * vector[32] +matrix[33][312] * vector[33] +matrix[34][312] * vector[34] +matrix[35][312] * vector[35] +matrix[36][312] * vector[36] +matrix[37][312] * vector[37] +matrix[38][312] * vector[38] +matrix[39][312] * vector[39] +matrix[40][312] * vector[40] +matrix[41][312] * vector[41] +matrix[42][312] * vector[42] +matrix[43][312] * vector[43] +matrix[44][312] * vector[44] +matrix[45][312] * vector[45] +matrix[46][312] * vector[46] +matrix[47][312] * vector[47] +matrix[48][312] * vector[48] +matrix[49][312] * vector[49] +matrix[50][312] * vector[50] +matrix[51][312] * vector[51] +matrix[52][312] * vector[52] +matrix[53][312] * vector[53] +matrix[54][312] * vector[54] +matrix[55][312] * vector[55] +matrix[56][312] * vector[56] +matrix[57][312] * vector[57] +matrix[58][312] * vector[58] +matrix[59][312] * vector[59] +matrix[60][312] * vector[60] +matrix[61][312] * vector[61] +matrix[62][312] * vector[62] +matrix[63][312] * vector[63] +matrix[64][312] * vector[64] +matrix[65][312] * vector[65] +matrix[66][312] * vector[66] +matrix[67][312] * vector[67] +matrix[68][312] * vector[68] +matrix[69][312] * vector[69] +matrix[70][312] * vector[70] +matrix[71][312] * vector[71] +matrix[72][312] * vector[72] +matrix[73][312] * vector[73] +matrix[74][312] * vector[74] +matrix[75][312] * vector[75] +matrix[76][312] * vector[76] +matrix[77][312] * vector[77] +matrix[78][312] * vector[78] +matrix[79][312] * vector[79] +matrix[80][312] * vector[80] +matrix[81][312] * vector[81] +matrix[82][312] * vector[82] +matrix[83][312] * vector[83] +matrix[84][312] * vector[84] +matrix[85][312] * vector[85] +matrix[86][312] * vector[86] +matrix[87][312] * vector[87] +matrix[88][312] * vector[88] +matrix[89][312] * vector[89] +matrix[90][312] * vector[90] +matrix[91][312] * vector[91] +matrix[92][312] * vector[92] +matrix[93][312] * vector[93] +matrix[94][312] * vector[94] +matrix[95][312] * vector[95] +matrix[96][312] * vector[96] +matrix[97][312] * vector[97] +matrix[98][312] * vector[98] +matrix[99][312] * vector[99] +b[312];
assign result[313] = matrix[0][313] * vector[0] +matrix[1][313] * vector[1] +matrix[2][313] * vector[2] +matrix[3][313] * vector[3] +matrix[4][313] * vector[4] +matrix[5][313] * vector[5] +matrix[6][313] * vector[6] +matrix[7][313] * vector[7] +matrix[8][313] * vector[8] +matrix[9][313] * vector[9] +matrix[10][313] * vector[10] +matrix[11][313] * vector[11] +matrix[12][313] * vector[12] +matrix[13][313] * vector[13] +matrix[14][313] * vector[14] +matrix[15][313] * vector[15] +matrix[16][313] * vector[16] +matrix[17][313] * vector[17] +matrix[18][313] * vector[18] +matrix[19][313] * vector[19] +matrix[20][313] * vector[20] +matrix[21][313] * vector[21] +matrix[22][313] * vector[22] +matrix[23][313] * vector[23] +matrix[24][313] * vector[24] +matrix[25][313] * vector[25] +matrix[26][313] * vector[26] +matrix[27][313] * vector[27] +matrix[28][313] * vector[28] +matrix[29][313] * vector[29] +matrix[30][313] * vector[30] +matrix[31][313] * vector[31] +matrix[32][313] * vector[32] +matrix[33][313] * vector[33] +matrix[34][313] * vector[34] +matrix[35][313] * vector[35] +matrix[36][313] * vector[36] +matrix[37][313] * vector[37] +matrix[38][313] * vector[38] +matrix[39][313] * vector[39] +matrix[40][313] * vector[40] +matrix[41][313] * vector[41] +matrix[42][313] * vector[42] +matrix[43][313] * vector[43] +matrix[44][313] * vector[44] +matrix[45][313] * vector[45] +matrix[46][313] * vector[46] +matrix[47][313] * vector[47] +matrix[48][313] * vector[48] +matrix[49][313] * vector[49] +matrix[50][313] * vector[50] +matrix[51][313] * vector[51] +matrix[52][313] * vector[52] +matrix[53][313] * vector[53] +matrix[54][313] * vector[54] +matrix[55][313] * vector[55] +matrix[56][313] * vector[56] +matrix[57][313] * vector[57] +matrix[58][313] * vector[58] +matrix[59][313] * vector[59] +matrix[60][313] * vector[60] +matrix[61][313] * vector[61] +matrix[62][313] * vector[62] +matrix[63][313] * vector[63] +matrix[64][313] * vector[64] +matrix[65][313] * vector[65] +matrix[66][313] * vector[66] +matrix[67][313] * vector[67] +matrix[68][313] * vector[68] +matrix[69][313] * vector[69] +matrix[70][313] * vector[70] +matrix[71][313] * vector[71] +matrix[72][313] * vector[72] +matrix[73][313] * vector[73] +matrix[74][313] * vector[74] +matrix[75][313] * vector[75] +matrix[76][313] * vector[76] +matrix[77][313] * vector[77] +matrix[78][313] * vector[78] +matrix[79][313] * vector[79] +matrix[80][313] * vector[80] +matrix[81][313] * vector[81] +matrix[82][313] * vector[82] +matrix[83][313] * vector[83] +matrix[84][313] * vector[84] +matrix[85][313] * vector[85] +matrix[86][313] * vector[86] +matrix[87][313] * vector[87] +matrix[88][313] * vector[88] +matrix[89][313] * vector[89] +matrix[90][313] * vector[90] +matrix[91][313] * vector[91] +matrix[92][313] * vector[92] +matrix[93][313] * vector[93] +matrix[94][313] * vector[94] +matrix[95][313] * vector[95] +matrix[96][313] * vector[96] +matrix[97][313] * vector[97] +matrix[98][313] * vector[98] +matrix[99][313] * vector[99] +b[313];
assign result[314] = matrix[0][314] * vector[0] +matrix[1][314] * vector[1] +matrix[2][314] * vector[2] +matrix[3][314] * vector[3] +matrix[4][314] * vector[4] +matrix[5][314] * vector[5] +matrix[6][314] * vector[6] +matrix[7][314] * vector[7] +matrix[8][314] * vector[8] +matrix[9][314] * vector[9] +matrix[10][314] * vector[10] +matrix[11][314] * vector[11] +matrix[12][314] * vector[12] +matrix[13][314] * vector[13] +matrix[14][314] * vector[14] +matrix[15][314] * vector[15] +matrix[16][314] * vector[16] +matrix[17][314] * vector[17] +matrix[18][314] * vector[18] +matrix[19][314] * vector[19] +matrix[20][314] * vector[20] +matrix[21][314] * vector[21] +matrix[22][314] * vector[22] +matrix[23][314] * vector[23] +matrix[24][314] * vector[24] +matrix[25][314] * vector[25] +matrix[26][314] * vector[26] +matrix[27][314] * vector[27] +matrix[28][314] * vector[28] +matrix[29][314] * vector[29] +matrix[30][314] * vector[30] +matrix[31][314] * vector[31] +matrix[32][314] * vector[32] +matrix[33][314] * vector[33] +matrix[34][314] * vector[34] +matrix[35][314] * vector[35] +matrix[36][314] * vector[36] +matrix[37][314] * vector[37] +matrix[38][314] * vector[38] +matrix[39][314] * vector[39] +matrix[40][314] * vector[40] +matrix[41][314] * vector[41] +matrix[42][314] * vector[42] +matrix[43][314] * vector[43] +matrix[44][314] * vector[44] +matrix[45][314] * vector[45] +matrix[46][314] * vector[46] +matrix[47][314] * vector[47] +matrix[48][314] * vector[48] +matrix[49][314] * vector[49] +matrix[50][314] * vector[50] +matrix[51][314] * vector[51] +matrix[52][314] * vector[52] +matrix[53][314] * vector[53] +matrix[54][314] * vector[54] +matrix[55][314] * vector[55] +matrix[56][314] * vector[56] +matrix[57][314] * vector[57] +matrix[58][314] * vector[58] +matrix[59][314] * vector[59] +matrix[60][314] * vector[60] +matrix[61][314] * vector[61] +matrix[62][314] * vector[62] +matrix[63][314] * vector[63] +matrix[64][314] * vector[64] +matrix[65][314] * vector[65] +matrix[66][314] * vector[66] +matrix[67][314] * vector[67] +matrix[68][314] * vector[68] +matrix[69][314] * vector[69] +matrix[70][314] * vector[70] +matrix[71][314] * vector[71] +matrix[72][314] * vector[72] +matrix[73][314] * vector[73] +matrix[74][314] * vector[74] +matrix[75][314] * vector[75] +matrix[76][314] * vector[76] +matrix[77][314] * vector[77] +matrix[78][314] * vector[78] +matrix[79][314] * vector[79] +matrix[80][314] * vector[80] +matrix[81][314] * vector[81] +matrix[82][314] * vector[82] +matrix[83][314] * vector[83] +matrix[84][314] * vector[84] +matrix[85][314] * vector[85] +matrix[86][314] * vector[86] +matrix[87][314] * vector[87] +matrix[88][314] * vector[88] +matrix[89][314] * vector[89] +matrix[90][314] * vector[90] +matrix[91][314] * vector[91] +matrix[92][314] * vector[92] +matrix[93][314] * vector[93] +matrix[94][314] * vector[94] +matrix[95][314] * vector[95] +matrix[96][314] * vector[96] +matrix[97][314] * vector[97] +matrix[98][314] * vector[98] +matrix[99][314] * vector[99] +b[314];
assign result[315] = matrix[0][315] * vector[0] +matrix[1][315] * vector[1] +matrix[2][315] * vector[2] +matrix[3][315] * vector[3] +matrix[4][315] * vector[4] +matrix[5][315] * vector[5] +matrix[6][315] * vector[6] +matrix[7][315] * vector[7] +matrix[8][315] * vector[8] +matrix[9][315] * vector[9] +matrix[10][315] * vector[10] +matrix[11][315] * vector[11] +matrix[12][315] * vector[12] +matrix[13][315] * vector[13] +matrix[14][315] * vector[14] +matrix[15][315] * vector[15] +matrix[16][315] * vector[16] +matrix[17][315] * vector[17] +matrix[18][315] * vector[18] +matrix[19][315] * vector[19] +matrix[20][315] * vector[20] +matrix[21][315] * vector[21] +matrix[22][315] * vector[22] +matrix[23][315] * vector[23] +matrix[24][315] * vector[24] +matrix[25][315] * vector[25] +matrix[26][315] * vector[26] +matrix[27][315] * vector[27] +matrix[28][315] * vector[28] +matrix[29][315] * vector[29] +matrix[30][315] * vector[30] +matrix[31][315] * vector[31] +matrix[32][315] * vector[32] +matrix[33][315] * vector[33] +matrix[34][315] * vector[34] +matrix[35][315] * vector[35] +matrix[36][315] * vector[36] +matrix[37][315] * vector[37] +matrix[38][315] * vector[38] +matrix[39][315] * vector[39] +matrix[40][315] * vector[40] +matrix[41][315] * vector[41] +matrix[42][315] * vector[42] +matrix[43][315] * vector[43] +matrix[44][315] * vector[44] +matrix[45][315] * vector[45] +matrix[46][315] * vector[46] +matrix[47][315] * vector[47] +matrix[48][315] * vector[48] +matrix[49][315] * vector[49] +matrix[50][315] * vector[50] +matrix[51][315] * vector[51] +matrix[52][315] * vector[52] +matrix[53][315] * vector[53] +matrix[54][315] * vector[54] +matrix[55][315] * vector[55] +matrix[56][315] * vector[56] +matrix[57][315] * vector[57] +matrix[58][315] * vector[58] +matrix[59][315] * vector[59] +matrix[60][315] * vector[60] +matrix[61][315] * vector[61] +matrix[62][315] * vector[62] +matrix[63][315] * vector[63] +matrix[64][315] * vector[64] +matrix[65][315] * vector[65] +matrix[66][315] * vector[66] +matrix[67][315] * vector[67] +matrix[68][315] * vector[68] +matrix[69][315] * vector[69] +matrix[70][315] * vector[70] +matrix[71][315] * vector[71] +matrix[72][315] * vector[72] +matrix[73][315] * vector[73] +matrix[74][315] * vector[74] +matrix[75][315] * vector[75] +matrix[76][315] * vector[76] +matrix[77][315] * vector[77] +matrix[78][315] * vector[78] +matrix[79][315] * vector[79] +matrix[80][315] * vector[80] +matrix[81][315] * vector[81] +matrix[82][315] * vector[82] +matrix[83][315] * vector[83] +matrix[84][315] * vector[84] +matrix[85][315] * vector[85] +matrix[86][315] * vector[86] +matrix[87][315] * vector[87] +matrix[88][315] * vector[88] +matrix[89][315] * vector[89] +matrix[90][315] * vector[90] +matrix[91][315] * vector[91] +matrix[92][315] * vector[92] +matrix[93][315] * vector[93] +matrix[94][315] * vector[94] +matrix[95][315] * vector[95] +matrix[96][315] * vector[96] +matrix[97][315] * vector[97] +matrix[98][315] * vector[98] +matrix[99][315] * vector[99] +b[315];
assign result[316] = matrix[0][316] * vector[0] +matrix[1][316] * vector[1] +matrix[2][316] * vector[2] +matrix[3][316] * vector[3] +matrix[4][316] * vector[4] +matrix[5][316] * vector[5] +matrix[6][316] * vector[6] +matrix[7][316] * vector[7] +matrix[8][316] * vector[8] +matrix[9][316] * vector[9] +matrix[10][316] * vector[10] +matrix[11][316] * vector[11] +matrix[12][316] * vector[12] +matrix[13][316] * vector[13] +matrix[14][316] * vector[14] +matrix[15][316] * vector[15] +matrix[16][316] * vector[16] +matrix[17][316] * vector[17] +matrix[18][316] * vector[18] +matrix[19][316] * vector[19] +matrix[20][316] * vector[20] +matrix[21][316] * vector[21] +matrix[22][316] * vector[22] +matrix[23][316] * vector[23] +matrix[24][316] * vector[24] +matrix[25][316] * vector[25] +matrix[26][316] * vector[26] +matrix[27][316] * vector[27] +matrix[28][316] * vector[28] +matrix[29][316] * vector[29] +matrix[30][316] * vector[30] +matrix[31][316] * vector[31] +matrix[32][316] * vector[32] +matrix[33][316] * vector[33] +matrix[34][316] * vector[34] +matrix[35][316] * vector[35] +matrix[36][316] * vector[36] +matrix[37][316] * vector[37] +matrix[38][316] * vector[38] +matrix[39][316] * vector[39] +matrix[40][316] * vector[40] +matrix[41][316] * vector[41] +matrix[42][316] * vector[42] +matrix[43][316] * vector[43] +matrix[44][316] * vector[44] +matrix[45][316] * vector[45] +matrix[46][316] * vector[46] +matrix[47][316] * vector[47] +matrix[48][316] * vector[48] +matrix[49][316] * vector[49] +matrix[50][316] * vector[50] +matrix[51][316] * vector[51] +matrix[52][316] * vector[52] +matrix[53][316] * vector[53] +matrix[54][316] * vector[54] +matrix[55][316] * vector[55] +matrix[56][316] * vector[56] +matrix[57][316] * vector[57] +matrix[58][316] * vector[58] +matrix[59][316] * vector[59] +matrix[60][316] * vector[60] +matrix[61][316] * vector[61] +matrix[62][316] * vector[62] +matrix[63][316] * vector[63] +matrix[64][316] * vector[64] +matrix[65][316] * vector[65] +matrix[66][316] * vector[66] +matrix[67][316] * vector[67] +matrix[68][316] * vector[68] +matrix[69][316] * vector[69] +matrix[70][316] * vector[70] +matrix[71][316] * vector[71] +matrix[72][316] * vector[72] +matrix[73][316] * vector[73] +matrix[74][316] * vector[74] +matrix[75][316] * vector[75] +matrix[76][316] * vector[76] +matrix[77][316] * vector[77] +matrix[78][316] * vector[78] +matrix[79][316] * vector[79] +matrix[80][316] * vector[80] +matrix[81][316] * vector[81] +matrix[82][316] * vector[82] +matrix[83][316] * vector[83] +matrix[84][316] * vector[84] +matrix[85][316] * vector[85] +matrix[86][316] * vector[86] +matrix[87][316] * vector[87] +matrix[88][316] * vector[88] +matrix[89][316] * vector[89] +matrix[90][316] * vector[90] +matrix[91][316] * vector[91] +matrix[92][316] * vector[92] +matrix[93][316] * vector[93] +matrix[94][316] * vector[94] +matrix[95][316] * vector[95] +matrix[96][316] * vector[96] +matrix[97][316] * vector[97] +matrix[98][316] * vector[98] +matrix[99][316] * vector[99] +b[316];
assign result[317] = matrix[0][317] * vector[0] +matrix[1][317] * vector[1] +matrix[2][317] * vector[2] +matrix[3][317] * vector[3] +matrix[4][317] * vector[4] +matrix[5][317] * vector[5] +matrix[6][317] * vector[6] +matrix[7][317] * vector[7] +matrix[8][317] * vector[8] +matrix[9][317] * vector[9] +matrix[10][317] * vector[10] +matrix[11][317] * vector[11] +matrix[12][317] * vector[12] +matrix[13][317] * vector[13] +matrix[14][317] * vector[14] +matrix[15][317] * vector[15] +matrix[16][317] * vector[16] +matrix[17][317] * vector[17] +matrix[18][317] * vector[18] +matrix[19][317] * vector[19] +matrix[20][317] * vector[20] +matrix[21][317] * vector[21] +matrix[22][317] * vector[22] +matrix[23][317] * vector[23] +matrix[24][317] * vector[24] +matrix[25][317] * vector[25] +matrix[26][317] * vector[26] +matrix[27][317] * vector[27] +matrix[28][317] * vector[28] +matrix[29][317] * vector[29] +matrix[30][317] * vector[30] +matrix[31][317] * vector[31] +matrix[32][317] * vector[32] +matrix[33][317] * vector[33] +matrix[34][317] * vector[34] +matrix[35][317] * vector[35] +matrix[36][317] * vector[36] +matrix[37][317] * vector[37] +matrix[38][317] * vector[38] +matrix[39][317] * vector[39] +matrix[40][317] * vector[40] +matrix[41][317] * vector[41] +matrix[42][317] * vector[42] +matrix[43][317] * vector[43] +matrix[44][317] * vector[44] +matrix[45][317] * vector[45] +matrix[46][317] * vector[46] +matrix[47][317] * vector[47] +matrix[48][317] * vector[48] +matrix[49][317] * vector[49] +matrix[50][317] * vector[50] +matrix[51][317] * vector[51] +matrix[52][317] * vector[52] +matrix[53][317] * vector[53] +matrix[54][317] * vector[54] +matrix[55][317] * vector[55] +matrix[56][317] * vector[56] +matrix[57][317] * vector[57] +matrix[58][317] * vector[58] +matrix[59][317] * vector[59] +matrix[60][317] * vector[60] +matrix[61][317] * vector[61] +matrix[62][317] * vector[62] +matrix[63][317] * vector[63] +matrix[64][317] * vector[64] +matrix[65][317] * vector[65] +matrix[66][317] * vector[66] +matrix[67][317] * vector[67] +matrix[68][317] * vector[68] +matrix[69][317] * vector[69] +matrix[70][317] * vector[70] +matrix[71][317] * vector[71] +matrix[72][317] * vector[72] +matrix[73][317] * vector[73] +matrix[74][317] * vector[74] +matrix[75][317] * vector[75] +matrix[76][317] * vector[76] +matrix[77][317] * vector[77] +matrix[78][317] * vector[78] +matrix[79][317] * vector[79] +matrix[80][317] * vector[80] +matrix[81][317] * vector[81] +matrix[82][317] * vector[82] +matrix[83][317] * vector[83] +matrix[84][317] * vector[84] +matrix[85][317] * vector[85] +matrix[86][317] * vector[86] +matrix[87][317] * vector[87] +matrix[88][317] * vector[88] +matrix[89][317] * vector[89] +matrix[90][317] * vector[90] +matrix[91][317] * vector[91] +matrix[92][317] * vector[92] +matrix[93][317] * vector[93] +matrix[94][317] * vector[94] +matrix[95][317] * vector[95] +matrix[96][317] * vector[96] +matrix[97][317] * vector[97] +matrix[98][317] * vector[98] +matrix[99][317] * vector[99] +b[317];
assign result[318] = matrix[0][318] * vector[0] +matrix[1][318] * vector[1] +matrix[2][318] * vector[2] +matrix[3][318] * vector[3] +matrix[4][318] * vector[4] +matrix[5][318] * vector[5] +matrix[6][318] * vector[6] +matrix[7][318] * vector[7] +matrix[8][318] * vector[8] +matrix[9][318] * vector[9] +matrix[10][318] * vector[10] +matrix[11][318] * vector[11] +matrix[12][318] * vector[12] +matrix[13][318] * vector[13] +matrix[14][318] * vector[14] +matrix[15][318] * vector[15] +matrix[16][318] * vector[16] +matrix[17][318] * vector[17] +matrix[18][318] * vector[18] +matrix[19][318] * vector[19] +matrix[20][318] * vector[20] +matrix[21][318] * vector[21] +matrix[22][318] * vector[22] +matrix[23][318] * vector[23] +matrix[24][318] * vector[24] +matrix[25][318] * vector[25] +matrix[26][318] * vector[26] +matrix[27][318] * vector[27] +matrix[28][318] * vector[28] +matrix[29][318] * vector[29] +matrix[30][318] * vector[30] +matrix[31][318] * vector[31] +matrix[32][318] * vector[32] +matrix[33][318] * vector[33] +matrix[34][318] * vector[34] +matrix[35][318] * vector[35] +matrix[36][318] * vector[36] +matrix[37][318] * vector[37] +matrix[38][318] * vector[38] +matrix[39][318] * vector[39] +matrix[40][318] * vector[40] +matrix[41][318] * vector[41] +matrix[42][318] * vector[42] +matrix[43][318] * vector[43] +matrix[44][318] * vector[44] +matrix[45][318] * vector[45] +matrix[46][318] * vector[46] +matrix[47][318] * vector[47] +matrix[48][318] * vector[48] +matrix[49][318] * vector[49] +matrix[50][318] * vector[50] +matrix[51][318] * vector[51] +matrix[52][318] * vector[52] +matrix[53][318] * vector[53] +matrix[54][318] * vector[54] +matrix[55][318] * vector[55] +matrix[56][318] * vector[56] +matrix[57][318] * vector[57] +matrix[58][318] * vector[58] +matrix[59][318] * vector[59] +matrix[60][318] * vector[60] +matrix[61][318] * vector[61] +matrix[62][318] * vector[62] +matrix[63][318] * vector[63] +matrix[64][318] * vector[64] +matrix[65][318] * vector[65] +matrix[66][318] * vector[66] +matrix[67][318] * vector[67] +matrix[68][318] * vector[68] +matrix[69][318] * vector[69] +matrix[70][318] * vector[70] +matrix[71][318] * vector[71] +matrix[72][318] * vector[72] +matrix[73][318] * vector[73] +matrix[74][318] * vector[74] +matrix[75][318] * vector[75] +matrix[76][318] * vector[76] +matrix[77][318] * vector[77] +matrix[78][318] * vector[78] +matrix[79][318] * vector[79] +matrix[80][318] * vector[80] +matrix[81][318] * vector[81] +matrix[82][318] * vector[82] +matrix[83][318] * vector[83] +matrix[84][318] * vector[84] +matrix[85][318] * vector[85] +matrix[86][318] * vector[86] +matrix[87][318] * vector[87] +matrix[88][318] * vector[88] +matrix[89][318] * vector[89] +matrix[90][318] * vector[90] +matrix[91][318] * vector[91] +matrix[92][318] * vector[92] +matrix[93][318] * vector[93] +matrix[94][318] * vector[94] +matrix[95][318] * vector[95] +matrix[96][318] * vector[96] +matrix[97][318] * vector[97] +matrix[98][318] * vector[98] +matrix[99][318] * vector[99] +b[318];
assign result[319] = matrix[0][319] * vector[0] +matrix[1][319] * vector[1] +matrix[2][319] * vector[2] +matrix[3][319] * vector[3] +matrix[4][319] * vector[4] +matrix[5][319] * vector[5] +matrix[6][319] * vector[6] +matrix[7][319] * vector[7] +matrix[8][319] * vector[8] +matrix[9][319] * vector[9] +matrix[10][319] * vector[10] +matrix[11][319] * vector[11] +matrix[12][319] * vector[12] +matrix[13][319] * vector[13] +matrix[14][319] * vector[14] +matrix[15][319] * vector[15] +matrix[16][319] * vector[16] +matrix[17][319] * vector[17] +matrix[18][319] * vector[18] +matrix[19][319] * vector[19] +matrix[20][319] * vector[20] +matrix[21][319] * vector[21] +matrix[22][319] * vector[22] +matrix[23][319] * vector[23] +matrix[24][319] * vector[24] +matrix[25][319] * vector[25] +matrix[26][319] * vector[26] +matrix[27][319] * vector[27] +matrix[28][319] * vector[28] +matrix[29][319] * vector[29] +matrix[30][319] * vector[30] +matrix[31][319] * vector[31] +matrix[32][319] * vector[32] +matrix[33][319] * vector[33] +matrix[34][319] * vector[34] +matrix[35][319] * vector[35] +matrix[36][319] * vector[36] +matrix[37][319] * vector[37] +matrix[38][319] * vector[38] +matrix[39][319] * vector[39] +matrix[40][319] * vector[40] +matrix[41][319] * vector[41] +matrix[42][319] * vector[42] +matrix[43][319] * vector[43] +matrix[44][319] * vector[44] +matrix[45][319] * vector[45] +matrix[46][319] * vector[46] +matrix[47][319] * vector[47] +matrix[48][319] * vector[48] +matrix[49][319] * vector[49] +matrix[50][319] * vector[50] +matrix[51][319] * vector[51] +matrix[52][319] * vector[52] +matrix[53][319] * vector[53] +matrix[54][319] * vector[54] +matrix[55][319] * vector[55] +matrix[56][319] * vector[56] +matrix[57][319] * vector[57] +matrix[58][319] * vector[58] +matrix[59][319] * vector[59] +matrix[60][319] * vector[60] +matrix[61][319] * vector[61] +matrix[62][319] * vector[62] +matrix[63][319] * vector[63] +matrix[64][319] * vector[64] +matrix[65][319] * vector[65] +matrix[66][319] * vector[66] +matrix[67][319] * vector[67] +matrix[68][319] * vector[68] +matrix[69][319] * vector[69] +matrix[70][319] * vector[70] +matrix[71][319] * vector[71] +matrix[72][319] * vector[72] +matrix[73][319] * vector[73] +matrix[74][319] * vector[74] +matrix[75][319] * vector[75] +matrix[76][319] * vector[76] +matrix[77][319] * vector[77] +matrix[78][319] * vector[78] +matrix[79][319] * vector[79] +matrix[80][319] * vector[80] +matrix[81][319] * vector[81] +matrix[82][319] * vector[82] +matrix[83][319] * vector[83] +matrix[84][319] * vector[84] +matrix[85][319] * vector[85] +matrix[86][319] * vector[86] +matrix[87][319] * vector[87] +matrix[88][319] * vector[88] +matrix[89][319] * vector[89] +matrix[90][319] * vector[90] +matrix[91][319] * vector[91] +matrix[92][319] * vector[92] +matrix[93][319] * vector[93] +matrix[94][319] * vector[94] +matrix[95][319] * vector[95] +matrix[96][319] * vector[96] +matrix[97][319] * vector[97] +matrix[98][319] * vector[98] +matrix[99][319] * vector[99] +b[319];
assign result[320] = matrix[0][320] * vector[0] +matrix[1][320] * vector[1] +matrix[2][320] * vector[2] +matrix[3][320] * vector[3] +matrix[4][320] * vector[4] +matrix[5][320] * vector[5] +matrix[6][320] * vector[6] +matrix[7][320] * vector[7] +matrix[8][320] * vector[8] +matrix[9][320] * vector[9] +matrix[10][320] * vector[10] +matrix[11][320] * vector[11] +matrix[12][320] * vector[12] +matrix[13][320] * vector[13] +matrix[14][320] * vector[14] +matrix[15][320] * vector[15] +matrix[16][320] * vector[16] +matrix[17][320] * vector[17] +matrix[18][320] * vector[18] +matrix[19][320] * vector[19] +matrix[20][320] * vector[20] +matrix[21][320] * vector[21] +matrix[22][320] * vector[22] +matrix[23][320] * vector[23] +matrix[24][320] * vector[24] +matrix[25][320] * vector[25] +matrix[26][320] * vector[26] +matrix[27][320] * vector[27] +matrix[28][320] * vector[28] +matrix[29][320] * vector[29] +matrix[30][320] * vector[30] +matrix[31][320] * vector[31] +matrix[32][320] * vector[32] +matrix[33][320] * vector[33] +matrix[34][320] * vector[34] +matrix[35][320] * vector[35] +matrix[36][320] * vector[36] +matrix[37][320] * vector[37] +matrix[38][320] * vector[38] +matrix[39][320] * vector[39] +matrix[40][320] * vector[40] +matrix[41][320] * vector[41] +matrix[42][320] * vector[42] +matrix[43][320] * vector[43] +matrix[44][320] * vector[44] +matrix[45][320] * vector[45] +matrix[46][320] * vector[46] +matrix[47][320] * vector[47] +matrix[48][320] * vector[48] +matrix[49][320] * vector[49] +matrix[50][320] * vector[50] +matrix[51][320] * vector[51] +matrix[52][320] * vector[52] +matrix[53][320] * vector[53] +matrix[54][320] * vector[54] +matrix[55][320] * vector[55] +matrix[56][320] * vector[56] +matrix[57][320] * vector[57] +matrix[58][320] * vector[58] +matrix[59][320] * vector[59] +matrix[60][320] * vector[60] +matrix[61][320] * vector[61] +matrix[62][320] * vector[62] +matrix[63][320] * vector[63] +matrix[64][320] * vector[64] +matrix[65][320] * vector[65] +matrix[66][320] * vector[66] +matrix[67][320] * vector[67] +matrix[68][320] * vector[68] +matrix[69][320] * vector[69] +matrix[70][320] * vector[70] +matrix[71][320] * vector[71] +matrix[72][320] * vector[72] +matrix[73][320] * vector[73] +matrix[74][320] * vector[74] +matrix[75][320] * vector[75] +matrix[76][320] * vector[76] +matrix[77][320] * vector[77] +matrix[78][320] * vector[78] +matrix[79][320] * vector[79] +matrix[80][320] * vector[80] +matrix[81][320] * vector[81] +matrix[82][320] * vector[82] +matrix[83][320] * vector[83] +matrix[84][320] * vector[84] +matrix[85][320] * vector[85] +matrix[86][320] * vector[86] +matrix[87][320] * vector[87] +matrix[88][320] * vector[88] +matrix[89][320] * vector[89] +matrix[90][320] * vector[90] +matrix[91][320] * vector[91] +matrix[92][320] * vector[92] +matrix[93][320] * vector[93] +matrix[94][320] * vector[94] +matrix[95][320] * vector[95] +matrix[96][320] * vector[96] +matrix[97][320] * vector[97] +matrix[98][320] * vector[98] +matrix[99][320] * vector[99] +b[320];
assign result[321] = matrix[0][321] * vector[0] +matrix[1][321] * vector[1] +matrix[2][321] * vector[2] +matrix[3][321] * vector[3] +matrix[4][321] * vector[4] +matrix[5][321] * vector[5] +matrix[6][321] * vector[6] +matrix[7][321] * vector[7] +matrix[8][321] * vector[8] +matrix[9][321] * vector[9] +matrix[10][321] * vector[10] +matrix[11][321] * vector[11] +matrix[12][321] * vector[12] +matrix[13][321] * vector[13] +matrix[14][321] * vector[14] +matrix[15][321] * vector[15] +matrix[16][321] * vector[16] +matrix[17][321] * vector[17] +matrix[18][321] * vector[18] +matrix[19][321] * vector[19] +matrix[20][321] * vector[20] +matrix[21][321] * vector[21] +matrix[22][321] * vector[22] +matrix[23][321] * vector[23] +matrix[24][321] * vector[24] +matrix[25][321] * vector[25] +matrix[26][321] * vector[26] +matrix[27][321] * vector[27] +matrix[28][321] * vector[28] +matrix[29][321] * vector[29] +matrix[30][321] * vector[30] +matrix[31][321] * vector[31] +matrix[32][321] * vector[32] +matrix[33][321] * vector[33] +matrix[34][321] * vector[34] +matrix[35][321] * vector[35] +matrix[36][321] * vector[36] +matrix[37][321] * vector[37] +matrix[38][321] * vector[38] +matrix[39][321] * vector[39] +matrix[40][321] * vector[40] +matrix[41][321] * vector[41] +matrix[42][321] * vector[42] +matrix[43][321] * vector[43] +matrix[44][321] * vector[44] +matrix[45][321] * vector[45] +matrix[46][321] * vector[46] +matrix[47][321] * vector[47] +matrix[48][321] * vector[48] +matrix[49][321] * vector[49] +matrix[50][321] * vector[50] +matrix[51][321] * vector[51] +matrix[52][321] * vector[52] +matrix[53][321] * vector[53] +matrix[54][321] * vector[54] +matrix[55][321] * vector[55] +matrix[56][321] * vector[56] +matrix[57][321] * vector[57] +matrix[58][321] * vector[58] +matrix[59][321] * vector[59] +matrix[60][321] * vector[60] +matrix[61][321] * vector[61] +matrix[62][321] * vector[62] +matrix[63][321] * vector[63] +matrix[64][321] * vector[64] +matrix[65][321] * vector[65] +matrix[66][321] * vector[66] +matrix[67][321] * vector[67] +matrix[68][321] * vector[68] +matrix[69][321] * vector[69] +matrix[70][321] * vector[70] +matrix[71][321] * vector[71] +matrix[72][321] * vector[72] +matrix[73][321] * vector[73] +matrix[74][321] * vector[74] +matrix[75][321] * vector[75] +matrix[76][321] * vector[76] +matrix[77][321] * vector[77] +matrix[78][321] * vector[78] +matrix[79][321] * vector[79] +matrix[80][321] * vector[80] +matrix[81][321] * vector[81] +matrix[82][321] * vector[82] +matrix[83][321] * vector[83] +matrix[84][321] * vector[84] +matrix[85][321] * vector[85] +matrix[86][321] * vector[86] +matrix[87][321] * vector[87] +matrix[88][321] * vector[88] +matrix[89][321] * vector[89] +matrix[90][321] * vector[90] +matrix[91][321] * vector[91] +matrix[92][321] * vector[92] +matrix[93][321] * vector[93] +matrix[94][321] * vector[94] +matrix[95][321] * vector[95] +matrix[96][321] * vector[96] +matrix[97][321] * vector[97] +matrix[98][321] * vector[98] +matrix[99][321] * vector[99] +b[321];
assign result[322] = matrix[0][322] * vector[0] +matrix[1][322] * vector[1] +matrix[2][322] * vector[2] +matrix[3][322] * vector[3] +matrix[4][322] * vector[4] +matrix[5][322] * vector[5] +matrix[6][322] * vector[6] +matrix[7][322] * vector[7] +matrix[8][322] * vector[8] +matrix[9][322] * vector[9] +matrix[10][322] * vector[10] +matrix[11][322] * vector[11] +matrix[12][322] * vector[12] +matrix[13][322] * vector[13] +matrix[14][322] * vector[14] +matrix[15][322] * vector[15] +matrix[16][322] * vector[16] +matrix[17][322] * vector[17] +matrix[18][322] * vector[18] +matrix[19][322] * vector[19] +matrix[20][322] * vector[20] +matrix[21][322] * vector[21] +matrix[22][322] * vector[22] +matrix[23][322] * vector[23] +matrix[24][322] * vector[24] +matrix[25][322] * vector[25] +matrix[26][322] * vector[26] +matrix[27][322] * vector[27] +matrix[28][322] * vector[28] +matrix[29][322] * vector[29] +matrix[30][322] * vector[30] +matrix[31][322] * vector[31] +matrix[32][322] * vector[32] +matrix[33][322] * vector[33] +matrix[34][322] * vector[34] +matrix[35][322] * vector[35] +matrix[36][322] * vector[36] +matrix[37][322] * vector[37] +matrix[38][322] * vector[38] +matrix[39][322] * vector[39] +matrix[40][322] * vector[40] +matrix[41][322] * vector[41] +matrix[42][322] * vector[42] +matrix[43][322] * vector[43] +matrix[44][322] * vector[44] +matrix[45][322] * vector[45] +matrix[46][322] * vector[46] +matrix[47][322] * vector[47] +matrix[48][322] * vector[48] +matrix[49][322] * vector[49] +matrix[50][322] * vector[50] +matrix[51][322] * vector[51] +matrix[52][322] * vector[52] +matrix[53][322] * vector[53] +matrix[54][322] * vector[54] +matrix[55][322] * vector[55] +matrix[56][322] * vector[56] +matrix[57][322] * vector[57] +matrix[58][322] * vector[58] +matrix[59][322] * vector[59] +matrix[60][322] * vector[60] +matrix[61][322] * vector[61] +matrix[62][322] * vector[62] +matrix[63][322] * vector[63] +matrix[64][322] * vector[64] +matrix[65][322] * vector[65] +matrix[66][322] * vector[66] +matrix[67][322] * vector[67] +matrix[68][322] * vector[68] +matrix[69][322] * vector[69] +matrix[70][322] * vector[70] +matrix[71][322] * vector[71] +matrix[72][322] * vector[72] +matrix[73][322] * vector[73] +matrix[74][322] * vector[74] +matrix[75][322] * vector[75] +matrix[76][322] * vector[76] +matrix[77][322] * vector[77] +matrix[78][322] * vector[78] +matrix[79][322] * vector[79] +matrix[80][322] * vector[80] +matrix[81][322] * vector[81] +matrix[82][322] * vector[82] +matrix[83][322] * vector[83] +matrix[84][322] * vector[84] +matrix[85][322] * vector[85] +matrix[86][322] * vector[86] +matrix[87][322] * vector[87] +matrix[88][322] * vector[88] +matrix[89][322] * vector[89] +matrix[90][322] * vector[90] +matrix[91][322] * vector[91] +matrix[92][322] * vector[92] +matrix[93][322] * vector[93] +matrix[94][322] * vector[94] +matrix[95][322] * vector[95] +matrix[96][322] * vector[96] +matrix[97][322] * vector[97] +matrix[98][322] * vector[98] +matrix[99][322] * vector[99] +b[322];
assign result[323] = matrix[0][323] * vector[0] +matrix[1][323] * vector[1] +matrix[2][323] * vector[2] +matrix[3][323] * vector[3] +matrix[4][323] * vector[4] +matrix[5][323] * vector[5] +matrix[6][323] * vector[6] +matrix[7][323] * vector[7] +matrix[8][323] * vector[8] +matrix[9][323] * vector[9] +matrix[10][323] * vector[10] +matrix[11][323] * vector[11] +matrix[12][323] * vector[12] +matrix[13][323] * vector[13] +matrix[14][323] * vector[14] +matrix[15][323] * vector[15] +matrix[16][323] * vector[16] +matrix[17][323] * vector[17] +matrix[18][323] * vector[18] +matrix[19][323] * vector[19] +matrix[20][323] * vector[20] +matrix[21][323] * vector[21] +matrix[22][323] * vector[22] +matrix[23][323] * vector[23] +matrix[24][323] * vector[24] +matrix[25][323] * vector[25] +matrix[26][323] * vector[26] +matrix[27][323] * vector[27] +matrix[28][323] * vector[28] +matrix[29][323] * vector[29] +matrix[30][323] * vector[30] +matrix[31][323] * vector[31] +matrix[32][323] * vector[32] +matrix[33][323] * vector[33] +matrix[34][323] * vector[34] +matrix[35][323] * vector[35] +matrix[36][323] * vector[36] +matrix[37][323] * vector[37] +matrix[38][323] * vector[38] +matrix[39][323] * vector[39] +matrix[40][323] * vector[40] +matrix[41][323] * vector[41] +matrix[42][323] * vector[42] +matrix[43][323] * vector[43] +matrix[44][323] * vector[44] +matrix[45][323] * vector[45] +matrix[46][323] * vector[46] +matrix[47][323] * vector[47] +matrix[48][323] * vector[48] +matrix[49][323] * vector[49] +matrix[50][323] * vector[50] +matrix[51][323] * vector[51] +matrix[52][323] * vector[52] +matrix[53][323] * vector[53] +matrix[54][323] * vector[54] +matrix[55][323] * vector[55] +matrix[56][323] * vector[56] +matrix[57][323] * vector[57] +matrix[58][323] * vector[58] +matrix[59][323] * vector[59] +matrix[60][323] * vector[60] +matrix[61][323] * vector[61] +matrix[62][323] * vector[62] +matrix[63][323] * vector[63] +matrix[64][323] * vector[64] +matrix[65][323] * vector[65] +matrix[66][323] * vector[66] +matrix[67][323] * vector[67] +matrix[68][323] * vector[68] +matrix[69][323] * vector[69] +matrix[70][323] * vector[70] +matrix[71][323] * vector[71] +matrix[72][323] * vector[72] +matrix[73][323] * vector[73] +matrix[74][323] * vector[74] +matrix[75][323] * vector[75] +matrix[76][323] * vector[76] +matrix[77][323] * vector[77] +matrix[78][323] * vector[78] +matrix[79][323] * vector[79] +matrix[80][323] * vector[80] +matrix[81][323] * vector[81] +matrix[82][323] * vector[82] +matrix[83][323] * vector[83] +matrix[84][323] * vector[84] +matrix[85][323] * vector[85] +matrix[86][323] * vector[86] +matrix[87][323] * vector[87] +matrix[88][323] * vector[88] +matrix[89][323] * vector[89] +matrix[90][323] * vector[90] +matrix[91][323] * vector[91] +matrix[92][323] * vector[92] +matrix[93][323] * vector[93] +matrix[94][323] * vector[94] +matrix[95][323] * vector[95] +matrix[96][323] * vector[96] +matrix[97][323] * vector[97] +matrix[98][323] * vector[98] +matrix[99][323] * vector[99] +b[323];
assign result[324] = matrix[0][324] * vector[0] +matrix[1][324] * vector[1] +matrix[2][324] * vector[2] +matrix[3][324] * vector[3] +matrix[4][324] * vector[4] +matrix[5][324] * vector[5] +matrix[6][324] * vector[6] +matrix[7][324] * vector[7] +matrix[8][324] * vector[8] +matrix[9][324] * vector[9] +matrix[10][324] * vector[10] +matrix[11][324] * vector[11] +matrix[12][324] * vector[12] +matrix[13][324] * vector[13] +matrix[14][324] * vector[14] +matrix[15][324] * vector[15] +matrix[16][324] * vector[16] +matrix[17][324] * vector[17] +matrix[18][324] * vector[18] +matrix[19][324] * vector[19] +matrix[20][324] * vector[20] +matrix[21][324] * vector[21] +matrix[22][324] * vector[22] +matrix[23][324] * vector[23] +matrix[24][324] * vector[24] +matrix[25][324] * vector[25] +matrix[26][324] * vector[26] +matrix[27][324] * vector[27] +matrix[28][324] * vector[28] +matrix[29][324] * vector[29] +matrix[30][324] * vector[30] +matrix[31][324] * vector[31] +matrix[32][324] * vector[32] +matrix[33][324] * vector[33] +matrix[34][324] * vector[34] +matrix[35][324] * vector[35] +matrix[36][324] * vector[36] +matrix[37][324] * vector[37] +matrix[38][324] * vector[38] +matrix[39][324] * vector[39] +matrix[40][324] * vector[40] +matrix[41][324] * vector[41] +matrix[42][324] * vector[42] +matrix[43][324] * vector[43] +matrix[44][324] * vector[44] +matrix[45][324] * vector[45] +matrix[46][324] * vector[46] +matrix[47][324] * vector[47] +matrix[48][324] * vector[48] +matrix[49][324] * vector[49] +matrix[50][324] * vector[50] +matrix[51][324] * vector[51] +matrix[52][324] * vector[52] +matrix[53][324] * vector[53] +matrix[54][324] * vector[54] +matrix[55][324] * vector[55] +matrix[56][324] * vector[56] +matrix[57][324] * vector[57] +matrix[58][324] * vector[58] +matrix[59][324] * vector[59] +matrix[60][324] * vector[60] +matrix[61][324] * vector[61] +matrix[62][324] * vector[62] +matrix[63][324] * vector[63] +matrix[64][324] * vector[64] +matrix[65][324] * vector[65] +matrix[66][324] * vector[66] +matrix[67][324] * vector[67] +matrix[68][324] * vector[68] +matrix[69][324] * vector[69] +matrix[70][324] * vector[70] +matrix[71][324] * vector[71] +matrix[72][324] * vector[72] +matrix[73][324] * vector[73] +matrix[74][324] * vector[74] +matrix[75][324] * vector[75] +matrix[76][324] * vector[76] +matrix[77][324] * vector[77] +matrix[78][324] * vector[78] +matrix[79][324] * vector[79] +matrix[80][324] * vector[80] +matrix[81][324] * vector[81] +matrix[82][324] * vector[82] +matrix[83][324] * vector[83] +matrix[84][324] * vector[84] +matrix[85][324] * vector[85] +matrix[86][324] * vector[86] +matrix[87][324] * vector[87] +matrix[88][324] * vector[88] +matrix[89][324] * vector[89] +matrix[90][324] * vector[90] +matrix[91][324] * vector[91] +matrix[92][324] * vector[92] +matrix[93][324] * vector[93] +matrix[94][324] * vector[94] +matrix[95][324] * vector[95] +matrix[96][324] * vector[96] +matrix[97][324] * vector[97] +matrix[98][324] * vector[98] +matrix[99][324] * vector[99] +b[324];
assign result[325] = matrix[0][325] * vector[0] +matrix[1][325] * vector[1] +matrix[2][325] * vector[2] +matrix[3][325] * vector[3] +matrix[4][325] * vector[4] +matrix[5][325] * vector[5] +matrix[6][325] * vector[6] +matrix[7][325] * vector[7] +matrix[8][325] * vector[8] +matrix[9][325] * vector[9] +matrix[10][325] * vector[10] +matrix[11][325] * vector[11] +matrix[12][325] * vector[12] +matrix[13][325] * vector[13] +matrix[14][325] * vector[14] +matrix[15][325] * vector[15] +matrix[16][325] * vector[16] +matrix[17][325] * vector[17] +matrix[18][325] * vector[18] +matrix[19][325] * vector[19] +matrix[20][325] * vector[20] +matrix[21][325] * vector[21] +matrix[22][325] * vector[22] +matrix[23][325] * vector[23] +matrix[24][325] * vector[24] +matrix[25][325] * vector[25] +matrix[26][325] * vector[26] +matrix[27][325] * vector[27] +matrix[28][325] * vector[28] +matrix[29][325] * vector[29] +matrix[30][325] * vector[30] +matrix[31][325] * vector[31] +matrix[32][325] * vector[32] +matrix[33][325] * vector[33] +matrix[34][325] * vector[34] +matrix[35][325] * vector[35] +matrix[36][325] * vector[36] +matrix[37][325] * vector[37] +matrix[38][325] * vector[38] +matrix[39][325] * vector[39] +matrix[40][325] * vector[40] +matrix[41][325] * vector[41] +matrix[42][325] * vector[42] +matrix[43][325] * vector[43] +matrix[44][325] * vector[44] +matrix[45][325] * vector[45] +matrix[46][325] * vector[46] +matrix[47][325] * vector[47] +matrix[48][325] * vector[48] +matrix[49][325] * vector[49] +matrix[50][325] * vector[50] +matrix[51][325] * vector[51] +matrix[52][325] * vector[52] +matrix[53][325] * vector[53] +matrix[54][325] * vector[54] +matrix[55][325] * vector[55] +matrix[56][325] * vector[56] +matrix[57][325] * vector[57] +matrix[58][325] * vector[58] +matrix[59][325] * vector[59] +matrix[60][325] * vector[60] +matrix[61][325] * vector[61] +matrix[62][325] * vector[62] +matrix[63][325] * vector[63] +matrix[64][325] * vector[64] +matrix[65][325] * vector[65] +matrix[66][325] * vector[66] +matrix[67][325] * vector[67] +matrix[68][325] * vector[68] +matrix[69][325] * vector[69] +matrix[70][325] * vector[70] +matrix[71][325] * vector[71] +matrix[72][325] * vector[72] +matrix[73][325] * vector[73] +matrix[74][325] * vector[74] +matrix[75][325] * vector[75] +matrix[76][325] * vector[76] +matrix[77][325] * vector[77] +matrix[78][325] * vector[78] +matrix[79][325] * vector[79] +matrix[80][325] * vector[80] +matrix[81][325] * vector[81] +matrix[82][325] * vector[82] +matrix[83][325] * vector[83] +matrix[84][325] * vector[84] +matrix[85][325] * vector[85] +matrix[86][325] * vector[86] +matrix[87][325] * vector[87] +matrix[88][325] * vector[88] +matrix[89][325] * vector[89] +matrix[90][325] * vector[90] +matrix[91][325] * vector[91] +matrix[92][325] * vector[92] +matrix[93][325] * vector[93] +matrix[94][325] * vector[94] +matrix[95][325] * vector[95] +matrix[96][325] * vector[96] +matrix[97][325] * vector[97] +matrix[98][325] * vector[98] +matrix[99][325] * vector[99] +b[325];
assign result[326] = matrix[0][326] * vector[0] +matrix[1][326] * vector[1] +matrix[2][326] * vector[2] +matrix[3][326] * vector[3] +matrix[4][326] * vector[4] +matrix[5][326] * vector[5] +matrix[6][326] * vector[6] +matrix[7][326] * vector[7] +matrix[8][326] * vector[8] +matrix[9][326] * vector[9] +matrix[10][326] * vector[10] +matrix[11][326] * vector[11] +matrix[12][326] * vector[12] +matrix[13][326] * vector[13] +matrix[14][326] * vector[14] +matrix[15][326] * vector[15] +matrix[16][326] * vector[16] +matrix[17][326] * vector[17] +matrix[18][326] * vector[18] +matrix[19][326] * vector[19] +matrix[20][326] * vector[20] +matrix[21][326] * vector[21] +matrix[22][326] * vector[22] +matrix[23][326] * vector[23] +matrix[24][326] * vector[24] +matrix[25][326] * vector[25] +matrix[26][326] * vector[26] +matrix[27][326] * vector[27] +matrix[28][326] * vector[28] +matrix[29][326] * vector[29] +matrix[30][326] * vector[30] +matrix[31][326] * vector[31] +matrix[32][326] * vector[32] +matrix[33][326] * vector[33] +matrix[34][326] * vector[34] +matrix[35][326] * vector[35] +matrix[36][326] * vector[36] +matrix[37][326] * vector[37] +matrix[38][326] * vector[38] +matrix[39][326] * vector[39] +matrix[40][326] * vector[40] +matrix[41][326] * vector[41] +matrix[42][326] * vector[42] +matrix[43][326] * vector[43] +matrix[44][326] * vector[44] +matrix[45][326] * vector[45] +matrix[46][326] * vector[46] +matrix[47][326] * vector[47] +matrix[48][326] * vector[48] +matrix[49][326] * vector[49] +matrix[50][326] * vector[50] +matrix[51][326] * vector[51] +matrix[52][326] * vector[52] +matrix[53][326] * vector[53] +matrix[54][326] * vector[54] +matrix[55][326] * vector[55] +matrix[56][326] * vector[56] +matrix[57][326] * vector[57] +matrix[58][326] * vector[58] +matrix[59][326] * vector[59] +matrix[60][326] * vector[60] +matrix[61][326] * vector[61] +matrix[62][326] * vector[62] +matrix[63][326] * vector[63] +matrix[64][326] * vector[64] +matrix[65][326] * vector[65] +matrix[66][326] * vector[66] +matrix[67][326] * vector[67] +matrix[68][326] * vector[68] +matrix[69][326] * vector[69] +matrix[70][326] * vector[70] +matrix[71][326] * vector[71] +matrix[72][326] * vector[72] +matrix[73][326] * vector[73] +matrix[74][326] * vector[74] +matrix[75][326] * vector[75] +matrix[76][326] * vector[76] +matrix[77][326] * vector[77] +matrix[78][326] * vector[78] +matrix[79][326] * vector[79] +matrix[80][326] * vector[80] +matrix[81][326] * vector[81] +matrix[82][326] * vector[82] +matrix[83][326] * vector[83] +matrix[84][326] * vector[84] +matrix[85][326] * vector[85] +matrix[86][326] * vector[86] +matrix[87][326] * vector[87] +matrix[88][326] * vector[88] +matrix[89][326] * vector[89] +matrix[90][326] * vector[90] +matrix[91][326] * vector[91] +matrix[92][326] * vector[92] +matrix[93][326] * vector[93] +matrix[94][326] * vector[94] +matrix[95][326] * vector[95] +matrix[96][326] * vector[96] +matrix[97][326] * vector[97] +matrix[98][326] * vector[98] +matrix[99][326] * vector[99] +b[326];
assign result[327] = matrix[0][327] * vector[0] +matrix[1][327] * vector[1] +matrix[2][327] * vector[2] +matrix[3][327] * vector[3] +matrix[4][327] * vector[4] +matrix[5][327] * vector[5] +matrix[6][327] * vector[6] +matrix[7][327] * vector[7] +matrix[8][327] * vector[8] +matrix[9][327] * vector[9] +matrix[10][327] * vector[10] +matrix[11][327] * vector[11] +matrix[12][327] * vector[12] +matrix[13][327] * vector[13] +matrix[14][327] * vector[14] +matrix[15][327] * vector[15] +matrix[16][327] * vector[16] +matrix[17][327] * vector[17] +matrix[18][327] * vector[18] +matrix[19][327] * vector[19] +matrix[20][327] * vector[20] +matrix[21][327] * vector[21] +matrix[22][327] * vector[22] +matrix[23][327] * vector[23] +matrix[24][327] * vector[24] +matrix[25][327] * vector[25] +matrix[26][327] * vector[26] +matrix[27][327] * vector[27] +matrix[28][327] * vector[28] +matrix[29][327] * vector[29] +matrix[30][327] * vector[30] +matrix[31][327] * vector[31] +matrix[32][327] * vector[32] +matrix[33][327] * vector[33] +matrix[34][327] * vector[34] +matrix[35][327] * vector[35] +matrix[36][327] * vector[36] +matrix[37][327] * vector[37] +matrix[38][327] * vector[38] +matrix[39][327] * vector[39] +matrix[40][327] * vector[40] +matrix[41][327] * vector[41] +matrix[42][327] * vector[42] +matrix[43][327] * vector[43] +matrix[44][327] * vector[44] +matrix[45][327] * vector[45] +matrix[46][327] * vector[46] +matrix[47][327] * vector[47] +matrix[48][327] * vector[48] +matrix[49][327] * vector[49] +matrix[50][327] * vector[50] +matrix[51][327] * vector[51] +matrix[52][327] * vector[52] +matrix[53][327] * vector[53] +matrix[54][327] * vector[54] +matrix[55][327] * vector[55] +matrix[56][327] * vector[56] +matrix[57][327] * vector[57] +matrix[58][327] * vector[58] +matrix[59][327] * vector[59] +matrix[60][327] * vector[60] +matrix[61][327] * vector[61] +matrix[62][327] * vector[62] +matrix[63][327] * vector[63] +matrix[64][327] * vector[64] +matrix[65][327] * vector[65] +matrix[66][327] * vector[66] +matrix[67][327] * vector[67] +matrix[68][327] * vector[68] +matrix[69][327] * vector[69] +matrix[70][327] * vector[70] +matrix[71][327] * vector[71] +matrix[72][327] * vector[72] +matrix[73][327] * vector[73] +matrix[74][327] * vector[74] +matrix[75][327] * vector[75] +matrix[76][327] * vector[76] +matrix[77][327] * vector[77] +matrix[78][327] * vector[78] +matrix[79][327] * vector[79] +matrix[80][327] * vector[80] +matrix[81][327] * vector[81] +matrix[82][327] * vector[82] +matrix[83][327] * vector[83] +matrix[84][327] * vector[84] +matrix[85][327] * vector[85] +matrix[86][327] * vector[86] +matrix[87][327] * vector[87] +matrix[88][327] * vector[88] +matrix[89][327] * vector[89] +matrix[90][327] * vector[90] +matrix[91][327] * vector[91] +matrix[92][327] * vector[92] +matrix[93][327] * vector[93] +matrix[94][327] * vector[94] +matrix[95][327] * vector[95] +matrix[96][327] * vector[96] +matrix[97][327] * vector[97] +matrix[98][327] * vector[98] +matrix[99][327] * vector[99] +b[327];
assign result[328] = matrix[0][328] * vector[0] +matrix[1][328] * vector[1] +matrix[2][328] * vector[2] +matrix[3][328] * vector[3] +matrix[4][328] * vector[4] +matrix[5][328] * vector[5] +matrix[6][328] * vector[6] +matrix[7][328] * vector[7] +matrix[8][328] * vector[8] +matrix[9][328] * vector[9] +matrix[10][328] * vector[10] +matrix[11][328] * vector[11] +matrix[12][328] * vector[12] +matrix[13][328] * vector[13] +matrix[14][328] * vector[14] +matrix[15][328] * vector[15] +matrix[16][328] * vector[16] +matrix[17][328] * vector[17] +matrix[18][328] * vector[18] +matrix[19][328] * vector[19] +matrix[20][328] * vector[20] +matrix[21][328] * vector[21] +matrix[22][328] * vector[22] +matrix[23][328] * vector[23] +matrix[24][328] * vector[24] +matrix[25][328] * vector[25] +matrix[26][328] * vector[26] +matrix[27][328] * vector[27] +matrix[28][328] * vector[28] +matrix[29][328] * vector[29] +matrix[30][328] * vector[30] +matrix[31][328] * vector[31] +matrix[32][328] * vector[32] +matrix[33][328] * vector[33] +matrix[34][328] * vector[34] +matrix[35][328] * vector[35] +matrix[36][328] * vector[36] +matrix[37][328] * vector[37] +matrix[38][328] * vector[38] +matrix[39][328] * vector[39] +matrix[40][328] * vector[40] +matrix[41][328] * vector[41] +matrix[42][328] * vector[42] +matrix[43][328] * vector[43] +matrix[44][328] * vector[44] +matrix[45][328] * vector[45] +matrix[46][328] * vector[46] +matrix[47][328] * vector[47] +matrix[48][328] * vector[48] +matrix[49][328] * vector[49] +matrix[50][328] * vector[50] +matrix[51][328] * vector[51] +matrix[52][328] * vector[52] +matrix[53][328] * vector[53] +matrix[54][328] * vector[54] +matrix[55][328] * vector[55] +matrix[56][328] * vector[56] +matrix[57][328] * vector[57] +matrix[58][328] * vector[58] +matrix[59][328] * vector[59] +matrix[60][328] * vector[60] +matrix[61][328] * vector[61] +matrix[62][328] * vector[62] +matrix[63][328] * vector[63] +matrix[64][328] * vector[64] +matrix[65][328] * vector[65] +matrix[66][328] * vector[66] +matrix[67][328] * vector[67] +matrix[68][328] * vector[68] +matrix[69][328] * vector[69] +matrix[70][328] * vector[70] +matrix[71][328] * vector[71] +matrix[72][328] * vector[72] +matrix[73][328] * vector[73] +matrix[74][328] * vector[74] +matrix[75][328] * vector[75] +matrix[76][328] * vector[76] +matrix[77][328] * vector[77] +matrix[78][328] * vector[78] +matrix[79][328] * vector[79] +matrix[80][328] * vector[80] +matrix[81][328] * vector[81] +matrix[82][328] * vector[82] +matrix[83][328] * vector[83] +matrix[84][328] * vector[84] +matrix[85][328] * vector[85] +matrix[86][328] * vector[86] +matrix[87][328] * vector[87] +matrix[88][328] * vector[88] +matrix[89][328] * vector[89] +matrix[90][328] * vector[90] +matrix[91][328] * vector[91] +matrix[92][328] * vector[92] +matrix[93][328] * vector[93] +matrix[94][328] * vector[94] +matrix[95][328] * vector[95] +matrix[96][328] * vector[96] +matrix[97][328] * vector[97] +matrix[98][328] * vector[98] +matrix[99][328] * vector[99] +b[328];
assign result[329] = matrix[0][329] * vector[0] +matrix[1][329] * vector[1] +matrix[2][329] * vector[2] +matrix[3][329] * vector[3] +matrix[4][329] * vector[4] +matrix[5][329] * vector[5] +matrix[6][329] * vector[6] +matrix[7][329] * vector[7] +matrix[8][329] * vector[8] +matrix[9][329] * vector[9] +matrix[10][329] * vector[10] +matrix[11][329] * vector[11] +matrix[12][329] * vector[12] +matrix[13][329] * vector[13] +matrix[14][329] * vector[14] +matrix[15][329] * vector[15] +matrix[16][329] * vector[16] +matrix[17][329] * vector[17] +matrix[18][329] * vector[18] +matrix[19][329] * vector[19] +matrix[20][329] * vector[20] +matrix[21][329] * vector[21] +matrix[22][329] * vector[22] +matrix[23][329] * vector[23] +matrix[24][329] * vector[24] +matrix[25][329] * vector[25] +matrix[26][329] * vector[26] +matrix[27][329] * vector[27] +matrix[28][329] * vector[28] +matrix[29][329] * vector[29] +matrix[30][329] * vector[30] +matrix[31][329] * vector[31] +matrix[32][329] * vector[32] +matrix[33][329] * vector[33] +matrix[34][329] * vector[34] +matrix[35][329] * vector[35] +matrix[36][329] * vector[36] +matrix[37][329] * vector[37] +matrix[38][329] * vector[38] +matrix[39][329] * vector[39] +matrix[40][329] * vector[40] +matrix[41][329] * vector[41] +matrix[42][329] * vector[42] +matrix[43][329] * vector[43] +matrix[44][329] * vector[44] +matrix[45][329] * vector[45] +matrix[46][329] * vector[46] +matrix[47][329] * vector[47] +matrix[48][329] * vector[48] +matrix[49][329] * vector[49] +matrix[50][329] * vector[50] +matrix[51][329] * vector[51] +matrix[52][329] * vector[52] +matrix[53][329] * vector[53] +matrix[54][329] * vector[54] +matrix[55][329] * vector[55] +matrix[56][329] * vector[56] +matrix[57][329] * vector[57] +matrix[58][329] * vector[58] +matrix[59][329] * vector[59] +matrix[60][329] * vector[60] +matrix[61][329] * vector[61] +matrix[62][329] * vector[62] +matrix[63][329] * vector[63] +matrix[64][329] * vector[64] +matrix[65][329] * vector[65] +matrix[66][329] * vector[66] +matrix[67][329] * vector[67] +matrix[68][329] * vector[68] +matrix[69][329] * vector[69] +matrix[70][329] * vector[70] +matrix[71][329] * vector[71] +matrix[72][329] * vector[72] +matrix[73][329] * vector[73] +matrix[74][329] * vector[74] +matrix[75][329] * vector[75] +matrix[76][329] * vector[76] +matrix[77][329] * vector[77] +matrix[78][329] * vector[78] +matrix[79][329] * vector[79] +matrix[80][329] * vector[80] +matrix[81][329] * vector[81] +matrix[82][329] * vector[82] +matrix[83][329] * vector[83] +matrix[84][329] * vector[84] +matrix[85][329] * vector[85] +matrix[86][329] * vector[86] +matrix[87][329] * vector[87] +matrix[88][329] * vector[88] +matrix[89][329] * vector[89] +matrix[90][329] * vector[90] +matrix[91][329] * vector[91] +matrix[92][329] * vector[92] +matrix[93][329] * vector[93] +matrix[94][329] * vector[94] +matrix[95][329] * vector[95] +matrix[96][329] * vector[96] +matrix[97][329] * vector[97] +matrix[98][329] * vector[98] +matrix[99][329] * vector[99] +b[329];
assign result[330] = matrix[0][330] * vector[0] +matrix[1][330] * vector[1] +matrix[2][330] * vector[2] +matrix[3][330] * vector[3] +matrix[4][330] * vector[4] +matrix[5][330] * vector[5] +matrix[6][330] * vector[6] +matrix[7][330] * vector[7] +matrix[8][330] * vector[8] +matrix[9][330] * vector[9] +matrix[10][330] * vector[10] +matrix[11][330] * vector[11] +matrix[12][330] * vector[12] +matrix[13][330] * vector[13] +matrix[14][330] * vector[14] +matrix[15][330] * vector[15] +matrix[16][330] * vector[16] +matrix[17][330] * vector[17] +matrix[18][330] * vector[18] +matrix[19][330] * vector[19] +matrix[20][330] * vector[20] +matrix[21][330] * vector[21] +matrix[22][330] * vector[22] +matrix[23][330] * vector[23] +matrix[24][330] * vector[24] +matrix[25][330] * vector[25] +matrix[26][330] * vector[26] +matrix[27][330] * vector[27] +matrix[28][330] * vector[28] +matrix[29][330] * vector[29] +matrix[30][330] * vector[30] +matrix[31][330] * vector[31] +matrix[32][330] * vector[32] +matrix[33][330] * vector[33] +matrix[34][330] * vector[34] +matrix[35][330] * vector[35] +matrix[36][330] * vector[36] +matrix[37][330] * vector[37] +matrix[38][330] * vector[38] +matrix[39][330] * vector[39] +matrix[40][330] * vector[40] +matrix[41][330] * vector[41] +matrix[42][330] * vector[42] +matrix[43][330] * vector[43] +matrix[44][330] * vector[44] +matrix[45][330] * vector[45] +matrix[46][330] * vector[46] +matrix[47][330] * vector[47] +matrix[48][330] * vector[48] +matrix[49][330] * vector[49] +matrix[50][330] * vector[50] +matrix[51][330] * vector[51] +matrix[52][330] * vector[52] +matrix[53][330] * vector[53] +matrix[54][330] * vector[54] +matrix[55][330] * vector[55] +matrix[56][330] * vector[56] +matrix[57][330] * vector[57] +matrix[58][330] * vector[58] +matrix[59][330] * vector[59] +matrix[60][330] * vector[60] +matrix[61][330] * vector[61] +matrix[62][330] * vector[62] +matrix[63][330] * vector[63] +matrix[64][330] * vector[64] +matrix[65][330] * vector[65] +matrix[66][330] * vector[66] +matrix[67][330] * vector[67] +matrix[68][330] * vector[68] +matrix[69][330] * vector[69] +matrix[70][330] * vector[70] +matrix[71][330] * vector[71] +matrix[72][330] * vector[72] +matrix[73][330] * vector[73] +matrix[74][330] * vector[74] +matrix[75][330] * vector[75] +matrix[76][330] * vector[76] +matrix[77][330] * vector[77] +matrix[78][330] * vector[78] +matrix[79][330] * vector[79] +matrix[80][330] * vector[80] +matrix[81][330] * vector[81] +matrix[82][330] * vector[82] +matrix[83][330] * vector[83] +matrix[84][330] * vector[84] +matrix[85][330] * vector[85] +matrix[86][330] * vector[86] +matrix[87][330] * vector[87] +matrix[88][330] * vector[88] +matrix[89][330] * vector[89] +matrix[90][330] * vector[90] +matrix[91][330] * vector[91] +matrix[92][330] * vector[92] +matrix[93][330] * vector[93] +matrix[94][330] * vector[94] +matrix[95][330] * vector[95] +matrix[96][330] * vector[96] +matrix[97][330] * vector[97] +matrix[98][330] * vector[98] +matrix[99][330] * vector[99] +b[330];
assign result[331] = matrix[0][331] * vector[0] +matrix[1][331] * vector[1] +matrix[2][331] * vector[2] +matrix[3][331] * vector[3] +matrix[4][331] * vector[4] +matrix[5][331] * vector[5] +matrix[6][331] * vector[6] +matrix[7][331] * vector[7] +matrix[8][331] * vector[8] +matrix[9][331] * vector[9] +matrix[10][331] * vector[10] +matrix[11][331] * vector[11] +matrix[12][331] * vector[12] +matrix[13][331] * vector[13] +matrix[14][331] * vector[14] +matrix[15][331] * vector[15] +matrix[16][331] * vector[16] +matrix[17][331] * vector[17] +matrix[18][331] * vector[18] +matrix[19][331] * vector[19] +matrix[20][331] * vector[20] +matrix[21][331] * vector[21] +matrix[22][331] * vector[22] +matrix[23][331] * vector[23] +matrix[24][331] * vector[24] +matrix[25][331] * vector[25] +matrix[26][331] * vector[26] +matrix[27][331] * vector[27] +matrix[28][331] * vector[28] +matrix[29][331] * vector[29] +matrix[30][331] * vector[30] +matrix[31][331] * vector[31] +matrix[32][331] * vector[32] +matrix[33][331] * vector[33] +matrix[34][331] * vector[34] +matrix[35][331] * vector[35] +matrix[36][331] * vector[36] +matrix[37][331] * vector[37] +matrix[38][331] * vector[38] +matrix[39][331] * vector[39] +matrix[40][331] * vector[40] +matrix[41][331] * vector[41] +matrix[42][331] * vector[42] +matrix[43][331] * vector[43] +matrix[44][331] * vector[44] +matrix[45][331] * vector[45] +matrix[46][331] * vector[46] +matrix[47][331] * vector[47] +matrix[48][331] * vector[48] +matrix[49][331] * vector[49] +matrix[50][331] * vector[50] +matrix[51][331] * vector[51] +matrix[52][331] * vector[52] +matrix[53][331] * vector[53] +matrix[54][331] * vector[54] +matrix[55][331] * vector[55] +matrix[56][331] * vector[56] +matrix[57][331] * vector[57] +matrix[58][331] * vector[58] +matrix[59][331] * vector[59] +matrix[60][331] * vector[60] +matrix[61][331] * vector[61] +matrix[62][331] * vector[62] +matrix[63][331] * vector[63] +matrix[64][331] * vector[64] +matrix[65][331] * vector[65] +matrix[66][331] * vector[66] +matrix[67][331] * vector[67] +matrix[68][331] * vector[68] +matrix[69][331] * vector[69] +matrix[70][331] * vector[70] +matrix[71][331] * vector[71] +matrix[72][331] * vector[72] +matrix[73][331] * vector[73] +matrix[74][331] * vector[74] +matrix[75][331] * vector[75] +matrix[76][331] * vector[76] +matrix[77][331] * vector[77] +matrix[78][331] * vector[78] +matrix[79][331] * vector[79] +matrix[80][331] * vector[80] +matrix[81][331] * vector[81] +matrix[82][331] * vector[82] +matrix[83][331] * vector[83] +matrix[84][331] * vector[84] +matrix[85][331] * vector[85] +matrix[86][331] * vector[86] +matrix[87][331] * vector[87] +matrix[88][331] * vector[88] +matrix[89][331] * vector[89] +matrix[90][331] * vector[90] +matrix[91][331] * vector[91] +matrix[92][331] * vector[92] +matrix[93][331] * vector[93] +matrix[94][331] * vector[94] +matrix[95][331] * vector[95] +matrix[96][331] * vector[96] +matrix[97][331] * vector[97] +matrix[98][331] * vector[98] +matrix[99][331] * vector[99] +b[331];
assign result[332] = matrix[0][332] * vector[0] +matrix[1][332] * vector[1] +matrix[2][332] * vector[2] +matrix[3][332] * vector[3] +matrix[4][332] * vector[4] +matrix[5][332] * vector[5] +matrix[6][332] * vector[6] +matrix[7][332] * vector[7] +matrix[8][332] * vector[8] +matrix[9][332] * vector[9] +matrix[10][332] * vector[10] +matrix[11][332] * vector[11] +matrix[12][332] * vector[12] +matrix[13][332] * vector[13] +matrix[14][332] * vector[14] +matrix[15][332] * vector[15] +matrix[16][332] * vector[16] +matrix[17][332] * vector[17] +matrix[18][332] * vector[18] +matrix[19][332] * vector[19] +matrix[20][332] * vector[20] +matrix[21][332] * vector[21] +matrix[22][332] * vector[22] +matrix[23][332] * vector[23] +matrix[24][332] * vector[24] +matrix[25][332] * vector[25] +matrix[26][332] * vector[26] +matrix[27][332] * vector[27] +matrix[28][332] * vector[28] +matrix[29][332] * vector[29] +matrix[30][332] * vector[30] +matrix[31][332] * vector[31] +matrix[32][332] * vector[32] +matrix[33][332] * vector[33] +matrix[34][332] * vector[34] +matrix[35][332] * vector[35] +matrix[36][332] * vector[36] +matrix[37][332] * vector[37] +matrix[38][332] * vector[38] +matrix[39][332] * vector[39] +matrix[40][332] * vector[40] +matrix[41][332] * vector[41] +matrix[42][332] * vector[42] +matrix[43][332] * vector[43] +matrix[44][332] * vector[44] +matrix[45][332] * vector[45] +matrix[46][332] * vector[46] +matrix[47][332] * vector[47] +matrix[48][332] * vector[48] +matrix[49][332] * vector[49] +matrix[50][332] * vector[50] +matrix[51][332] * vector[51] +matrix[52][332] * vector[52] +matrix[53][332] * vector[53] +matrix[54][332] * vector[54] +matrix[55][332] * vector[55] +matrix[56][332] * vector[56] +matrix[57][332] * vector[57] +matrix[58][332] * vector[58] +matrix[59][332] * vector[59] +matrix[60][332] * vector[60] +matrix[61][332] * vector[61] +matrix[62][332] * vector[62] +matrix[63][332] * vector[63] +matrix[64][332] * vector[64] +matrix[65][332] * vector[65] +matrix[66][332] * vector[66] +matrix[67][332] * vector[67] +matrix[68][332] * vector[68] +matrix[69][332] * vector[69] +matrix[70][332] * vector[70] +matrix[71][332] * vector[71] +matrix[72][332] * vector[72] +matrix[73][332] * vector[73] +matrix[74][332] * vector[74] +matrix[75][332] * vector[75] +matrix[76][332] * vector[76] +matrix[77][332] * vector[77] +matrix[78][332] * vector[78] +matrix[79][332] * vector[79] +matrix[80][332] * vector[80] +matrix[81][332] * vector[81] +matrix[82][332] * vector[82] +matrix[83][332] * vector[83] +matrix[84][332] * vector[84] +matrix[85][332] * vector[85] +matrix[86][332] * vector[86] +matrix[87][332] * vector[87] +matrix[88][332] * vector[88] +matrix[89][332] * vector[89] +matrix[90][332] * vector[90] +matrix[91][332] * vector[91] +matrix[92][332] * vector[92] +matrix[93][332] * vector[93] +matrix[94][332] * vector[94] +matrix[95][332] * vector[95] +matrix[96][332] * vector[96] +matrix[97][332] * vector[97] +matrix[98][332] * vector[98] +matrix[99][332] * vector[99] +b[332];
assign result[333] = matrix[0][333] * vector[0] +matrix[1][333] * vector[1] +matrix[2][333] * vector[2] +matrix[3][333] * vector[3] +matrix[4][333] * vector[4] +matrix[5][333] * vector[5] +matrix[6][333] * vector[6] +matrix[7][333] * vector[7] +matrix[8][333] * vector[8] +matrix[9][333] * vector[9] +matrix[10][333] * vector[10] +matrix[11][333] * vector[11] +matrix[12][333] * vector[12] +matrix[13][333] * vector[13] +matrix[14][333] * vector[14] +matrix[15][333] * vector[15] +matrix[16][333] * vector[16] +matrix[17][333] * vector[17] +matrix[18][333] * vector[18] +matrix[19][333] * vector[19] +matrix[20][333] * vector[20] +matrix[21][333] * vector[21] +matrix[22][333] * vector[22] +matrix[23][333] * vector[23] +matrix[24][333] * vector[24] +matrix[25][333] * vector[25] +matrix[26][333] * vector[26] +matrix[27][333] * vector[27] +matrix[28][333] * vector[28] +matrix[29][333] * vector[29] +matrix[30][333] * vector[30] +matrix[31][333] * vector[31] +matrix[32][333] * vector[32] +matrix[33][333] * vector[33] +matrix[34][333] * vector[34] +matrix[35][333] * vector[35] +matrix[36][333] * vector[36] +matrix[37][333] * vector[37] +matrix[38][333] * vector[38] +matrix[39][333] * vector[39] +matrix[40][333] * vector[40] +matrix[41][333] * vector[41] +matrix[42][333] * vector[42] +matrix[43][333] * vector[43] +matrix[44][333] * vector[44] +matrix[45][333] * vector[45] +matrix[46][333] * vector[46] +matrix[47][333] * vector[47] +matrix[48][333] * vector[48] +matrix[49][333] * vector[49] +matrix[50][333] * vector[50] +matrix[51][333] * vector[51] +matrix[52][333] * vector[52] +matrix[53][333] * vector[53] +matrix[54][333] * vector[54] +matrix[55][333] * vector[55] +matrix[56][333] * vector[56] +matrix[57][333] * vector[57] +matrix[58][333] * vector[58] +matrix[59][333] * vector[59] +matrix[60][333] * vector[60] +matrix[61][333] * vector[61] +matrix[62][333] * vector[62] +matrix[63][333] * vector[63] +matrix[64][333] * vector[64] +matrix[65][333] * vector[65] +matrix[66][333] * vector[66] +matrix[67][333] * vector[67] +matrix[68][333] * vector[68] +matrix[69][333] * vector[69] +matrix[70][333] * vector[70] +matrix[71][333] * vector[71] +matrix[72][333] * vector[72] +matrix[73][333] * vector[73] +matrix[74][333] * vector[74] +matrix[75][333] * vector[75] +matrix[76][333] * vector[76] +matrix[77][333] * vector[77] +matrix[78][333] * vector[78] +matrix[79][333] * vector[79] +matrix[80][333] * vector[80] +matrix[81][333] * vector[81] +matrix[82][333] * vector[82] +matrix[83][333] * vector[83] +matrix[84][333] * vector[84] +matrix[85][333] * vector[85] +matrix[86][333] * vector[86] +matrix[87][333] * vector[87] +matrix[88][333] * vector[88] +matrix[89][333] * vector[89] +matrix[90][333] * vector[90] +matrix[91][333] * vector[91] +matrix[92][333] * vector[92] +matrix[93][333] * vector[93] +matrix[94][333] * vector[94] +matrix[95][333] * vector[95] +matrix[96][333] * vector[96] +matrix[97][333] * vector[97] +matrix[98][333] * vector[98] +matrix[99][333] * vector[99] +b[333];
assign result[334] = matrix[0][334] * vector[0] +matrix[1][334] * vector[1] +matrix[2][334] * vector[2] +matrix[3][334] * vector[3] +matrix[4][334] * vector[4] +matrix[5][334] * vector[5] +matrix[6][334] * vector[6] +matrix[7][334] * vector[7] +matrix[8][334] * vector[8] +matrix[9][334] * vector[9] +matrix[10][334] * vector[10] +matrix[11][334] * vector[11] +matrix[12][334] * vector[12] +matrix[13][334] * vector[13] +matrix[14][334] * vector[14] +matrix[15][334] * vector[15] +matrix[16][334] * vector[16] +matrix[17][334] * vector[17] +matrix[18][334] * vector[18] +matrix[19][334] * vector[19] +matrix[20][334] * vector[20] +matrix[21][334] * vector[21] +matrix[22][334] * vector[22] +matrix[23][334] * vector[23] +matrix[24][334] * vector[24] +matrix[25][334] * vector[25] +matrix[26][334] * vector[26] +matrix[27][334] * vector[27] +matrix[28][334] * vector[28] +matrix[29][334] * vector[29] +matrix[30][334] * vector[30] +matrix[31][334] * vector[31] +matrix[32][334] * vector[32] +matrix[33][334] * vector[33] +matrix[34][334] * vector[34] +matrix[35][334] * vector[35] +matrix[36][334] * vector[36] +matrix[37][334] * vector[37] +matrix[38][334] * vector[38] +matrix[39][334] * vector[39] +matrix[40][334] * vector[40] +matrix[41][334] * vector[41] +matrix[42][334] * vector[42] +matrix[43][334] * vector[43] +matrix[44][334] * vector[44] +matrix[45][334] * vector[45] +matrix[46][334] * vector[46] +matrix[47][334] * vector[47] +matrix[48][334] * vector[48] +matrix[49][334] * vector[49] +matrix[50][334] * vector[50] +matrix[51][334] * vector[51] +matrix[52][334] * vector[52] +matrix[53][334] * vector[53] +matrix[54][334] * vector[54] +matrix[55][334] * vector[55] +matrix[56][334] * vector[56] +matrix[57][334] * vector[57] +matrix[58][334] * vector[58] +matrix[59][334] * vector[59] +matrix[60][334] * vector[60] +matrix[61][334] * vector[61] +matrix[62][334] * vector[62] +matrix[63][334] * vector[63] +matrix[64][334] * vector[64] +matrix[65][334] * vector[65] +matrix[66][334] * vector[66] +matrix[67][334] * vector[67] +matrix[68][334] * vector[68] +matrix[69][334] * vector[69] +matrix[70][334] * vector[70] +matrix[71][334] * vector[71] +matrix[72][334] * vector[72] +matrix[73][334] * vector[73] +matrix[74][334] * vector[74] +matrix[75][334] * vector[75] +matrix[76][334] * vector[76] +matrix[77][334] * vector[77] +matrix[78][334] * vector[78] +matrix[79][334] * vector[79] +matrix[80][334] * vector[80] +matrix[81][334] * vector[81] +matrix[82][334] * vector[82] +matrix[83][334] * vector[83] +matrix[84][334] * vector[84] +matrix[85][334] * vector[85] +matrix[86][334] * vector[86] +matrix[87][334] * vector[87] +matrix[88][334] * vector[88] +matrix[89][334] * vector[89] +matrix[90][334] * vector[90] +matrix[91][334] * vector[91] +matrix[92][334] * vector[92] +matrix[93][334] * vector[93] +matrix[94][334] * vector[94] +matrix[95][334] * vector[95] +matrix[96][334] * vector[96] +matrix[97][334] * vector[97] +matrix[98][334] * vector[98] +matrix[99][334] * vector[99] +b[334];
assign result[335] = matrix[0][335] * vector[0] +matrix[1][335] * vector[1] +matrix[2][335] * vector[2] +matrix[3][335] * vector[3] +matrix[4][335] * vector[4] +matrix[5][335] * vector[5] +matrix[6][335] * vector[6] +matrix[7][335] * vector[7] +matrix[8][335] * vector[8] +matrix[9][335] * vector[9] +matrix[10][335] * vector[10] +matrix[11][335] * vector[11] +matrix[12][335] * vector[12] +matrix[13][335] * vector[13] +matrix[14][335] * vector[14] +matrix[15][335] * vector[15] +matrix[16][335] * vector[16] +matrix[17][335] * vector[17] +matrix[18][335] * vector[18] +matrix[19][335] * vector[19] +matrix[20][335] * vector[20] +matrix[21][335] * vector[21] +matrix[22][335] * vector[22] +matrix[23][335] * vector[23] +matrix[24][335] * vector[24] +matrix[25][335] * vector[25] +matrix[26][335] * vector[26] +matrix[27][335] * vector[27] +matrix[28][335] * vector[28] +matrix[29][335] * vector[29] +matrix[30][335] * vector[30] +matrix[31][335] * vector[31] +matrix[32][335] * vector[32] +matrix[33][335] * vector[33] +matrix[34][335] * vector[34] +matrix[35][335] * vector[35] +matrix[36][335] * vector[36] +matrix[37][335] * vector[37] +matrix[38][335] * vector[38] +matrix[39][335] * vector[39] +matrix[40][335] * vector[40] +matrix[41][335] * vector[41] +matrix[42][335] * vector[42] +matrix[43][335] * vector[43] +matrix[44][335] * vector[44] +matrix[45][335] * vector[45] +matrix[46][335] * vector[46] +matrix[47][335] * vector[47] +matrix[48][335] * vector[48] +matrix[49][335] * vector[49] +matrix[50][335] * vector[50] +matrix[51][335] * vector[51] +matrix[52][335] * vector[52] +matrix[53][335] * vector[53] +matrix[54][335] * vector[54] +matrix[55][335] * vector[55] +matrix[56][335] * vector[56] +matrix[57][335] * vector[57] +matrix[58][335] * vector[58] +matrix[59][335] * vector[59] +matrix[60][335] * vector[60] +matrix[61][335] * vector[61] +matrix[62][335] * vector[62] +matrix[63][335] * vector[63] +matrix[64][335] * vector[64] +matrix[65][335] * vector[65] +matrix[66][335] * vector[66] +matrix[67][335] * vector[67] +matrix[68][335] * vector[68] +matrix[69][335] * vector[69] +matrix[70][335] * vector[70] +matrix[71][335] * vector[71] +matrix[72][335] * vector[72] +matrix[73][335] * vector[73] +matrix[74][335] * vector[74] +matrix[75][335] * vector[75] +matrix[76][335] * vector[76] +matrix[77][335] * vector[77] +matrix[78][335] * vector[78] +matrix[79][335] * vector[79] +matrix[80][335] * vector[80] +matrix[81][335] * vector[81] +matrix[82][335] * vector[82] +matrix[83][335] * vector[83] +matrix[84][335] * vector[84] +matrix[85][335] * vector[85] +matrix[86][335] * vector[86] +matrix[87][335] * vector[87] +matrix[88][335] * vector[88] +matrix[89][335] * vector[89] +matrix[90][335] * vector[90] +matrix[91][335] * vector[91] +matrix[92][335] * vector[92] +matrix[93][335] * vector[93] +matrix[94][335] * vector[94] +matrix[95][335] * vector[95] +matrix[96][335] * vector[96] +matrix[97][335] * vector[97] +matrix[98][335] * vector[98] +matrix[99][335] * vector[99] +b[335];
assign result[336] = matrix[0][336] * vector[0] +matrix[1][336] * vector[1] +matrix[2][336] * vector[2] +matrix[3][336] * vector[3] +matrix[4][336] * vector[4] +matrix[5][336] * vector[5] +matrix[6][336] * vector[6] +matrix[7][336] * vector[7] +matrix[8][336] * vector[8] +matrix[9][336] * vector[9] +matrix[10][336] * vector[10] +matrix[11][336] * vector[11] +matrix[12][336] * vector[12] +matrix[13][336] * vector[13] +matrix[14][336] * vector[14] +matrix[15][336] * vector[15] +matrix[16][336] * vector[16] +matrix[17][336] * vector[17] +matrix[18][336] * vector[18] +matrix[19][336] * vector[19] +matrix[20][336] * vector[20] +matrix[21][336] * vector[21] +matrix[22][336] * vector[22] +matrix[23][336] * vector[23] +matrix[24][336] * vector[24] +matrix[25][336] * vector[25] +matrix[26][336] * vector[26] +matrix[27][336] * vector[27] +matrix[28][336] * vector[28] +matrix[29][336] * vector[29] +matrix[30][336] * vector[30] +matrix[31][336] * vector[31] +matrix[32][336] * vector[32] +matrix[33][336] * vector[33] +matrix[34][336] * vector[34] +matrix[35][336] * vector[35] +matrix[36][336] * vector[36] +matrix[37][336] * vector[37] +matrix[38][336] * vector[38] +matrix[39][336] * vector[39] +matrix[40][336] * vector[40] +matrix[41][336] * vector[41] +matrix[42][336] * vector[42] +matrix[43][336] * vector[43] +matrix[44][336] * vector[44] +matrix[45][336] * vector[45] +matrix[46][336] * vector[46] +matrix[47][336] * vector[47] +matrix[48][336] * vector[48] +matrix[49][336] * vector[49] +matrix[50][336] * vector[50] +matrix[51][336] * vector[51] +matrix[52][336] * vector[52] +matrix[53][336] * vector[53] +matrix[54][336] * vector[54] +matrix[55][336] * vector[55] +matrix[56][336] * vector[56] +matrix[57][336] * vector[57] +matrix[58][336] * vector[58] +matrix[59][336] * vector[59] +matrix[60][336] * vector[60] +matrix[61][336] * vector[61] +matrix[62][336] * vector[62] +matrix[63][336] * vector[63] +matrix[64][336] * vector[64] +matrix[65][336] * vector[65] +matrix[66][336] * vector[66] +matrix[67][336] * vector[67] +matrix[68][336] * vector[68] +matrix[69][336] * vector[69] +matrix[70][336] * vector[70] +matrix[71][336] * vector[71] +matrix[72][336] * vector[72] +matrix[73][336] * vector[73] +matrix[74][336] * vector[74] +matrix[75][336] * vector[75] +matrix[76][336] * vector[76] +matrix[77][336] * vector[77] +matrix[78][336] * vector[78] +matrix[79][336] * vector[79] +matrix[80][336] * vector[80] +matrix[81][336] * vector[81] +matrix[82][336] * vector[82] +matrix[83][336] * vector[83] +matrix[84][336] * vector[84] +matrix[85][336] * vector[85] +matrix[86][336] * vector[86] +matrix[87][336] * vector[87] +matrix[88][336] * vector[88] +matrix[89][336] * vector[89] +matrix[90][336] * vector[90] +matrix[91][336] * vector[91] +matrix[92][336] * vector[92] +matrix[93][336] * vector[93] +matrix[94][336] * vector[94] +matrix[95][336] * vector[95] +matrix[96][336] * vector[96] +matrix[97][336] * vector[97] +matrix[98][336] * vector[98] +matrix[99][336] * vector[99] +b[336];
assign result[337] = matrix[0][337] * vector[0] +matrix[1][337] * vector[1] +matrix[2][337] * vector[2] +matrix[3][337] * vector[3] +matrix[4][337] * vector[4] +matrix[5][337] * vector[5] +matrix[6][337] * vector[6] +matrix[7][337] * vector[7] +matrix[8][337] * vector[8] +matrix[9][337] * vector[9] +matrix[10][337] * vector[10] +matrix[11][337] * vector[11] +matrix[12][337] * vector[12] +matrix[13][337] * vector[13] +matrix[14][337] * vector[14] +matrix[15][337] * vector[15] +matrix[16][337] * vector[16] +matrix[17][337] * vector[17] +matrix[18][337] * vector[18] +matrix[19][337] * vector[19] +matrix[20][337] * vector[20] +matrix[21][337] * vector[21] +matrix[22][337] * vector[22] +matrix[23][337] * vector[23] +matrix[24][337] * vector[24] +matrix[25][337] * vector[25] +matrix[26][337] * vector[26] +matrix[27][337] * vector[27] +matrix[28][337] * vector[28] +matrix[29][337] * vector[29] +matrix[30][337] * vector[30] +matrix[31][337] * vector[31] +matrix[32][337] * vector[32] +matrix[33][337] * vector[33] +matrix[34][337] * vector[34] +matrix[35][337] * vector[35] +matrix[36][337] * vector[36] +matrix[37][337] * vector[37] +matrix[38][337] * vector[38] +matrix[39][337] * vector[39] +matrix[40][337] * vector[40] +matrix[41][337] * vector[41] +matrix[42][337] * vector[42] +matrix[43][337] * vector[43] +matrix[44][337] * vector[44] +matrix[45][337] * vector[45] +matrix[46][337] * vector[46] +matrix[47][337] * vector[47] +matrix[48][337] * vector[48] +matrix[49][337] * vector[49] +matrix[50][337] * vector[50] +matrix[51][337] * vector[51] +matrix[52][337] * vector[52] +matrix[53][337] * vector[53] +matrix[54][337] * vector[54] +matrix[55][337] * vector[55] +matrix[56][337] * vector[56] +matrix[57][337] * vector[57] +matrix[58][337] * vector[58] +matrix[59][337] * vector[59] +matrix[60][337] * vector[60] +matrix[61][337] * vector[61] +matrix[62][337] * vector[62] +matrix[63][337] * vector[63] +matrix[64][337] * vector[64] +matrix[65][337] * vector[65] +matrix[66][337] * vector[66] +matrix[67][337] * vector[67] +matrix[68][337] * vector[68] +matrix[69][337] * vector[69] +matrix[70][337] * vector[70] +matrix[71][337] * vector[71] +matrix[72][337] * vector[72] +matrix[73][337] * vector[73] +matrix[74][337] * vector[74] +matrix[75][337] * vector[75] +matrix[76][337] * vector[76] +matrix[77][337] * vector[77] +matrix[78][337] * vector[78] +matrix[79][337] * vector[79] +matrix[80][337] * vector[80] +matrix[81][337] * vector[81] +matrix[82][337] * vector[82] +matrix[83][337] * vector[83] +matrix[84][337] * vector[84] +matrix[85][337] * vector[85] +matrix[86][337] * vector[86] +matrix[87][337] * vector[87] +matrix[88][337] * vector[88] +matrix[89][337] * vector[89] +matrix[90][337] * vector[90] +matrix[91][337] * vector[91] +matrix[92][337] * vector[92] +matrix[93][337] * vector[93] +matrix[94][337] * vector[94] +matrix[95][337] * vector[95] +matrix[96][337] * vector[96] +matrix[97][337] * vector[97] +matrix[98][337] * vector[98] +matrix[99][337] * vector[99] +b[337];
assign result[338] = matrix[0][338] * vector[0] +matrix[1][338] * vector[1] +matrix[2][338] * vector[2] +matrix[3][338] * vector[3] +matrix[4][338] * vector[4] +matrix[5][338] * vector[5] +matrix[6][338] * vector[6] +matrix[7][338] * vector[7] +matrix[8][338] * vector[8] +matrix[9][338] * vector[9] +matrix[10][338] * vector[10] +matrix[11][338] * vector[11] +matrix[12][338] * vector[12] +matrix[13][338] * vector[13] +matrix[14][338] * vector[14] +matrix[15][338] * vector[15] +matrix[16][338] * vector[16] +matrix[17][338] * vector[17] +matrix[18][338] * vector[18] +matrix[19][338] * vector[19] +matrix[20][338] * vector[20] +matrix[21][338] * vector[21] +matrix[22][338] * vector[22] +matrix[23][338] * vector[23] +matrix[24][338] * vector[24] +matrix[25][338] * vector[25] +matrix[26][338] * vector[26] +matrix[27][338] * vector[27] +matrix[28][338] * vector[28] +matrix[29][338] * vector[29] +matrix[30][338] * vector[30] +matrix[31][338] * vector[31] +matrix[32][338] * vector[32] +matrix[33][338] * vector[33] +matrix[34][338] * vector[34] +matrix[35][338] * vector[35] +matrix[36][338] * vector[36] +matrix[37][338] * vector[37] +matrix[38][338] * vector[38] +matrix[39][338] * vector[39] +matrix[40][338] * vector[40] +matrix[41][338] * vector[41] +matrix[42][338] * vector[42] +matrix[43][338] * vector[43] +matrix[44][338] * vector[44] +matrix[45][338] * vector[45] +matrix[46][338] * vector[46] +matrix[47][338] * vector[47] +matrix[48][338] * vector[48] +matrix[49][338] * vector[49] +matrix[50][338] * vector[50] +matrix[51][338] * vector[51] +matrix[52][338] * vector[52] +matrix[53][338] * vector[53] +matrix[54][338] * vector[54] +matrix[55][338] * vector[55] +matrix[56][338] * vector[56] +matrix[57][338] * vector[57] +matrix[58][338] * vector[58] +matrix[59][338] * vector[59] +matrix[60][338] * vector[60] +matrix[61][338] * vector[61] +matrix[62][338] * vector[62] +matrix[63][338] * vector[63] +matrix[64][338] * vector[64] +matrix[65][338] * vector[65] +matrix[66][338] * vector[66] +matrix[67][338] * vector[67] +matrix[68][338] * vector[68] +matrix[69][338] * vector[69] +matrix[70][338] * vector[70] +matrix[71][338] * vector[71] +matrix[72][338] * vector[72] +matrix[73][338] * vector[73] +matrix[74][338] * vector[74] +matrix[75][338] * vector[75] +matrix[76][338] * vector[76] +matrix[77][338] * vector[77] +matrix[78][338] * vector[78] +matrix[79][338] * vector[79] +matrix[80][338] * vector[80] +matrix[81][338] * vector[81] +matrix[82][338] * vector[82] +matrix[83][338] * vector[83] +matrix[84][338] * vector[84] +matrix[85][338] * vector[85] +matrix[86][338] * vector[86] +matrix[87][338] * vector[87] +matrix[88][338] * vector[88] +matrix[89][338] * vector[89] +matrix[90][338] * vector[90] +matrix[91][338] * vector[91] +matrix[92][338] * vector[92] +matrix[93][338] * vector[93] +matrix[94][338] * vector[94] +matrix[95][338] * vector[95] +matrix[96][338] * vector[96] +matrix[97][338] * vector[97] +matrix[98][338] * vector[98] +matrix[99][338] * vector[99] +b[338];
assign result[339] = matrix[0][339] * vector[0] +matrix[1][339] * vector[1] +matrix[2][339] * vector[2] +matrix[3][339] * vector[3] +matrix[4][339] * vector[4] +matrix[5][339] * vector[5] +matrix[6][339] * vector[6] +matrix[7][339] * vector[7] +matrix[8][339] * vector[8] +matrix[9][339] * vector[9] +matrix[10][339] * vector[10] +matrix[11][339] * vector[11] +matrix[12][339] * vector[12] +matrix[13][339] * vector[13] +matrix[14][339] * vector[14] +matrix[15][339] * vector[15] +matrix[16][339] * vector[16] +matrix[17][339] * vector[17] +matrix[18][339] * vector[18] +matrix[19][339] * vector[19] +matrix[20][339] * vector[20] +matrix[21][339] * vector[21] +matrix[22][339] * vector[22] +matrix[23][339] * vector[23] +matrix[24][339] * vector[24] +matrix[25][339] * vector[25] +matrix[26][339] * vector[26] +matrix[27][339] * vector[27] +matrix[28][339] * vector[28] +matrix[29][339] * vector[29] +matrix[30][339] * vector[30] +matrix[31][339] * vector[31] +matrix[32][339] * vector[32] +matrix[33][339] * vector[33] +matrix[34][339] * vector[34] +matrix[35][339] * vector[35] +matrix[36][339] * vector[36] +matrix[37][339] * vector[37] +matrix[38][339] * vector[38] +matrix[39][339] * vector[39] +matrix[40][339] * vector[40] +matrix[41][339] * vector[41] +matrix[42][339] * vector[42] +matrix[43][339] * vector[43] +matrix[44][339] * vector[44] +matrix[45][339] * vector[45] +matrix[46][339] * vector[46] +matrix[47][339] * vector[47] +matrix[48][339] * vector[48] +matrix[49][339] * vector[49] +matrix[50][339] * vector[50] +matrix[51][339] * vector[51] +matrix[52][339] * vector[52] +matrix[53][339] * vector[53] +matrix[54][339] * vector[54] +matrix[55][339] * vector[55] +matrix[56][339] * vector[56] +matrix[57][339] * vector[57] +matrix[58][339] * vector[58] +matrix[59][339] * vector[59] +matrix[60][339] * vector[60] +matrix[61][339] * vector[61] +matrix[62][339] * vector[62] +matrix[63][339] * vector[63] +matrix[64][339] * vector[64] +matrix[65][339] * vector[65] +matrix[66][339] * vector[66] +matrix[67][339] * vector[67] +matrix[68][339] * vector[68] +matrix[69][339] * vector[69] +matrix[70][339] * vector[70] +matrix[71][339] * vector[71] +matrix[72][339] * vector[72] +matrix[73][339] * vector[73] +matrix[74][339] * vector[74] +matrix[75][339] * vector[75] +matrix[76][339] * vector[76] +matrix[77][339] * vector[77] +matrix[78][339] * vector[78] +matrix[79][339] * vector[79] +matrix[80][339] * vector[80] +matrix[81][339] * vector[81] +matrix[82][339] * vector[82] +matrix[83][339] * vector[83] +matrix[84][339] * vector[84] +matrix[85][339] * vector[85] +matrix[86][339] * vector[86] +matrix[87][339] * vector[87] +matrix[88][339] * vector[88] +matrix[89][339] * vector[89] +matrix[90][339] * vector[90] +matrix[91][339] * vector[91] +matrix[92][339] * vector[92] +matrix[93][339] * vector[93] +matrix[94][339] * vector[94] +matrix[95][339] * vector[95] +matrix[96][339] * vector[96] +matrix[97][339] * vector[97] +matrix[98][339] * vector[98] +matrix[99][339] * vector[99] +b[339];
assign result[340] = matrix[0][340] * vector[0] +matrix[1][340] * vector[1] +matrix[2][340] * vector[2] +matrix[3][340] * vector[3] +matrix[4][340] * vector[4] +matrix[5][340] * vector[5] +matrix[6][340] * vector[6] +matrix[7][340] * vector[7] +matrix[8][340] * vector[8] +matrix[9][340] * vector[9] +matrix[10][340] * vector[10] +matrix[11][340] * vector[11] +matrix[12][340] * vector[12] +matrix[13][340] * vector[13] +matrix[14][340] * vector[14] +matrix[15][340] * vector[15] +matrix[16][340] * vector[16] +matrix[17][340] * vector[17] +matrix[18][340] * vector[18] +matrix[19][340] * vector[19] +matrix[20][340] * vector[20] +matrix[21][340] * vector[21] +matrix[22][340] * vector[22] +matrix[23][340] * vector[23] +matrix[24][340] * vector[24] +matrix[25][340] * vector[25] +matrix[26][340] * vector[26] +matrix[27][340] * vector[27] +matrix[28][340] * vector[28] +matrix[29][340] * vector[29] +matrix[30][340] * vector[30] +matrix[31][340] * vector[31] +matrix[32][340] * vector[32] +matrix[33][340] * vector[33] +matrix[34][340] * vector[34] +matrix[35][340] * vector[35] +matrix[36][340] * vector[36] +matrix[37][340] * vector[37] +matrix[38][340] * vector[38] +matrix[39][340] * vector[39] +matrix[40][340] * vector[40] +matrix[41][340] * vector[41] +matrix[42][340] * vector[42] +matrix[43][340] * vector[43] +matrix[44][340] * vector[44] +matrix[45][340] * vector[45] +matrix[46][340] * vector[46] +matrix[47][340] * vector[47] +matrix[48][340] * vector[48] +matrix[49][340] * vector[49] +matrix[50][340] * vector[50] +matrix[51][340] * vector[51] +matrix[52][340] * vector[52] +matrix[53][340] * vector[53] +matrix[54][340] * vector[54] +matrix[55][340] * vector[55] +matrix[56][340] * vector[56] +matrix[57][340] * vector[57] +matrix[58][340] * vector[58] +matrix[59][340] * vector[59] +matrix[60][340] * vector[60] +matrix[61][340] * vector[61] +matrix[62][340] * vector[62] +matrix[63][340] * vector[63] +matrix[64][340] * vector[64] +matrix[65][340] * vector[65] +matrix[66][340] * vector[66] +matrix[67][340] * vector[67] +matrix[68][340] * vector[68] +matrix[69][340] * vector[69] +matrix[70][340] * vector[70] +matrix[71][340] * vector[71] +matrix[72][340] * vector[72] +matrix[73][340] * vector[73] +matrix[74][340] * vector[74] +matrix[75][340] * vector[75] +matrix[76][340] * vector[76] +matrix[77][340] * vector[77] +matrix[78][340] * vector[78] +matrix[79][340] * vector[79] +matrix[80][340] * vector[80] +matrix[81][340] * vector[81] +matrix[82][340] * vector[82] +matrix[83][340] * vector[83] +matrix[84][340] * vector[84] +matrix[85][340] * vector[85] +matrix[86][340] * vector[86] +matrix[87][340] * vector[87] +matrix[88][340] * vector[88] +matrix[89][340] * vector[89] +matrix[90][340] * vector[90] +matrix[91][340] * vector[91] +matrix[92][340] * vector[92] +matrix[93][340] * vector[93] +matrix[94][340] * vector[94] +matrix[95][340] * vector[95] +matrix[96][340] * vector[96] +matrix[97][340] * vector[97] +matrix[98][340] * vector[98] +matrix[99][340] * vector[99] +b[340];
assign result[341] = matrix[0][341] * vector[0] +matrix[1][341] * vector[1] +matrix[2][341] * vector[2] +matrix[3][341] * vector[3] +matrix[4][341] * vector[4] +matrix[5][341] * vector[5] +matrix[6][341] * vector[6] +matrix[7][341] * vector[7] +matrix[8][341] * vector[8] +matrix[9][341] * vector[9] +matrix[10][341] * vector[10] +matrix[11][341] * vector[11] +matrix[12][341] * vector[12] +matrix[13][341] * vector[13] +matrix[14][341] * vector[14] +matrix[15][341] * vector[15] +matrix[16][341] * vector[16] +matrix[17][341] * vector[17] +matrix[18][341] * vector[18] +matrix[19][341] * vector[19] +matrix[20][341] * vector[20] +matrix[21][341] * vector[21] +matrix[22][341] * vector[22] +matrix[23][341] * vector[23] +matrix[24][341] * vector[24] +matrix[25][341] * vector[25] +matrix[26][341] * vector[26] +matrix[27][341] * vector[27] +matrix[28][341] * vector[28] +matrix[29][341] * vector[29] +matrix[30][341] * vector[30] +matrix[31][341] * vector[31] +matrix[32][341] * vector[32] +matrix[33][341] * vector[33] +matrix[34][341] * vector[34] +matrix[35][341] * vector[35] +matrix[36][341] * vector[36] +matrix[37][341] * vector[37] +matrix[38][341] * vector[38] +matrix[39][341] * vector[39] +matrix[40][341] * vector[40] +matrix[41][341] * vector[41] +matrix[42][341] * vector[42] +matrix[43][341] * vector[43] +matrix[44][341] * vector[44] +matrix[45][341] * vector[45] +matrix[46][341] * vector[46] +matrix[47][341] * vector[47] +matrix[48][341] * vector[48] +matrix[49][341] * vector[49] +matrix[50][341] * vector[50] +matrix[51][341] * vector[51] +matrix[52][341] * vector[52] +matrix[53][341] * vector[53] +matrix[54][341] * vector[54] +matrix[55][341] * vector[55] +matrix[56][341] * vector[56] +matrix[57][341] * vector[57] +matrix[58][341] * vector[58] +matrix[59][341] * vector[59] +matrix[60][341] * vector[60] +matrix[61][341] * vector[61] +matrix[62][341] * vector[62] +matrix[63][341] * vector[63] +matrix[64][341] * vector[64] +matrix[65][341] * vector[65] +matrix[66][341] * vector[66] +matrix[67][341] * vector[67] +matrix[68][341] * vector[68] +matrix[69][341] * vector[69] +matrix[70][341] * vector[70] +matrix[71][341] * vector[71] +matrix[72][341] * vector[72] +matrix[73][341] * vector[73] +matrix[74][341] * vector[74] +matrix[75][341] * vector[75] +matrix[76][341] * vector[76] +matrix[77][341] * vector[77] +matrix[78][341] * vector[78] +matrix[79][341] * vector[79] +matrix[80][341] * vector[80] +matrix[81][341] * vector[81] +matrix[82][341] * vector[82] +matrix[83][341] * vector[83] +matrix[84][341] * vector[84] +matrix[85][341] * vector[85] +matrix[86][341] * vector[86] +matrix[87][341] * vector[87] +matrix[88][341] * vector[88] +matrix[89][341] * vector[89] +matrix[90][341] * vector[90] +matrix[91][341] * vector[91] +matrix[92][341] * vector[92] +matrix[93][341] * vector[93] +matrix[94][341] * vector[94] +matrix[95][341] * vector[95] +matrix[96][341] * vector[96] +matrix[97][341] * vector[97] +matrix[98][341] * vector[98] +matrix[99][341] * vector[99] +b[341];
assign result[342] = matrix[0][342] * vector[0] +matrix[1][342] * vector[1] +matrix[2][342] * vector[2] +matrix[3][342] * vector[3] +matrix[4][342] * vector[4] +matrix[5][342] * vector[5] +matrix[6][342] * vector[6] +matrix[7][342] * vector[7] +matrix[8][342] * vector[8] +matrix[9][342] * vector[9] +matrix[10][342] * vector[10] +matrix[11][342] * vector[11] +matrix[12][342] * vector[12] +matrix[13][342] * vector[13] +matrix[14][342] * vector[14] +matrix[15][342] * vector[15] +matrix[16][342] * vector[16] +matrix[17][342] * vector[17] +matrix[18][342] * vector[18] +matrix[19][342] * vector[19] +matrix[20][342] * vector[20] +matrix[21][342] * vector[21] +matrix[22][342] * vector[22] +matrix[23][342] * vector[23] +matrix[24][342] * vector[24] +matrix[25][342] * vector[25] +matrix[26][342] * vector[26] +matrix[27][342] * vector[27] +matrix[28][342] * vector[28] +matrix[29][342] * vector[29] +matrix[30][342] * vector[30] +matrix[31][342] * vector[31] +matrix[32][342] * vector[32] +matrix[33][342] * vector[33] +matrix[34][342] * vector[34] +matrix[35][342] * vector[35] +matrix[36][342] * vector[36] +matrix[37][342] * vector[37] +matrix[38][342] * vector[38] +matrix[39][342] * vector[39] +matrix[40][342] * vector[40] +matrix[41][342] * vector[41] +matrix[42][342] * vector[42] +matrix[43][342] * vector[43] +matrix[44][342] * vector[44] +matrix[45][342] * vector[45] +matrix[46][342] * vector[46] +matrix[47][342] * vector[47] +matrix[48][342] * vector[48] +matrix[49][342] * vector[49] +matrix[50][342] * vector[50] +matrix[51][342] * vector[51] +matrix[52][342] * vector[52] +matrix[53][342] * vector[53] +matrix[54][342] * vector[54] +matrix[55][342] * vector[55] +matrix[56][342] * vector[56] +matrix[57][342] * vector[57] +matrix[58][342] * vector[58] +matrix[59][342] * vector[59] +matrix[60][342] * vector[60] +matrix[61][342] * vector[61] +matrix[62][342] * vector[62] +matrix[63][342] * vector[63] +matrix[64][342] * vector[64] +matrix[65][342] * vector[65] +matrix[66][342] * vector[66] +matrix[67][342] * vector[67] +matrix[68][342] * vector[68] +matrix[69][342] * vector[69] +matrix[70][342] * vector[70] +matrix[71][342] * vector[71] +matrix[72][342] * vector[72] +matrix[73][342] * vector[73] +matrix[74][342] * vector[74] +matrix[75][342] * vector[75] +matrix[76][342] * vector[76] +matrix[77][342] * vector[77] +matrix[78][342] * vector[78] +matrix[79][342] * vector[79] +matrix[80][342] * vector[80] +matrix[81][342] * vector[81] +matrix[82][342] * vector[82] +matrix[83][342] * vector[83] +matrix[84][342] * vector[84] +matrix[85][342] * vector[85] +matrix[86][342] * vector[86] +matrix[87][342] * vector[87] +matrix[88][342] * vector[88] +matrix[89][342] * vector[89] +matrix[90][342] * vector[90] +matrix[91][342] * vector[91] +matrix[92][342] * vector[92] +matrix[93][342] * vector[93] +matrix[94][342] * vector[94] +matrix[95][342] * vector[95] +matrix[96][342] * vector[96] +matrix[97][342] * vector[97] +matrix[98][342] * vector[98] +matrix[99][342] * vector[99] +b[342];
assign result[343] = matrix[0][343] * vector[0] +matrix[1][343] * vector[1] +matrix[2][343] * vector[2] +matrix[3][343] * vector[3] +matrix[4][343] * vector[4] +matrix[5][343] * vector[5] +matrix[6][343] * vector[6] +matrix[7][343] * vector[7] +matrix[8][343] * vector[8] +matrix[9][343] * vector[9] +matrix[10][343] * vector[10] +matrix[11][343] * vector[11] +matrix[12][343] * vector[12] +matrix[13][343] * vector[13] +matrix[14][343] * vector[14] +matrix[15][343] * vector[15] +matrix[16][343] * vector[16] +matrix[17][343] * vector[17] +matrix[18][343] * vector[18] +matrix[19][343] * vector[19] +matrix[20][343] * vector[20] +matrix[21][343] * vector[21] +matrix[22][343] * vector[22] +matrix[23][343] * vector[23] +matrix[24][343] * vector[24] +matrix[25][343] * vector[25] +matrix[26][343] * vector[26] +matrix[27][343] * vector[27] +matrix[28][343] * vector[28] +matrix[29][343] * vector[29] +matrix[30][343] * vector[30] +matrix[31][343] * vector[31] +matrix[32][343] * vector[32] +matrix[33][343] * vector[33] +matrix[34][343] * vector[34] +matrix[35][343] * vector[35] +matrix[36][343] * vector[36] +matrix[37][343] * vector[37] +matrix[38][343] * vector[38] +matrix[39][343] * vector[39] +matrix[40][343] * vector[40] +matrix[41][343] * vector[41] +matrix[42][343] * vector[42] +matrix[43][343] * vector[43] +matrix[44][343] * vector[44] +matrix[45][343] * vector[45] +matrix[46][343] * vector[46] +matrix[47][343] * vector[47] +matrix[48][343] * vector[48] +matrix[49][343] * vector[49] +matrix[50][343] * vector[50] +matrix[51][343] * vector[51] +matrix[52][343] * vector[52] +matrix[53][343] * vector[53] +matrix[54][343] * vector[54] +matrix[55][343] * vector[55] +matrix[56][343] * vector[56] +matrix[57][343] * vector[57] +matrix[58][343] * vector[58] +matrix[59][343] * vector[59] +matrix[60][343] * vector[60] +matrix[61][343] * vector[61] +matrix[62][343] * vector[62] +matrix[63][343] * vector[63] +matrix[64][343] * vector[64] +matrix[65][343] * vector[65] +matrix[66][343] * vector[66] +matrix[67][343] * vector[67] +matrix[68][343] * vector[68] +matrix[69][343] * vector[69] +matrix[70][343] * vector[70] +matrix[71][343] * vector[71] +matrix[72][343] * vector[72] +matrix[73][343] * vector[73] +matrix[74][343] * vector[74] +matrix[75][343] * vector[75] +matrix[76][343] * vector[76] +matrix[77][343] * vector[77] +matrix[78][343] * vector[78] +matrix[79][343] * vector[79] +matrix[80][343] * vector[80] +matrix[81][343] * vector[81] +matrix[82][343] * vector[82] +matrix[83][343] * vector[83] +matrix[84][343] * vector[84] +matrix[85][343] * vector[85] +matrix[86][343] * vector[86] +matrix[87][343] * vector[87] +matrix[88][343] * vector[88] +matrix[89][343] * vector[89] +matrix[90][343] * vector[90] +matrix[91][343] * vector[91] +matrix[92][343] * vector[92] +matrix[93][343] * vector[93] +matrix[94][343] * vector[94] +matrix[95][343] * vector[95] +matrix[96][343] * vector[96] +matrix[97][343] * vector[97] +matrix[98][343] * vector[98] +matrix[99][343] * vector[99] +b[343];
assign result[344] = matrix[0][344] * vector[0] +matrix[1][344] * vector[1] +matrix[2][344] * vector[2] +matrix[3][344] * vector[3] +matrix[4][344] * vector[4] +matrix[5][344] * vector[5] +matrix[6][344] * vector[6] +matrix[7][344] * vector[7] +matrix[8][344] * vector[8] +matrix[9][344] * vector[9] +matrix[10][344] * vector[10] +matrix[11][344] * vector[11] +matrix[12][344] * vector[12] +matrix[13][344] * vector[13] +matrix[14][344] * vector[14] +matrix[15][344] * vector[15] +matrix[16][344] * vector[16] +matrix[17][344] * vector[17] +matrix[18][344] * vector[18] +matrix[19][344] * vector[19] +matrix[20][344] * vector[20] +matrix[21][344] * vector[21] +matrix[22][344] * vector[22] +matrix[23][344] * vector[23] +matrix[24][344] * vector[24] +matrix[25][344] * vector[25] +matrix[26][344] * vector[26] +matrix[27][344] * vector[27] +matrix[28][344] * vector[28] +matrix[29][344] * vector[29] +matrix[30][344] * vector[30] +matrix[31][344] * vector[31] +matrix[32][344] * vector[32] +matrix[33][344] * vector[33] +matrix[34][344] * vector[34] +matrix[35][344] * vector[35] +matrix[36][344] * vector[36] +matrix[37][344] * vector[37] +matrix[38][344] * vector[38] +matrix[39][344] * vector[39] +matrix[40][344] * vector[40] +matrix[41][344] * vector[41] +matrix[42][344] * vector[42] +matrix[43][344] * vector[43] +matrix[44][344] * vector[44] +matrix[45][344] * vector[45] +matrix[46][344] * vector[46] +matrix[47][344] * vector[47] +matrix[48][344] * vector[48] +matrix[49][344] * vector[49] +matrix[50][344] * vector[50] +matrix[51][344] * vector[51] +matrix[52][344] * vector[52] +matrix[53][344] * vector[53] +matrix[54][344] * vector[54] +matrix[55][344] * vector[55] +matrix[56][344] * vector[56] +matrix[57][344] * vector[57] +matrix[58][344] * vector[58] +matrix[59][344] * vector[59] +matrix[60][344] * vector[60] +matrix[61][344] * vector[61] +matrix[62][344] * vector[62] +matrix[63][344] * vector[63] +matrix[64][344] * vector[64] +matrix[65][344] * vector[65] +matrix[66][344] * vector[66] +matrix[67][344] * vector[67] +matrix[68][344] * vector[68] +matrix[69][344] * vector[69] +matrix[70][344] * vector[70] +matrix[71][344] * vector[71] +matrix[72][344] * vector[72] +matrix[73][344] * vector[73] +matrix[74][344] * vector[74] +matrix[75][344] * vector[75] +matrix[76][344] * vector[76] +matrix[77][344] * vector[77] +matrix[78][344] * vector[78] +matrix[79][344] * vector[79] +matrix[80][344] * vector[80] +matrix[81][344] * vector[81] +matrix[82][344] * vector[82] +matrix[83][344] * vector[83] +matrix[84][344] * vector[84] +matrix[85][344] * vector[85] +matrix[86][344] * vector[86] +matrix[87][344] * vector[87] +matrix[88][344] * vector[88] +matrix[89][344] * vector[89] +matrix[90][344] * vector[90] +matrix[91][344] * vector[91] +matrix[92][344] * vector[92] +matrix[93][344] * vector[93] +matrix[94][344] * vector[94] +matrix[95][344] * vector[95] +matrix[96][344] * vector[96] +matrix[97][344] * vector[97] +matrix[98][344] * vector[98] +matrix[99][344] * vector[99] +b[344];
assign result[345] = matrix[0][345] * vector[0] +matrix[1][345] * vector[1] +matrix[2][345] * vector[2] +matrix[3][345] * vector[3] +matrix[4][345] * vector[4] +matrix[5][345] * vector[5] +matrix[6][345] * vector[6] +matrix[7][345] * vector[7] +matrix[8][345] * vector[8] +matrix[9][345] * vector[9] +matrix[10][345] * vector[10] +matrix[11][345] * vector[11] +matrix[12][345] * vector[12] +matrix[13][345] * vector[13] +matrix[14][345] * vector[14] +matrix[15][345] * vector[15] +matrix[16][345] * vector[16] +matrix[17][345] * vector[17] +matrix[18][345] * vector[18] +matrix[19][345] * vector[19] +matrix[20][345] * vector[20] +matrix[21][345] * vector[21] +matrix[22][345] * vector[22] +matrix[23][345] * vector[23] +matrix[24][345] * vector[24] +matrix[25][345] * vector[25] +matrix[26][345] * vector[26] +matrix[27][345] * vector[27] +matrix[28][345] * vector[28] +matrix[29][345] * vector[29] +matrix[30][345] * vector[30] +matrix[31][345] * vector[31] +matrix[32][345] * vector[32] +matrix[33][345] * vector[33] +matrix[34][345] * vector[34] +matrix[35][345] * vector[35] +matrix[36][345] * vector[36] +matrix[37][345] * vector[37] +matrix[38][345] * vector[38] +matrix[39][345] * vector[39] +matrix[40][345] * vector[40] +matrix[41][345] * vector[41] +matrix[42][345] * vector[42] +matrix[43][345] * vector[43] +matrix[44][345] * vector[44] +matrix[45][345] * vector[45] +matrix[46][345] * vector[46] +matrix[47][345] * vector[47] +matrix[48][345] * vector[48] +matrix[49][345] * vector[49] +matrix[50][345] * vector[50] +matrix[51][345] * vector[51] +matrix[52][345] * vector[52] +matrix[53][345] * vector[53] +matrix[54][345] * vector[54] +matrix[55][345] * vector[55] +matrix[56][345] * vector[56] +matrix[57][345] * vector[57] +matrix[58][345] * vector[58] +matrix[59][345] * vector[59] +matrix[60][345] * vector[60] +matrix[61][345] * vector[61] +matrix[62][345] * vector[62] +matrix[63][345] * vector[63] +matrix[64][345] * vector[64] +matrix[65][345] * vector[65] +matrix[66][345] * vector[66] +matrix[67][345] * vector[67] +matrix[68][345] * vector[68] +matrix[69][345] * vector[69] +matrix[70][345] * vector[70] +matrix[71][345] * vector[71] +matrix[72][345] * vector[72] +matrix[73][345] * vector[73] +matrix[74][345] * vector[74] +matrix[75][345] * vector[75] +matrix[76][345] * vector[76] +matrix[77][345] * vector[77] +matrix[78][345] * vector[78] +matrix[79][345] * vector[79] +matrix[80][345] * vector[80] +matrix[81][345] * vector[81] +matrix[82][345] * vector[82] +matrix[83][345] * vector[83] +matrix[84][345] * vector[84] +matrix[85][345] * vector[85] +matrix[86][345] * vector[86] +matrix[87][345] * vector[87] +matrix[88][345] * vector[88] +matrix[89][345] * vector[89] +matrix[90][345] * vector[90] +matrix[91][345] * vector[91] +matrix[92][345] * vector[92] +matrix[93][345] * vector[93] +matrix[94][345] * vector[94] +matrix[95][345] * vector[95] +matrix[96][345] * vector[96] +matrix[97][345] * vector[97] +matrix[98][345] * vector[98] +matrix[99][345] * vector[99] +b[345];
assign result[346] = matrix[0][346] * vector[0] +matrix[1][346] * vector[1] +matrix[2][346] * vector[2] +matrix[3][346] * vector[3] +matrix[4][346] * vector[4] +matrix[5][346] * vector[5] +matrix[6][346] * vector[6] +matrix[7][346] * vector[7] +matrix[8][346] * vector[8] +matrix[9][346] * vector[9] +matrix[10][346] * vector[10] +matrix[11][346] * vector[11] +matrix[12][346] * vector[12] +matrix[13][346] * vector[13] +matrix[14][346] * vector[14] +matrix[15][346] * vector[15] +matrix[16][346] * vector[16] +matrix[17][346] * vector[17] +matrix[18][346] * vector[18] +matrix[19][346] * vector[19] +matrix[20][346] * vector[20] +matrix[21][346] * vector[21] +matrix[22][346] * vector[22] +matrix[23][346] * vector[23] +matrix[24][346] * vector[24] +matrix[25][346] * vector[25] +matrix[26][346] * vector[26] +matrix[27][346] * vector[27] +matrix[28][346] * vector[28] +matrix[29][346] * vector[29] +matrix[30][346] * vector[30] +matrix[31][346] * vector[31] +matrix[32][346] * vector[32] +matrix[33][346] * vector[33] +matrix[34][346] * vector[34] +matrix[35][346] * vector[35] +matrix[36][346] * vector[36] +matrix[37][346] * vector[37] +matrix[38][346] * vector[38] +matrix[39][346] * vector[39] +matrix[40][346] * vector[40] +matrix[41][346] * vector[41] +matrix[42][346] * vector[42] +matrix[43][346] * vector[43] +matrix[44][346] * vector[44] +matrix[45][346] * vector[45] +matrix[46][346] * vector[46] +matrix[47][346] * vector[47] +matrix[48][346] * vector[48] +matrix[49][346] * vector[49] +matrix[50][346] * vector[50] +matrix[51][346] * vector[51] +matrix[52][346] * vector[52] +matrix[53][346] * vector[53] +matrix[54][346] * vector[54] +matrix[55][346] * vector[55] +matrix[56][346] * vector[56] +matrix[57][346] * vector[57] +matrix[58][346] * vector[58] +matrix[59][346] * vector[59] +matrix[60][346] * vector[60] +matrix[61][346] * vector[61] +matrix[62][346] * vector[62] +matrix[63][346] * vector[63] +matrix[64][346] * vector[64] +matrix[65][346] * vector[65] +matrix[66][346] * vector[66] +matrix[67][346] * vector[67] +matrix[68][346] * vector[68] +matrix[69][346] * vector[69] +matrix[70][346] * vector[70] +matrix[71][346] * vector[71] +matrix[72][346] * vector[72] +matrix[73][346] * vector[73] +matrix[74][346] * vector[74] +matrix[75][346] * vector[75] +matrix[76][346] * vector[76] +matrix[77][346] * vector[77] +matrix[78][346] * vector[78] +matrix[79][346] * vector[79] +matrix[80][346] * vector[80] +matrix[81][346] * vector[81] +matrix[82][346] * vector[82] +matrix[83][346] * vector[83] +matrix[84][346] * vector[84] +matrix[85][346] * vector[85] +matrix[86][346] * vector[86] +matrix[87][346] * vector[87] +matrix[88][346] * vector[88] +matrix[89][346] * vector[89] +matrix[90][346] * vector[90] +matrix[91][346] * vector[91] +matrix[92][346] * vector[92] +matrix[93][346] * vector[93] +matrix[94][346] * vector[94] +matrix[95][346] * vector[95] +matrix[96][346] * vector[96] +matrix[97][346] * vector[97] +matrix[98][346] * vector[98] +matrix[99][346] * vector[99] +b[346];
assign result[347] = matrix[0][347] * vector[0] +matrix[1][347] * vector[1] +matrix[2][347] * vector[2] +matrix[3][347] * vector[3] +matrix[4][347] * vector[4] +matrix[5][347] * vector[5] +matrix[6][347] * vector[6] +matrix[7][347] * vector[7] +matrix[8][347] * vector[8] +matrix[9][347] * vector[9] +matrix[10][347] * vector[10] +matrix[11][347] * vector[11] +matrix[12][347] * vector[12] +matrix[13][347] * vector[13] +matrix[14][347] * vector[14] +matrix[15][347] * vector[15] +matrix[16][347] * vector[16] +matrix[17][347] * vector[17] +matrix[18][347] * vector[18] +matrix[19][347] * vector[19] +matrix[20][347] * vector[20] +matrix[21][347] * vector[21] +matrix[22][347] * vector[22] +matrix[23][347] * vector[23] +matrix[24][347] * vector[24] +matrix[25][347] * vector[25] +matrix[26][347] * vector[26] +matrix[27][347] * vector[27] +matrix[28][347] * vector[28] +matrix[29][347] * vector[29] +matrix[30][347] * vector[30] +matrix[31][347] * vector[31] +matrix[32][347] * vector[32] +matrix[33][347] * vector[33] +matrix[34][347] * vector[34] +matrix[35][347] * vector[35] +matrix[36][347] * vector[36] +matrix[37][347] * vector[37] +matrix[38][347] * vector[38] +matrix[39][347] * vector[39] +matrix[40][347] * vector[40] +matrix[41][347] * vector[41] +matrix[42][347] * vector[42] +matrix[43][347] * vector[43] +matrix[44][347] * vector[44] +matrix[45][347] * vector[45] +matrix[46][347] * vector[46] +matrix[47][347] * vector[47] +matrix[48][347] * vector[48] +matrix[49][347] * vector[49] +matrix[50][347] * vector[50] +matrix[51][347] * vector[51] +matrix[52][347] * vector[52] +matrix[53][347] * vector[53] +matrix[54][347] * vector[54] +matrix[55][347] * vector[55] +matrix[56][347] * vector[56] +matrix[57][347] * vector[57] +matrix[58][347] * vector[58] +matrix[59][347] * vector[59] +matrix[60][347] * vector[60] +matrix[61][347] * vector[61] +matrix[62][347] * vector[62] +matrix[63][347] * vector[63] +matrix[64][347] * vector[64] +matrix[65][347] * vector[65] +matrix[66][347] * vector[66] +matrix[67][347] * vector[67] +matrix[68][347] * vector[68] +matrix[69][347] * vector[69] +matrix[70][347] * vector[70] +matrix[71][347] * vector[71] +matrix[72][347] * vector[72] +matrix[73][347] * vector[73] +matrix[74][347] * vector[74] +matrix[75][347] * vector[75] +matrix[76][347] * vector[76] +matrix[77][347] * vector[77] +matrix[78][347] * vector[78] +matrix[79][347] * vector[79] +matrix[80][347] * vector[80] +matrix[81][347] * vector[81] +matrix[82][347] * vector[82] +matrix[83][347] * vector[83] +matrix[84][347] * vector[84] +matrix[85][347] * vector[85] +matrix[86][347] * vector[86] +matrix[87][347] * vector[87] +matrix[88][347] * vector[88] +matrix[89][347] * vector[89] +matrix[90][347] * vector[90] +matrix[91][347] * vector[91] +matrix[92][347] * vector[92] +matrix[93][347] * vector[93] +matrix[94][347] * vector[94] +matrix[95][347] * vector[95] +matrix[96][347] * vector[96] +matrix[97][347] * vector[97] +matrix[98][347] * vector[98] +matrix[99][347] * vector[99] +b[347];
assign result[348] = matrix[0][348] * vector[0] +matrix[1][348] * vector[1] +matrix[2][348] * vector[2] +matrix[3][348] * vector[3] +matrix[4][348] * vector[4] +matrix[5][348] * vector[5] +matrix[6][348] * vector[6] +matrix[7][348] * vector[7] +matrix[8][348] * vector[8] +matrix[9][348] * vector[9] +matrix[10][348] * vector[10] +matrix[11][348] * vector[11] +matrix[12][348] * vector[12] +matrix[13][348] * vector[13] +matrix[14][348] * vector[14] +matrix[15][348] * vector[15] +matrix[16][348] * vector[16] +matrix[17][348] * vector[17] +matrix[18][348] * vector[18] +matrix[19][348] * vector[19] +matrix[20][348] * vector[20] +matrix[21][348] * vector[21] +matrix[22][348] * vector[22] +matrix[23][348] * vector[23] +matrix[24][348] * vector[24] +matrix[25][348] * vector[25] +matrix[26][348] * vector[26] +matrix[27][348] * vector[27] +matrix[28][348] * vector[28] +matrix[29][348] * vector[29] +matrix[30][348] * vector[30] +matrix[31][348] * vector[31] +matrix[32][348] * vector[32] +matrix[33][348] * vector[33] +matrix[34][348] * vector[34] +matrix[35][348] * vector[35] +matrix[36][348] * vector[36] +matrix[37][348] * vector[37] +matrix[38][348] * vector[38] +matrix[39][348] * vector[39] +matrix[40][348] * vector[40] +matrix[41][348] * vector[41] +matrix[42][348] * vector[42] +matrix[43][348] * vector[43] +matrix[44][348] * vector[44] +matrix[45][348] * vector[45] +matrix[46][348] * vector[46] +matrix[47][348] * vector[47] +matrix[48][348] * vector[48] +matrix[49][348] * vector[49] +matrix[50][348] * vector[50] +matrix[51][348] * vector[51] +matrix[52][348] * vector[52] +matrix[53][348] * vector[53] +matrix[54][348] * vector[54] +matrix[55][348] * vector[55] +matrix[56][348] * vector[56] +matrix[57][348] * vector[57] +matrix[58][348] * vector[58] +matrix[59][348] * vector[59] +matrix[60][348] * vector[60] +matrix[61][348] * vector[61] +matrix[62][348] * vector[62] +matrix[63][348] * vector[63] +matrix[64][348] * vector[64] +matrix[65][348] * vector[65] +matrix[66][348] * vector[66] +matrix[67][348] * vector[67] +matrix[68][348] * vector[68] +matrix[69][348] * vector[69] +matrix[70][348] * vector[70] +matrix[71][348] * vector[71] +matrix[72][348] * vector[72] +matrix[73][348] * vector[73] +matrix[74][348] * vector[74] +matrix[75][348] * vector[75] +matrix[76][348] * vector[76] +matrix[77][348] * vector[77] +matrix[78][348] * vector[78] +matrix[79][348] * vector[79] +matrix[80][348] * vector[80] +matrix[81][348] * vector[81] +matrix[82][348] * vector[82] +matrix[83][348] * vector[83] +matrix[84][348] * vector[84] +matrix[85][348] * vector[85] +matrix[86][348] * vector[86] +matrix[87][348] * vector[87] +matrix[88][348] * vector[88] +matrix[89][348] * vector[89] +matrix[90][348] * vector[90] +matrix[91][348] * vector[91] +matrix[92][348] * vector[92] +matrix[93][348] * vector[93] +matrix[94][348] * vector[94] +matrix[95][348] * vector[95] +matrix[96][348] * vector[96] +matrix[97][348] * vector[97] +matrix[98][348] * vector[98] +matrix[99][348] * vector[99] +b[348];
assign result[349] = matrix[0][349] * vector[0] +matrix[1][349] * vector[1] +matrix[2][349] * vector[2] +matrix[3][349] * vector[3] +matrix[4][349] * vector[4] +matrix[5][349] * vector[5] +matrix[6][349] * vector[6] +matrix[7][349] * vector[7] +matrix[8][349] * vector[8] +matrix[9][349] * vector[9] +matrix[10][349] * vector[10] +matrix[11][349] * vector[11] +matrix[12][349] * vector[12] +matrix[13][349] * vector[13] +matrix[14][349] * vector[14] +matrix[15][349] * vector[15] +matrix[16][349] * vector[16] +matrix[17][349] * vector[17] +matrix[18][349] * vector[18] +matrix[19][349] * vector[19] +matrix[20][349] * vector[20] +matrix[21][349] * vector[21] +matrix[22][349] * vector[22] +matrix[23][349] * vector[23] +matrix[24][349] * vector[24] +matrix[25][349] * vector[25] +matrix[26][349] * vector[26] +matrix[27][349] * vector[27] +matrix[28][349] * vector[28] +matrix[29][349] * vector[29] +matrix[30][349] * vector[30] +matrix[31][349] * vector[31] +matrix[32][349] * vector[32] +matrix[33][349] * vector[33] +matrix[34][349] * vector[34] +matrix[35][349] * vector[35] +matrix[36][349] * vector[36] +matrix[37][349] * vector[37] +matrix[38][349] * vector[38] +matrix[39][349] * vector[39] +matrix[40][349] * vector[40] +matrix[41][349] * vector[41] +matrix[42][349] * vector[42] +matrix[43][349] * vector[43] +matrix[44][349] * vector[44] +matrix[45][349] * vector[45] +matrix[46][349] * vector[46] +matrix[47][349] * vector[47] +matrix[48][349] * vector[48] +matrix[49][349] * vector[49] +matrix[50][349] * vector[50] +matrix[51][349] * vector[51] +matrix[52][349] * vector[52] +matrix[53][349] * vector[53] +matrix[54][349] * vector[54] +matrix[55][349] * vector[55] +matrix[56][349] * vector[56] +matrix[57][349] * vector[57] +matrix[58][349] * vector[58] +matrix[59][349] * vector[59] +matrix[60][349] * vector[60] +matrix[61][349] * vector[61] +matrix[62][349] * vector[62] +matrix[63][349] * vector[63] +matrix[64][349] * vector[64] +matrix[65][349] * vector[65] +matrix[66][349] * vector[66] +matrix[67][349] * vector[67] +matrix[68][349] * vector[68] +matrix[69][349] * vector[69] +matrix[70][349] * vector[70] +matrix[71][349] * vector[71] +matrix[72][349] * vector[72] +matrix[73][349] * vector[73] +matrix[74][349] * vector[74] +matrix[75][349] * vector[75] +matrix[76][349] * vector[76] +matrix[77][349] * vector[77] +matrix[78][349] * vector[78] +matrix[79][349] * vector[79] +matrix[80][349] * vector[80] +matrix[81][349] * vector[81] +matrix[82][349] * vector[82] +matrix[83][349] * vector[83] +matrix[84][349] * vector[84] +matrix[85][349] * vector[85] +matrix[86][349] * vector[86] +matrix[87][349] * vector[87] +matrix[88][349] * vector[88] +matrix[89][349] * vector[89] +matrix[90][349] * vector[90] +matrix[91][349] * vector[91] +matrix[92][349] * vector[92] +matrix[93][349] * vector[93] +matrix[94][349] * vector[94] +matrix[95][349] * vector[95] +matrix[96][349] * vector[96] +matrix[97][349] * vector[97] +matrix[98][349] * vector[98] +matrix[99][349] * vector[99] +b[349];
assign result[350] = matrix[0][350] * vector[0] +matrix[1][350] * vector[1] +matrix[2][350] * vector[2] +matrix[3][350] * vector[3] +matrix[4][350] * vector[4] +matrix[5][350] * vector[5] +matrix[6][350] * vector[6] +matrix[7][350] * vector[7] +matrix[8][350] * vector[8] +matrix[9][350] * vector[9] +matrix[10][350] * vector[10] +matrix[11][350] * vector[11] +matrix[12][350] * vector[12] +matrix[13][350] * vector[13] +matrix[14][350] * vector[14] +matrix[15][350] * vector[15] +matrix[16][350] * vector[16] +matrix[17][350] * vector[17] +matrix[18][350] * vector[18] +matrix[19][350] * vector[19] +matrix[20][350] * vector[20] +matrix[21][350] * vector[21] +matrix[22][350] * vector[22] +matrix[23][350] * vector[23] +matrix[24][350] * vector[24] +matrix[25][350] * vector[25] +matrix[26][350] * vector[26] +matrix[27][350] * vector[27] +matrix[28][350] * vector[28] +matrix[29][350] * vector[29] +matrix[30][350] * vector[30] +matrix[31][350] * vector[31] +matrix[32][350] * vector[32] +matrix[33][350] * vector[33] +matrix[34][350] * vector[34] +matrix[35][350] * vector[35] +matrix[36][350] * vector[36] +matrix[37][350] * vector[37] +matrix[38][350] * vector[38] +matrix[39][350] * vector[39] +matrix[40][350] * vector[40] +matrix[41][350] * vector[41] +matrix[42][350] * vector[42] +matrix[43][350] * vector[43] +matrix[44][350] * vector[44] +matrix[45][350] * vector[45] +matrix[46][350] * vector[46] +matrix[47][350] * vector[47] +matrix[48][350] * vector[48] +matrix[49][350] * vector[49] +matrix[50][350] * vector[50] +matrix[51][350] * vector[51] +matrix[52][350] * vector[52] +matrix[53][350] * vector[53] +matrix[54][350] * vector[54] +matrix[55][350] * vector[55] +matrix[56][350] * vector[56] +matrix[57][350] * vector[57] +matrix[58][350] * vector[58] +matrix[59][350] * vector[59] +matrix[60][350] * vector[60] +matrix[61][350] * vector[61] +matrix[62][350] * vector[62] +matrix[63][350] * vector[63] +matrix[64][350] * vector[64] +matrix[65][350] * vector[65] +matrix[66][350] * vector[66] +matrix[67][350] * vector[67] +matrix[68][350] * vector[68] +matrix[69][350] * vector[69] +matrix[70][350] * vector[70] +matrix[71][350] * vector[71] +matrix[72][350] * vector[72] +matrix[73][350] * vector[73] +matrix[74][350] * vector[74] +matrix[75][350] * vector[75] +matrix[76][350] * vector[76] +matrix[77][350] * vector[77] +matrix[78][350] * vector[78] +matrix[79][350] * vector[79] +matrix[80][350] * vector[80] +matrix[81][350] * vector[81] +matrix[82][350] * vector[82] +matrix[83][350] * vector[83] +matrix[84][350] * vector[84] +matrix[85][350] * vector[85] +matrix[86][350] * vector[86] +matrix[87][350] * vector[87] +matrix[88][350] * vector[88] +matrix[89][350] * vector[89] +matrix[90][350] * vector[90] +matrix[91][350] * vector[91] +matrix[92][350] * vector[92] +matrix[93][350] * vector[93] +matrix[94][350] * vector[94] +matrix[95][350] * vector[95] +matrix[96][350] * vector[96] +matrix[97][350] * vector[97] +matrix[98][350] * vector[98] +matrix[99][350] * vector[99] +b[350];
assign result[351] = matrix[0][351] * vector[0] +matrix[1][351] * vector[1] +matrix[2][351] * vector[2] +matrix[3][351] * vector[3] +matrix[4][351] * vector[4] +matrix[5][351] * vector[5] +matrix[6][351] * vector[6] +matrix[7][351] * vector[7] +matrix[8][351] * vector[8] +matrix[9][351] * vector[9] +matrix[10][351] * vector[10] +matrix[11][351] * vector[11] +matrix[12][351] * vector[12] +matrix[13][351] * vector[13] +matrix[14][351] * vector[14] +matrix[15][351] * vector[15] +matrix[16][351] * vector[16] +matrix[17][351] * vector[17] +matrix[18][351] * vector[18] +matrix[19][351] * vector[19] +matrix[20][351] * vector[20] +matrix[21][351] * vector[21] +matrix[22][351] * vector[22] +matrix[23][351] * vector[23] +matrix[24][351] * vector[24] +matrix[25][351] * vector[25] +matrix[26][351] * vector[26] +matrix[27][351] * vector[27] +matrix[28][351] * vector[28] +matrix[29][351] * vector[29] +matrix[30][351] * vector[30] +matrix[31][351] * vector[31] +matrix[32][351] * vector[32] +matrix[33][351] * vector[33] +matrix[34][351] * vector[34] +matrix[35][351] * vector[35] +matrix[36][351] * vector[36] +matrix[37][351] * vector[37] +matrix[38][351] * vector[38] +matrix[39][351] * vector[39] +matrix[40][351] * vector[40] +matrix[41][351] * vector[41] +matrix[42][351] * vector[42] +matrix[43][351] * vector[43] +matrix[44][351] * vector[44] +matrix[45][351] * vector[45] +matrix[46][351] * vector[46] +matrix[47][351] * vector[47] +matrix[48][351] * vector[48] +matrix[49][351] * vector[49] +matrix[50][351] * vector[50] +matrix[51][351] * vector[51] +matrix[52][351] * vector[52] +matrix[53][351] * vector[53] +matrix[54][351] * vector[54] +matrix[55][351] * vector[55] +matrix[56][351] * vector[56] +matrix[57][351] * vector[57] +matrix[58][351] * vector[58] +matrix[59][351] * vector[59] +matrix[60][351] * vector[60] +matrix[61][351] * vector[61] +matrix[62][351] * vector[62] +matrix[63][351] * vector[63] +matrix[64][351] * vector[64] +matrix[65][351] * vector[65] +matrix[66][351] * vector[66] +matrix[67][351] * vector[67] +matrix[68][351] * vector[68] +matrix[69][351] * vector[69] +matrix[70][351] * vector[70] +matrix[71][351] * vector[71] +matrix[72][351] * vector[72] +matrix[73][351] * vector[73] +matrix[74][351] * vector[74] +matrix[75][351] * vector[75] +matrix[76][351] * vector[76] +matrix[77][351] * vector[77] +matrix[78][351] * vector[78] +matrix[79][351] * vector[79] +matrix[80][351] * vector[80] +matrix[81][351] * vector[81] +matrix[82][351] * vector[82] +matrix[83][351] * vector[83] +matrix[84][351] * vector[84] +matrix[85][351] * vector[85] +matrix[86][351] * vector[86] +matrix[87][351] * vector[87] +matrix[88][351] * vector[88] +matrix[89][351] * vector[89] +matrix[90][351] * vector[90] +matrix[91][351] * vector[91] +matrix[92][351] * vector[92] +matrix[93][351] * vector[93] +matrix[94][351] * vector[94] +matrix[95][351] * vector[95] +matrix[96][351] * vector[96] +matrix[97][351] * vector[97] +matrix[98][351] * vector[98] +matrix[99][351] * vector[99] +b[351];
assign result[352] = matrix[0][352] * vector[0] +matrix[1][352] * vector[1] +matrix[2][352] * vector[2] +matrix[3][352] * vector[3] +matrix[4][352] * vector[4] +matrix[5][352] * vector[5] +matrix[6][352] * vector[6] +matrix[7][352] * vector[7] +matrix[8][352] * vector[8] +matrix[9][352] * vector[9] +matrix[10][352] * vector[10] +matrix[11][352] * vector[11] +matrix[12][352] * vector[12] +matrix[13][352] * vector[13] +matrix[14][352] * vector[14] +matrix[15][352] * vector[15] +matrix[16][352] * vector[16] +matrix[17][352] * vector[17] +matrix[18][352] * vector[18] +matrix[19][352] * vector[19] +matrix[20][352] * vector[20] +matrix[21][352] * vector[21] +matrix[22][352] * vector[22] +matrix[23][352] * vector[23] +matrix[24][352] * vector[24] +matrix[25][352] * vector[25] +matrix[26][352] * vector[26] +matrix[27][352] * vector[27] +matrix[28][352] * vector[28] +matrix[29][352] * vector[29] +matrix[30][352] * vector[30] +matrix[31][352] * vector[31] +matrix[32][352] * vector[32] +matrix[33][352] * vector[33] +matrix[34][352] * vector[34] +matrix[35][352] * vector[35] +matrix[36][352] * vector[36] +matrix[37][352] * vector[37] +matrix[38][352] * vector[38] +matrix[39][352] * vector[39] +matrix[40][352] * vector[40] +matrix[41][352] * vector[41] +matrix[42][352] * vector[42] +matrix[43][352] * vector[43] +matrix[44][352] * vector[44] +matrix[45][352] * vector[45] +matrix[46][352] * vector[46] +matrix[47][352] * vector[47] +matrix[48][352] * vector[48] +matrix[49][352] * vector[49] +matrix[50][352] * vector[50] +matrix[51][352] * vector[51] +matrix[52][352] * vector[52] +matrix[53][352] * vector[53] +matrix[54][352] * vector[54] +matrix[55][352] * vector[55] +matrix[56][352] * vector[56] +matrix[57][352] * vector[57] +matrix[58][352] * vector[58] +matrix[59][352] * vector[59] +matrix[60][352] * vector[60] +matrix[61][352] * vector[61] +matrix[62][352] * vector[62] +matrix[63][352] * vector[63] +matrix[64][352] * vector[64] +matrix[65][352] * vector[65] +matrix[66][352] * vector[66] +matrix[67][352] * vector[67] +matrix[68][352] * vector[68] +matrix[69][352] * vector[69] +matrix[70][352] * vector[70] +matrix[71][352] * vector[71] +matrix[72][352] * vector[72] +matrix[73][352] * vector[73] +matrix[74][352] * vector[74] +matrix[75][352] * vector[75] +matrix[76][352] * vector[76] +matrix[77][352] * vector[77] +matrix[78][352] * vector[78] +matrix[79][352] * vector[79] +matrix[80][352] * vector[80] +matrix[81][352] * vector[81] +matrix[82][352] * vector[82] +matrix[83][352] * vector[83] +matrix[84][352] * vector[84] +matrix[85][352] * vector[85] +matrix[86][352] * vector[86] +matrix[87][352] * vector[87] +matrix[88][352] * vector[88] +matrix[89][352] * vector[89] +matrix[90][352] * vector[90] +matrix[91][352] * vector[91] +matrix[92][352] * vector[92] +matrix[93][352] * vector[93] +matrix[94][352] * vector[94] +matrix[95][352] * vector[95] +matrix[96][352] * vector[96] +matrix[97][352] * vector[97] +matrix[98][352] * vector[98] +matrix[99][352] * vector[99] +b[352];
assign result[353] = matrix[0][353] * vector[0] +matrix[1][353] * vector[1] +matrix[2][353] * vector[2] +matrix[3][353] * vector[3] +matrix[4][353] * vector[4] +matrix[5][353] * vector[5] +matrix[6][353] * vector[6] +matrix[7][353] * vector[7] +matrix[8][353] * vector[8] +matrix[9][353] * vector[9] +matrix[10][353] * vector[10] +matrix[11][353] * vector[11] +matrix[12][353] * vector[12] +matrix[13][353] * vector[13] +matrix[14][353] * vector[14] +matrix[15][353] * vector[15] +matrix[16][353] * vector[16] +matrix[17][353] * vector[17] +matrix[18][353] * vector[18] +matrix[19][353] * vector[19] +matrix[20][353] * vector[20] +matrix[21][353] * vector[21] +matrix[22][353] * vector[22] +matrix[23][353] * vector[23] +matrix[24][353] * vector[24] +matrix[25][353] * vector[25] +matrix[26][353] * vector[26] +matrix[27][353] * vector[27] +matrix[28][353] * vector[28] +matrix[29][353] * vector[29] +matrix[30][353] * vector[30] +matrix[31][353] * vector[31] +matrix[32][353] * vector[32] +matrix[33][353] * vector[33] +matrix[34][353] * vector[34] +matrix[35][353] * vector[35] +matrix[36][353] * vector[36] +matrix[37][353] * vector[37] +matrix[38][353] * vector[38] +matrix[39][353] * vector[39] +matrix[40][353] * vector[40] +matrix[41][353] * vector[41] +matrix[42][353] * vector[42] +matrix[43][353] * vector[43] +matrix[44][353] * vector[44] +matrix[45][353] * vector[45] +matrix[46][353] * vector[46] +matrix[47][353] * vector[47] +matrix[48][353] * vector[48] +matrix[49][353] * vector[49] +matrix[50][353] * vector[50] +matrix[51][353] * vector[51] +matrix[52][353] * vector[52] +matrix[53][353] * vector[53] +matrix[54][353] * vector[54] +matrix[55][353] * vector[55] +matrix[56][353] * vector[56] +matrix[57][353] * vector[57] +matrix[58][353] * vector[58] +matrix[59][353] * vector[59] +matrix[60][353] * vector[60] +matrix[61][353] * vector[61] +matrix[62][353] * vector[62] +matrix[63][353] * vector[63] +matrix[64][353] * vector[64] +matrix[65][353] * vector[65] +matrix[66][353] * vector[66] +matrix[67][353] * vector[67] +matrix[68][353] * vector[68] +matrix[69][353] * vector[69] +matrix[70][353] * vector[70] +matrix[71][353] * vector[71] +matrix[72][353] * vector[72] +matrix[73][353] * vector[73] +matrix[74][353] * vector[74] +matrix[75][353] * vector[75] +matrix[76][353] * vector[76] +matrix[77][353] * vector[77] +matrix[78][353] * vector[78] +matrix[79][353] * vector[79] +matrix[80][353] * vector[80] +matrix[81][353] * vector[81] +matrix[82][353] * vector[82] +matrix[83][353] * vector[83] +matrix[84][353] * vector[84] +matrix[85][353] * vector[85] +matrix[86][353] * vector[86] +matrix[87][353] * vector[87] +matrix[88][353] * vector[88] +matrix[89][353] * vector[89] +matrix[90][353] * vector[90] +matrix[91][353] * vector[91] +matrix[92][353] * vector[92] +matrix[93][353] * vector[93] +matrix[94][353] * vector[94] +matrix[95][353] * vector[95] +matrix[96][353] * vector[96] +matrix[97][353] * vector[97] +matrix[98][353] * vector[98] +matrix[99][353] * vector[99] +b[353];
assign result[354] = matrix[0][354] * vector[0] +matrix[1][354] * vector[1] +matrix[2][354] * vector[2] +matrix[3][354] * vector[3] +matrix[4][354] * vector[4] +matrix[5][354] * vector[5] +matrix[6][354] * vector[6] +matrix[7][354] * vector[7] +matrix[8][354] * vector[8] +matrix[9][354] * vector[9] +matrix[10][354] * vector[10] +matrix[11][354] * vector[11] +matrix[12][354] * vector[12] +matrix[13][354] * vector[13] +matrix[14][354] * vector[14] +matrix[15][354] * vector[15] +matrix[16][354] * vector[16] +matrix[17][354] * vector[17] +matrix[18][354] * vector[18] +matrix[19][354] * vector[19] +matrix[20][354] * vector[20] +matrix[21][354] * vector[21] +matrix[22][354] * vector[22] +matrix[23][354] * vector[23] +matrix[24][354] * vector[24] +matrix[25][354] * vector[25] +matrix[26][354] * vector[26] +matrix[27][354] * vector[27] +matrix[28][354] * vector[28] +matrix[29][354] * vector[29] +matrix[30][354] * vector[30] +matrix[31][354] * vector[31] +matrix[32][354] * vector[32] +matrix[33][354] * vector[33] +matrix[34][354] * vector[34] +matrix[35][354] * vector[35] +matrix[36][354] * vector[36] +matrix[37][354] * vector[37] +matrix[38][354] * vector[38] +matrix[39][354] * vector[39] +matrix[40][354] * vector[40] +matrix[41][354] * vector[41] +matrix[42][354] * vector[42] +matrix[43][354] * vector[43] +matrix[44][354] * vector[44] +matrix[45][354] * vector[45] +matrix[46][354] * vector[46] +matrix[47][354] * vector[47] +matrix[48][354] * vector[48] +matrix[49][354] * vector[49] +matrix[50][354] * vector[50] +matrix[51][354] * vector[51] +matrix[52][354] * vector[52] +matrix[53][354] * vector[53] +matrix[54][354] * vector[54] +matrix[55][354] * vector[55] +matrix[56][354] * vector[56] +matrix[57][354] * vector[57] +matrix[58][354] * vector[58] +matrix[59][354] * vector[59] +matrix[60][354] * vector[60] +matrix[61][354] * vector[61] +matrix[62][354] * vector[62] +matrix[63][354] * vector[63] +matrix[64][354] * vector[64] +matrix[65][354] * vector[65] +matrix[66][354] * vector[66] +matrix[67][354] * vector[67] +matrix[68][354] * vector[68] +matrix[69][354] * vector[69] +matrix[70][354] * vector[70] +matrix[71][354] * vector[71] +matrix[72][354] * vector[72] +matrix[73][354] * vector[73] +matrix[74][354] * vector[74] +matrix[75][354] * vector[75] +matrix[76][354] * vector[76] +matrix[77][354] * vector[77] +matrix[78][354] * vector[78] +matrix[79][354] * vector[79] +matrix[80][354] * vector[80] +matrix[81][354] * vector[81] +matrix[82][354] * vector[82] +matrix[83][354] * vector[83] +matrix[84][354] * vector[84] +matrix[85][354] * vector[85] +matrix[86][354] * vector[86] +matrix[87][354] * vector[87] +matrix[88][354] * vector[88] +matrix[89][354] * vector[89] +matrix[90][354] * vector[90] +matrix[91][354] * vector[91] +matrix[92][354] * vector[92] +matrix[93][354] * vector[93] +matrix[94][354] * vector[94] +matrix[95][354] * vector[95] +matrix[96][354] * vector[96] +matrix[97][354] * vector[97] +matrix[98][354] * vector[98] +matrix[99][354] * vector[99] +b[354];
assign result[355] = matrix[0][355] * vector[0] +matrix[1][355] * vector[1] +matrix[2][355] * vector[2] +matrix[3][355] * vector[3] +matrix[4][355] * vector[4] +matrix[5][355] * vector[5] +matrix[6][355] * vector[6] +matrix[7][355] * vector[7] +matrix[8][355] * vector[8] +matrix[9][355] * vector[9] +matrix[10][355] * vector[10] +matrix[11][355] * vector[11] +matrix[12][355] * vector[12] +matrix[13][355] * vector[13] +matrix[14][355] * vector[14] +matrix[15][355] * vector[15] +matrix[16][355] * vector[16] +matrix[17][355] * vector[17] +matrix[18][355] * vector[18] +matrix[19][355] * vector[19] +matrix[20][355] * vector[20] +matrix[21][355] * vector[21] +matrix[22][355] * vector[22] +matrix[23][355] * vector[23] +matrix[24][355] * vector[24] +matrix[25][355] * vector[25] +matrix[26][355] * vector[26] +matrix[27][355] * vector[27] +matrix[28][355] * vector[28] +matrix[29][355] * vector[29] +matrix[30][355] * vector[30] +matrix[31][355] * vector[31] +matrix[32][355] * vector[32] +matrix[33][355] * vector[33] +matrix[34][355] * vector[34] +matrix[35][355] * vector[35] +matrix[36][355] * vector[36] +matrix[37][355] * vector[37] +matrix[38][355] * vector[38] +matrix[39][355] * vector[39] +matrix[40][355] * vector[40] +matrix[41][355] * vector[41] +matrix[42][355] * vector[42] +matrix[43][355] * vector[43] +matrix[44][355] * vector[44] +matrix[45][355] * vector[45] +matrix[46][355] * vector[46] +matrix[47][355] * vector[47] +matrix[48][355] * vector[48] +matrix[49][355] * vector[49] +matrix[50][355] * vector[50] +matrix[51][355] * vector[51] +matrix[52][355] * vector[52] +matrix[53][355] * vector[53] +matrix[54][355] * vector[54] +matrix[55][355] * vector[55] +matrix[56][355] * vector[56] +matrix[57][355] * vector[57] +matrix[58][355] * vector[58] +matrix[59][355] * vector[59] +matrix[60][355] * vector[60] +matrix[61][355] * vector[61] +matrix[62][355] * vector[62] +matrix[63][355] * vector[63] +matrix[64][355] * vector[64] +matrix[65][355] * vector[65] +matrix[66][355] * vector[66] +matrix[67][355] * vector[67] +matrix[68][355] * vector[68] +matrix[69][355] * vector[69] +matrix[70][355] * vector[70] +matrix[71][355] * vector[71] +matrix[72][355] * vector[72] +matrix[73][355] * vector[73] +matrix[74][355] * vector[74] +matrix[75][355] * vector[75] +matrix[76][355] * vector[76] +matrix[77][355] * vector[77] +matrix[78][355] * vector[78] +matrix[79][355] * vector[79] +matrix[80][355] * vector[80] +matrix[81][355] * vector[81] +matrix[82][355] * vector[82] +matrix[83][355] * vector[83] +matrix[84][355] * vector[84] +matrix[85][355] * vector[85] +matrix[86][355] * vector[86] +matrix[87][355] * vector[87] +matrix[88][355] * vector[88] +matrix[89][355] * vector[89] +matrix[90][355] * vector[90] +matrix[91][355] * vector[91] +matrix[92][355] * vector[92] +matrix[93][355] * vector[93] +matrix[94][355] * vector[94] +matrix[95][355] * vector[95] +matrix[96][355] * vector[96] +matrix[97][355] * vector[97] +matrix[98][355] * vector[98] +matrix[99][355] * vector[99] +b[355];
assign result[356] = matrix[0][356] * vector[0] +matrix[1][356] * vector[1] +matrix[2][356] * vector[2] +matrix[3][356] * vector[3] +matrix[4][356] * vector[4] +matrix[5][356] * vector[5] +matrix[6][356] * vector[6] +matrix[7][356] * vector[7] +matrix[8][356] * vector[8] +matrix[9][356] * vector[9] +matrix[10][356] * vector[10] +matrix[11][356] * vector[11] +matrix[12][356] * vector[12] +matrix[13][356] * vector[13] +matrix[14][356] * vector[14] +matrix[15][356] * vector[15] +matrix[16][356] * vector[16] +matrix[17][356] * vector[17] +matrix[18][356] * vector[18] +matrix[19][356] * vector[19] +matrix[20][356] * vector[20] +matrix[21][356] * vector[21] +matrix[22][356] * vector[22] +matrix[23][356] * vector[23] +matrix[24][356] * vector[24] +matrix[25][356] * vector[25] +matrix[26][356] * vector[26] +matrix[27][356] * vector[27] +matrix[28][356] * vector[28] +matrix[29][356] * vector[29] +matrix[30][356] * vector[30] +matrix[31][356] * vector[31] +matrix[32][356] * vector[32] +matrix[33][356] * vector[33] +matrix[34][356] * vector[34] +matrix[35][356] * vector[35] +matrix[36][356] * vector[36] +matrix[37][356] * vector[37] +matrix[38][356] * vector[38] +matrix[39][356] * vector[39] +matrix[40][356] * vector[40] +matrix[41][356] * vector[41] +matrix[42][356] * vector[42] +matrix[43][356] * vector[43] +matrix[44][356] * vector[44] +matrix[45][356] * vector[45] +matrix[46][356] * vector[46] +matrix[47][356] * vector[47] +matrix[48][356] * vector[48] +matrix[49][356] * vector[49] +matrix[50][356] * vector[50] +matrix[51][356] * vector[51] +matrix[52][356] * vector[52] +matrix[53][356] * vector[53] +matrix[54][356] * vector[54] +matrix[55][356] * vector[55] +matrix[56][356] * vector[56] +matrix[57][356] * vector[57] +matrix[58][356] * vector[58] +matrix[59][356] * vector[59] +matrix[60][356] * vector[60] +matrix[61][356] * vector[61] +matrix[62][356] * vector[62] +matrix[63][356] * vector[63] +matrix[64][356] * vector[64] +matrix[65][356] * vector[65] +matrix[66][356] * vector[66] +matrix[67][356] * vector[67] +matrix[68][356] * vector[68] +matrix[69][356] * vector[69] +matrix[70][356] * vector[70] +matrix[71][356] * vector[71] +matrix[72][356] * vector[72] +matrix[73][356] * vector[73] +matrix[74][356] * vector[74] +matrix[75][356] * vector[75] +matrix[76][356] * vector[76] +matrix[77][356] * vector[77] +matrix[78][356] * vector[78] +matrix[79][356] * vector[79] +matrix[80][356] * vector[80] +matrix[81][356] * vector[81] +matrix[82][356] * vector[82] +matrix[83][356] * vector[83] +matrix[84][356] * vector[84] +matrix[85][356] * vector[85] +matrix[86][356] * vector[86] +matrix[87][356] * vector[87] +matrix[88][356] * vector[88] +matrix[89][356] * vector[89] +matrix[90][356] * vector[90] +matrix[91][356] * vector[91] +matrix[92][356] * vector[92] +matrix[93][356] * vector[93] +matrix[94][356] * vector[94] +matrix[95][356] * vector[95] +matrix[96][356] * vector[96] +matrix[97][356] * vector[97] +matrix[98][356] * vector[98] +matrix[99][356] * vector[99] +b[356];
assign result[357] = matrix[0][357] * vector[0] +matrix[1][357] * vector[1] +matrix[2][357] * vector[2] +matrix[3][357] * vector[3] +matrix[4][357] * vector[4] +matrix[5][357] * vector[5] +matrix[6][357] * vector[6] +matrix[7][357] * vector[7] +matrix[8][357] * vector[8] +matrix[9][357] * vector[9] +matrix[10][357] * vector[10] +matrix[11][357] * vector[11] +matrix[12][357] * vector[12] +matrix[13][357] * vector[13] +matrix[14][357] * vector[14] +matrix[15][357] * vector[15] +matrix[16][357] * vector[16] +matrix[17][357] * vector[17] +matrix[18][357] * vector[18] +matrix[19][357] * vector[19] +matrix[20][357] * vector[20] +matrix[21][357] * vector[21] +matrix[22][357] * vector[22] +matrix[23][357] * vector[23] +matrix[24][357] * vector[24] +matrix[25][357] * vector[25] +matrix[26][357] * vector[26] +matrix[27][357] * vector[27] +matrix[28][357] * vector[28] +matrix[29][357] * vector[29] +matrix[30][357] * vector[30] +matrix[31][357] * vector[31] +matrix[32][357] * vector[32] +matrix[33][357] * vector[33] +matrix[34][357] * vector[34] +matrix[35][357] * vector[35] +matrix[36][357] * vector[36] +matrix[37][357] * vector[37] +matrix[38][357] * vector[38] +matrix[39][357] * vector[39] +matrix[40][357] * vector[40] +matrix[41][357] * vector[41] +matrix[42][357] * vector[42] +matrix[43][357] * vector[43] +matrix[44][357] * vector[44] +matrix[45][357] * vector[45] +matrix[46][357] * vector[46] +matrix[47][357] * vector[47] +matrix[48][357] * vector[48] +matrix[49][357] * vector[49] +matrix[50][357] * vector[50] +matrix[51][357] * vector[51] +matrix[52][357] * vector[52] +matrix[53][357] * vector[53] +matrix[54][357] * vector[54] +matrix[55][357] * vector[55] +matrix[56][357] * vector[56] +matrix[57][357] * vector[57] +matrix[58][357] * vector[58] +matrix[59][357] * vector[59] +matrix[60][357] * vector[60] +matrix[61][357] * vector[61] +matrix[62][357] * vector[62] +matrix[63][357] * vector[63] +matrix[64][357] * vector[64] +matrix[65][357] * vector[65] +matrix[66][357] * vector[66] +matrix[67][357] * vector[67] +matrix[68][357] * vector[68] +matrix[69][357] * vector[69] +matrix[70][357] * vector[70] +matrix[71][357] * vector[71] +matrix[72][357] * vector[72] +matrix[73][357] * vector[73] +matrix[74][357] * vector[74] +matrix[75][357] * vector[75] +matrix[76][357] * vector[76] +matrix[77][357] * vector[77] +matrix[78][357] * vector[78] +matrix[79][357] * vector[79] +matrix[80][357] * vector[80] +matrix[81][357] * vector[81] +matrix[82][357] * vector[82] +matrix[83][357] * vector[83] +matrix[84][357] * vector[84] +matrix[85][357] * vector[85] +matrix[86][357] * vector[86] +matrix[87][357] * vector[87] +matrix[88][357] * vector[88] +matrix[89][357] * vector[89] +matrix[90][357] * vector[90] +matrix[91][357] * vector[91] +matrix[92][357] * vector[92] +matrix[93][357] * vector[93] +matrix[94][357] * vector[94] +matrix[95][357] * vector[95] +matrix[96][357] * vector[96] +matrix[97][357] * vector[97] +matrix[98][357] * vector[98] +matrix[99][357] * vector[99] +b[357];
assign result[358] = matrix[0][358] * vector[0] +matrix[1][358] * vector[1] +matrix[2][358] * vector[2] +matrix[3][358] * vector[3] +matrix[4][358] * vector[4] +matrix[5][358] * vector[5] +matrix[6][358] * vector[6] +matrix[7][358] * vector[7] +matrix[8][358] * vector[8] +matrix[9][358] * vector[9] +matrix[10][358] * vector[10] +matrix[11][358] * vector[11] +matrix[12][358] * vector[12] +matrix[13][358] * vector[13] +matrix[14][358] * vector[14] +matrix[15][358] * vector[15] +matrix[16][358] * vector[16] +matrix[17][358] * vector[17] +matrix[18][358] * vector[18] +matrix[19][358] * vector[19] +matrix[20][358] * vector[20] +matrix[21][358] * vector[21] +matrix[22][358] * vector[22] +matrix[23][358] * vector[23] +matrix[24][358] * vector[24] +matrix[25][358] * vector[25] +matrix[26][358] * vector[26] +matrix[27][358] * vector[27] +matrix[28][358] * vector[28] +matrix[29][358] * vector[29] +matrix[30][358] * vector[30] +matrix[31][358] * vector[31] +matrix[32][358] * vector[32] +matrix[33][358] * vector[33] +matrix[34][358] * vector[34] +matrix[35][358] * vector[35] +matrix[36][358] * vector[36] +matrix[37][358] * vector[37] +matrix[38][358] * vector[38] +matrix[39][358] * vector[39] +matrix[40][358] * vector[40] +matrix[41][358] * vector[41] +matrix[42][358] * vector[42] +matrix[43][358] * vector[43] +matrix[44][358] * vector[44] +matrix[45][358] * vector[45] +matrix[46][358] * vector[46] +matrix[47][358] * vector[47] +matrix[48][358] * vector[48] +matrix[49][358] * vector[49] +matrix[50][358] * vector[50] +matrix[51][358] * vector[51] +matrix[52][358] * vector[52] +matrix[53][358] * vector[53] +matrix[54][358] * vector[54] +matrix[55][358] * vector[55] +matrix[56][358] * vector[56] +matrix[57][358] * vector[57] +matrix[58][358] * vector[58] +matrix[59][358] * vector[59] +matrix[60][358] * vector[60] +matrix[61][358] * vector[61] +matrix[62][358] * vector[62] +matrix[63][358] * vector[63] +matrix[64][358] * vector[64] +matrix[65][358] * vector[65] +matrix[66][358] * vector[66] +matrix[67][358] * vector[67] +matrix[68][358] * vector[68] +matrix[69][358] * vector[69] +matrix[70][358] * vector[70] +matrix[71][358] * vector[71] +matrix[72][358] * vector[72] +matrix[73][358] * vector[73] +matrix[74][358] * vector[74] +matrix[75][358] * vector[75] +matrix[76][358] * vector[76] +matrix[77][358] * vector[77] +matrix[78][358] * vector[78] +matrix[79][358] * vector[79] +matrix[80][358] * vector[80] +matrix[81][358] * vector[81] +matrix[82][358] * vector[82] +matrix[83][358] * vector[83] +matrix[84][358] * vector[84] +matrix[85][358] * vector[85] +matrix[86][358] * vector[86] +matrix[87][358] * vector[87] +matrix[88][358] * vector[88] +matrix[89][358] * vector[89] +matrix[90][358] * vector[90] +matrix[91][358] * vector[91] +matrix[92][358] * vector[92] +matrix[93][358] * vector[93] +matrix[94][358] * vector[94] +matrix[95][358] * vector[95] +matrix[96][358] * vector[96] +matrix[97][358] * vector[97] +matrix[98][358] * vector[98] +matrix[99][358] * vector[99] +b[358];
assign result[359] = matrix[0][359] * vector[0] +matrix[1][359] * vector[1] +matrix[2][359] * vector[2] +matrix[3][359] * vector[3] +matrix[4][359] * vector[4] +matrix[5][359] * vector[5] +matrix[6][359] * vector[6] +matrix[7][359] * vector[7] +matrix[8][359] * vector[8] +matrix[9][359] * vector[9] +matrix[10][359] * vector[10] +matrix[11][359] * vector[11] +matrix[12][359] * vector[12] +matrix[13][359] * vector[13] +matrix[14][359] * vector[14] +matrix[15][359] * vector[15] +matrix[16][359] * vector[16] +matrix[17][359] * vector[17] +matrix[18][359] * vector[18] +matrix[19][359] * vector[19] +matrix[20][359] * vector[20] +matrix[21][359] * vector[21] +matrix[22][359] * vector[22] +matrix[23][359] * vector[23] +matrix[24][359] * vector[24] +matrix[25][359] * vector[25] +matrix[26][359] * vector[26] +matrix[27][359] * vector[27] +matrix[28][359] * vector[28] +matrix[29][359] * vector[29] +matrix[30][359] * vector[30] +matrix[31][359] * vector[31] +matrix[32][359] * vector[32] +matrix[33][359] * vector[33] +matrix[34][359] * vector[34] +matrix[35][359] * vector[35] +matrix[36][359] * vector[36] +matrix[37][359] * vector[37] +matrix[38][359] * vector[38] +matrix[39][359] * vector[39] +matrix[40][359] * vector[40] +matrix[41][359] * vector[41] +matrix[42][359] * vector[42] +matrix[43][359] * vector[43] +matrix[44][359] * vector[44] +matrix[45][359] * vector[45] +matrix[46][359] * vector[46] +matrix[47][359] * vector[47] +matrix[48][359] * vector[48] +matrix[49][359] * vector[49] +matrix[50][359] * vector[50] +matrix[51][359] * vector[51] +matrix[52][359] * vector[52] +matrix[53][359] * vector[53] +matrix[54][359] * vector[54] +matrix[55][359] * vector[55] +matrix[56][359] * vector[56] +matrix[57][359] * vector[57] +matrix[58][359] * vector[58] +matrix[59][359] * vector[59] +matrix[60][359] * vector[60] +matrix[61][359] * vector[61] +matrix[62][359] * vector[62] +matrix[63][359] * vector[63] +matrix[64][359] * vector[64] +matrix[65][359] * vector[65] +matrix[66][359] * vector[66] +matrix[67][359] * vector[67] +matrix[68][359] * vector[68] +matrix[69][359] * vector[69] +matrix[70][359] * vector[70] +matrix[71][359] * vector[71] +matrix[72][359] * vector[72] +matrix[73][359] * vector[73] +matrix[74][359] * vector[74] +matrix[75][359] * vector[75] +matrix[76][359] * vector[76] +matrix[77][359] * vector[77] +matrix[78][359] * vector[78] +matrix[79][359] * vector[79] +matrix[80][359] * vector[80] +matrix[81][359] * vector[81] +matrix[82][359] * vector[82] +matrix[83][359] * vector[83] +matrix[84][359] * vector[84] +matrix[85][359] * vector[85] +matrix[86][359] * vector[86] +matrix[87][359] * vector[87] +matrix[88][359] * vector[88] +matrix[89][359] * vector[89] +matrix[90][359] * vector[90] +matrix[91][359] * vector[91] +matrix[92][359] * vector[92] +matrix[93][359] * vector[93] +matrix[94][359] * vector[94] +matrix[95][359] * vector[95] +matrix[96][359] * vector[96] +matrix[97][359] * vector[97] +matrix[98][359] * vector[98] +matrix[99][359] * vector[99] +b[359];
assign result[360] = matrix[0][360] * vector[0] +matrix[1][360] * vector[1] +matrix[2][360] * vector[2] +matrix[3][360] * vector[3] +matrix[4][360] * vector[4] +matrix[5][360] * vector[5] +matrix[6][360] * vector[6] +matrix[7][360] * vector[7] +matrix[8][360] * vector[8] +matrix[9][360] * vector[9] +matrix[10][360] * vector[10] +matrix[11][360] * vector[11] +matrix[12][360] * vector[12] +matrix[13][360] * vector[13] +matrix[14][360] * vector[14] +matrix[15][360] * vector[15] +matrix[16][360] * vector[16] +matrix[17][360] * vector[17] +matrix[18][360] * vector[18] +matrix[19][360] * vector[19] +matrix[20][360] * vector[20] +matrix[21][360] * vector[21] +matrix[22][360] * vector[22] +matrix[23][360] * vector[23] +matrix[24][360] * vector[24] +matrix[25][360] * vector[25] +matrix[26][360] * vector[26] +matrix[27][360] * vector[27] +matrix[28][360] * vector[28] +matrix[29][360] * vector[29] +matrix[30][360] * vector[30] +matrix[31][360] * vector[31] +matrix[32][360] * vector[32] +matrix[33][360] * vector[33] +matrix[34][360] * vector[34] +matrix[35][360] * vector[35] +matrix[36][360] * vector[36] +matrix[37][360] * vector[37] +matrix[38][360] * vector[38] +matrix[39][360] * vector[39] +matrix[40][360] * vector[40] +matrix[41][360] * vector[41] +matrix[42][360] * vector[42] +matrix[43][360] * vector[43] +matrix[44][360] * vector[44] +matrix[45][360] * vector[45] +matrix[46][360] * vector[46] +matrix[47][360] * vector[47] +matrix[48][360] * vector[48] +matrix[49][360] * vector[49] +matrix[50][360] * vector[50] +matrix[51][360] * vector[51] +matrix[52][360] * vector[52] +matrix[53][360] * vector[53] +matrix[54][360] * vector[54] +matrix[55][360] * vector[55] +matrix[56][360] * vector[56] +matrix[57][360] * vector[57] +matrix[58][360] * vector[58] +matrix[59][360] * vector[59] +matrix[60][360] * vector[60] +matrix[61][360] * vector[61] +matrix[62][360] * vector[62] +matrix[63][360] * vector[63] +matrix[64][360] * vector[64] +matrix[65][360] * vector[65] +matrix[66][360] * vector[66] +matrix[67][360] * vector[67] +matrix[68][360] * vector[68] +matrix[69][360] * vector[69] +matrix[70][360] * vector[70] +matrix[71][360] * vector[71] +matrix[72][360] * vector[72] +matrix[73][360] * vector[73] +matrix[74][360] * vector[74] +matrix[75][360] * vector[75] +matrix[76][360] * vector[76] +matrix[77][360] * vector[77] +matrix[78][360] * vector[78] +matrix[79][360] * vector[79] +matrix[80][360] * vector[80] +matrix[81][360] * vector[81] +matrix[82][360] * vector[82] +matrix[83][360] * vector[83] +matrix[84][360] * vector[84] +matrix[85][360] * vector[85] +matrix[86][360] * vector[86] +matrix[87][360] * vector[87] +matrix[88][360] * vector[88] +matrix[89][360] * vector[89] +matrix[90][360] * vector[90] +matrix[91][360] * vector[91] +matrix[92][360] * vector[92] +matrix[93][360] * vector[93] +matrix[94][360] * vector[94] +matrix[95][360] * vector[95] +matrix[96][360] * vector[96] +matrix[97][360] * vector[97] +matrix[98][360] * vector[98] +matrix[99][360] * vector[99] +b[360];
assign result[361] = matrix[0][361] * vector[0] +matrix[1][361] * vector[1] +matrix[2][361] * vector[2] +matrix[3][361] * vector[3] +matrix[4][361] * vector[4] +matrix[5][361] * vector[5] +matrix[6][361] * vector[6] +matrix[7][361] * vector[7] +matrix[8][361] * vector[8] +matrix[9][361] * vector[9] +matrix[10][361] * vector[10] +matrix[11][361] * vector[11] +matrix[12][361] * vector[12] +matrix[13][361] * vector[13] +matrix[14][361] * vector[14] +matrix[15][361] * vector[15] +matrix[16][361] * vector[16] +matrix[17][361] * vector[17] +matrix[18][361] * vector[18] +matrix[19][361] * vector[19] +matrix[20][361] * vector[20] +matrix[21][361] * vector[21] +matrix[22][361] * vector[22] +matrix[23][361] * vector[23] +matrix[24][361] * vector[24] +matrix[25][361] * vector[25] +matrix[26][361] * vector[26] +matrix[27][361] * vector[27] +matrix[28][361] * vector[28] +matrix[29][361] * vector[29] +matrix[30][361] * vector[30] +matrix[31][361] * vector[31] +matrix[32][361] * vector[32] +matrix[33][361] * vector[33] +matrix[34][361] * vector[34] +matrix[35][361] * vector[35] +matrix[36][361] * vector[36] +matrix[37][361] * vector[37] +matrix[38][361] * vector[38] +matrix[39][361] * vector[39] +matrix[40][361] * vector[40] +matrix[41][361] * vector[41] +matrix[42][361] * vector[42] +matrix[43][361] * vector[43] +matrix[44][361] * vector[44] +matrix[45][361] * vector[45] +matrix[46][361] * vector[46] +matrix[47][361] * vector[47] +matrix[48][361] * vector[48] +matrix[49][361] * vector[49] +matrix[50][361] * vector[50] +matrix[51][361] * vector[51] +matrix[52][361] * vector[52] +matrix[53][361] * vector[53] +matrix[54][361] * vector[54] +matrix[55][361] * vector[55] +matrix[56][361] * vector[56] +matrix[57][361] * vector[57] +matrix[58][361] * vector[58] +matrix[59][361] * vector[59] +matrix[60][361] * vector[60] +matrix[61][361] * vector[61] +matrix[62][361] * vector[62] +matrix[63][361] * vector[63] +matrix[64][361] * vector[64] +matrix[65][361] * vector[65] +matrix[66][361] * vector[66] +matrix[67][361] * vector[67] +matrix[68][361] * vector[68] +matrix[69][361] * vector[69] +matrix[70][361] * vector[70] +matrix[71][361] * vector[71] +matrix[72][361] * vector[72] +matrix[73][361] * vector[73] +matrix[74][361] * vector[74] +matrix[75][361] * vector[75] +matrix[76][361] * vector[76] +matrix[77][361] * vector[77] +matrix[78][361] * vector[78] +matrix[79][361] * vector[79] +matrix[80][361] * vector[80] +matrix[81][361] * vector[81] +matrix[82][361] * vector[82] +matrix[83][361] * vector[83] +matrix[84][361] * vector[84] +matrix[85][361] * vector[85] +matrix[86][361] * vector[86] +matrix[87][361] * vector[87] +matrix[88][361] * vector[88] +matrix[89][361] * vector[89] +matrix[90][361] * vector[90] +matrix[91][361] * vector[91] +matrix[92][361] * vector[92] +matrix[93][361] * vector[93] +matrix[94][361] * vector[94] +matrix[95][361] * vector[95] +matrix[96][361] * vector[96] +matrix[97][361] * vector[97] +matrix[98][361] * vector[98] +matrix[99][361] * vector[99] +b[361];
assign result[362] = matrix[0][362] * vector[0] +matrix[1][362] * vector[1] +matrix[2][362] * vector[2] +matrix[3][362] * vector[3] +matrix[4][362] * vector[4] +matrix[5][362] * vector[5] +matrix[6][362] * vector[6] +matrix[7][362] * vector[7] +matrix[8][362] * vector[8] +matrix[9][362] * vector[9] +matrix[10][362] * vector[10] +matrix[11][362] * vector[11] +matrix[12][362] * vector[12] +matrix[13][362] * vector[13] +matrix[14][362] * vector[14] +matrix[15][362] * vector[15] +matrix[16][362] * vector[16] +matrix[17][362] * vector[17] +matrix[18][362] * vector[18] +matrix[19][362] * vector[19] +matrix[20][362] * vector[20] +matrix[21][362] * vector[21] +matrix[22][362] * vector[22] +matrix[23][362] * vector[23] +matrix[24][362] * vector[24] +matrix[25][362] * vector[25] +matrix[26][362] * vector[26] +matrix[27][362] * vector[27] +matrix[28][362] * vector[28] +matrix[29][362] * vector[29] +matrix[30][362] * vector[30] +matrix[31][362] * vector[31] +matrix[32][362] * vector[32] +matrix[33][362] * vector[33] +matrix[34][362] * vector[34] +matrix[35][362] * vector[35] +matrix[36][362] * vector[36] +matrix[37][362] * vector[37] +matrix[38][362] * vector[38] +matrix[39][362] * vector[39] +matrix[40][362] * vector[40] +matrix[41][362] * vector[41] +matrix[42][362] * vector[42] +matrix[43][362] * vector[43] +matrix[44][362] * vector[44] +matrix[45][362] * vector[45] +matrix[46][362] * vector[46] +matrix[47][362] * vector[47] +matrix[48][362] * vector[48] +matrix[49][362] * vector[49] +matrix[50][362] * vector[50] +matrix[51][362] * vector[51] +matrix[52][362] * vector[52] +matrix[53][362] * vector[53] +matrix[54][362] * vector[54] +matrix[55][362] * vector[55] +matrix[56][362] * vector[56] +matrix[57][362] * vector[57] +matrix[58][362] * vector[58] +matrix[59][362] * vector[59] +matrix[60][362] * vector[60] +matrix[61][362] * vector[61] +matrix[62][362] * vector[62] +matrix[63][362] * vector[63] +matrix[64][362] * vector[64] +matrix[65][362] * vector[65] +matrix[66][362] * vector[66] +matrix[67][362] * vector[67] +matrix[68][362] * vector[68] +matrix[69][362] * vector[69] +matrix[70][362] * vector[70] +matrix[71][362] * vector[71] +matrix[72][362] * vector[72] +matrix[73][362] * vector[73] +matrix[74][362] * vector[74] +matrix[75][362] * vector[75] +matrix[76][362] * vector[76] +matrix[77][362] * vector[77] +matrix[78][362] * vector[78] +matrix[79][362] * vector[79] +matrix[80][362] * vector[80] +matrix[81][362] * vector[81] +matrix[82][362] * vector[82] +matrix[83][362] * vector[83] +matrix[84][362] * vector[84] +matrix[85][362] * vector[85] +matrix[86][362] * vector[86] +matrix[87][362] * vector[87] +matrix[88][362] * vector[88] +matrix[89][362] * vector[89] +matrix[90][362] * vector[90] +matrix[91][362] * vector[91] +matrix[92][362] * vector[92] +matrix[93][362] * vector[93] +matrix[94][362] * vector[94] +matrix[95][362] * vector[95] +matrix[96][362] * vector[96] +matrix[97][362] * vector[97] +matrix[98][362] * vector[98] +matrix[99][362] * vector[99] +b[362];
assign result[363] = matrix[0][363] * vector[0] +matrix[1][363] * vector[1] +matrix[2][363] * vector[2] +matrix[3][363] * vector[3] +matrix[4][363] * vector[4] +matrix[5][363] * vector[5] +matrix[6][363] * vector[6] +matrix[7][363] * vector[7] +matrix[8][363] * vector[8] +matrix[9][363] * vector[9] +matrix[10][363] * vector[10] +matrix[11][363] * vector[11] +matrix[12][363] * vector[12] +matrix[13][363] * vector[13] +matrix[14][363] * vector[14] +matrix[15][363] * vector[15] +matrix[16][363] * vector[16] +matrix[17][363] * vector[17] +matrix[18][363] * vector[18] +matrix[19][363] * vector[19] +matrix[20][363] * vector[20] +matrix[21][363] * vector[21] +matrix[22][363] * vector[22] +matrix[23][363] * vector[23] +matrix[24][363] * vector[24] +matrix[25][363] * vector[25] +matrix[26][363] * vector[26] +matrix[27][363] * vector[27] +matrix[28][363] * vector[28] +matrix[29][363] * vector[29] +matrix[30][363] * vector[30] +matrix[31][363] * vector[31] +matrix[32][363] * vector[32] +matrix[33][363] * vector[33] +matrix[34][363] * vector[34] +matrix[35][363] * vector[35] +matrix[36][363] * vector[36] +matrix[37][363] * vector[37] +matrix[38][363] * vector[38] +matrix[39][363] * vector[39] +matrix[40][363] * vector[40] +matrix[41][363] * vector[41] +matrix[42][363] * vector[42] +matrix[43][363] * vector[43] +matrix[44][363] * vector[44] +matrix[45][363] * vector[45] +matrix[46][363] * vector[46] +matrix[47][363] * vector[47] +matrix[48][363] * vector[48] +matrix[49][363] * vector[49] +matrix[50][363] * vector[50] +matrix[51][363] * vector[51] +matrix[52][363] * vector[52] +matrix[53][363] * vector[53] +matrix[54][363] * vector[54] +matrix[55][363] * vector[55] +matrix[56][363] * vector[56] +matrix[57][363] * vector[57] +matrix[58][363] * vector[58] +matrix[59][363] * vector[59] +matrix[60][363] * vector[60] +matrix[61][363] * vector[61] +matrix[62][363] * vector[62] +matrix[63][363] * vector[63] +matrix[64][363] * vector[64] +matrix[65][363] * vector[65] +matrix[66][363] * vector[66] +matrix[67][363] * vector[67] +matrix[68][363] * vector[68] +matrix[69][363] * vector[69] +matrix[70][363] * vector[70] +matrix[71][363] * vector[71] +matrix[72][363] * vector[72] +matrix[73][363] * vector[73] +matrix[74][363] * vector[74] +matrix[75][363] * vector[75] +matrix[76][363] * vector[76] +matrix[77][363] * vector[77] +matrix[78][363] * vector[78] +matrix[79][363] * vector[79] +matrix[80][363] * vector[80] +matrix[81][363] * vector[81] +matrix[82][363] * vector[82] +matrix[83][363] * vector[83] +matrix[84][363] * vector[84] +matrix[85][363] * vector[85] +matrix[86][363] * vector[86] +matrix[87][363] * vector[87] +matrix[88][363] * vector[88] +matrix[89][363] * vector[89] +matrix[90][363] * vector[90] +matrix[91][363] * vector[91] +matrix[92][363] * vector[92] +matrix[93][363] * vector[93] +matrix[94][363] * vector[94] +matrix[95][363] * vector[95] +matrix[96][363] * vector[96] +matrix[97][363] * vector[97] +matrix[98][363] * vector[98] +matrix[99][363] * vector[99] +b[363];
assign result[364] = matrix[0][364] * vector[0] +matrix[1][364] * vector[1] +matrix[2][364] * vector[2] +matrix[3][364] * vector[3] +matrix[4][364] * vector[4] +matrix[5][364] * vector[5] +matrix[6][364] * vector[6] +matrix[7][364] * vector[7] +matrix[8][364] * vector[8] +matrix[9][364] * vector[9] +matrix[10][364] * vector[10] +matrix[11][364] * vector[11] +matrix[12][364] * vector[12] +matrix[13][364] * vector[13] +matrix[14][364] * vector[14] +matrix[15][364] * vector[15] +matrix[16][364] * vector[16] +matrix[17][364] * vector[17] +matrix[18][364] * vector[18] +matrix[19][364] * vector[19] +matrix[20][364] * vector[20] +matrix[21][364] * vector[21] +matrix[22][364] * vector[22] +matrix[23][364] * vector[23] +matrix[24][364] * vector[24] +matrix[25][364] * vector[25] +matrix[26][364] * vector[26] +matrix[27][364] * vector[27] +matrix[28][364] * vector[28] +matrix[29][364] * vector[29] +matrix[30][364] * vector[30] +matrix[31][364] * vector[31] +matrix[32][364] * vector[32] +matrix[33][364] * vector[33] +matrix[34][364] * vector[34] +matrix[35][364] * vector[35] +matrix[36][364] * vector[36] +matrix[37][364] * vector[37] +matrix[38][364] * vector[38] +matrix[39][364] * vector[39] +matrix[40][364] * vector[40] +matrix[41][364] * vector[41] +matrix[42][364] * vector[42] +matrix[43][364] * vector[43] +matrix[44][364] * vector[44] +matrix[45][364] * vector[45] +matrix[46][364] * vector[46] +matrix[47][364] * vector[47] +matrix[48][364] * vector[48] +matrix[49][364] * vector[49] +matrix[50][364] * vector[50] +matrix[51][364] * vector[51] +matrix[52][364] * vector[52] +matrix[53][364] * vector[53] +matrix[54][364] * vector[54] +matrix[55][364] * vector[55] +matrix[56][364] * vector[56] +matrix[57][364] * vector[57] +matrix[58][364] * vector[58] +matrix[59][364] * vector[59] +matrix[60][364] * vector[60] +matrix[61][364] * vector[61] +matrix[62][364] * vector[62] +matrix[63][364] * vector[63] +matrix[64][364] * vector[64] +matrix[65][364] * vector[65] +matrix[66][364] * vector[66] +matrix[67][364] * vector[67] +matrix[68][364] * vector[68] +matrix[69][364] * vector[69] +matrix[70][364] * vector[70] +matrix[71][364] * vector[71] +matrix[72][364] * vector[72] +matrix[73][364] * vector[73] +matrix[74][364] * vector[74] +matrix[75][364] * vector[75] +matrix[76][364] * vector[76] +matrix[77][364] * vector[77] +matrix[78][364] * vector[78] +matrix[79][364] * vector[79] +matrix[80][364] * vector[80] +matrix[81][364] * vector[81] +matrix[82][364] * vector[82] +matrix[83][364] * vector[83] +matrix[84][364] * vector[84] +matrix[85][364] * vector[85] +matrix[86][364] * vector[86] +matrix[87][364] * vector[87] +matrix[88][364] * vector[88] +matrix[89][364] * vector[89] +matrix[90][364] * vector[90] +matrix[91][364] * vector[91] +matrix[92][364] * vector[92] +matrix[93][364] * vector[93] +matrix[94][364] * vector[94] +matrix[95][364] * vector[95] +matrix[96][364] * vector[96] +matrix[97][364] * vector[97] +matrix[98][364] * vector[98] +matrix[99][364] * vector[99] +b[364];
assign result[365] = matrix[0][365] * vector[0] +matrix[1][365] * vector[1] +matrix[2][365] * vector[2] +matrix[3][365] * vector[3] +matrix[4][365] * vector[4] +matrix[5][365] * vector[5] +matrix[6][365] * vector[6] +matrix[7][365] * vector[7] +matrix[8][365] * vector[8] +matrix[9][365] * vector[9] +matrix[10][365] * vector[10] +matrix[11][365] * vector[11] +matrix[12][365] * vector[12] +matrix[13][365] * vector[13] +matrix[14][365] * vector[14] +matrix[15][365] * vector[15] +matrix[16][365] * vector[16] +matrix[17][365] * vector[17] +matrix[18][365] * vector[18] +matrix[19][365] * vector[19] +matrix[20][365] * vector[20] +matrix[21][365] * vector[21] +matrix[22][365] * vector[22] +matrix[23][365] * vector[23] +matrix[24][365] * vector[24] +matrix[25][365] * vector[25] +matrix[26][365] * vector[26] +matrix[27][365] * vector[27] +matrix[28][365] * vector[28] +matrix[29][365] * vector[29] +matrix[30][365] * vector[30] +matrix[31][365] * vector[31] +matrix[32][365] * vector[32] +matrix[33][365] * vector[33] +matrix[34][365] * vector[34] +matrix[35][365] * vector[35] +matrix[36][365] * vector[36] +matrix[37][365] * vector[37] +matrix[38][365] * vector[38] +matrix[39][365] * vector[39] +matrix[40][365] * vector[40] +matrix[41][365] * vector[41] +matrix[42][365] * vector[42] +matrix[43][365] * vector[43] +matrix[44][365] * vector[44] +matrix[45][365] * vector[45] +matrix[46][365] * vector[46] +matrix[47][365] * vector[47] +matrix[48][365] * vector[48] +matrix[49][365] * vector[49] +matrix[50][365] * vector[50] +matrix[51][365] * vector[51] +matrix[52][365] * vector[52] +matrix[53][365] * vector[53] +matrix[54][365] * vector[54] +matrix[55][365] * vector[55] +matrix[56][365] * vector[56] +matrix[57][365] * vector[57] +matrix[58][365] * vector[58] +matrix[59][365] * vector[59] +matrix[60][365] * vector[60] +matrix[61][365] * vector[61] +matrix[62][365] * vector[62] +matrix[63][365] * vector[63] +matrix[64][365] * vector[64] +matrix[65][365] * vector[65] +matrix[66][365] * vector[66] +matrix[67][365] * vector[67] +matrix[68][365] * vector[68] +matrix[69][365] * vector[69] +matrix[70][365] * vector[70] +matrix[71][365] * vector[71] +matrix[72][365] * vector[72] +matrix[73][365] * vector[73] +matrix[74][365] * vector[74] +matrix[75][365] * vector[75] +matrix[76][365] * vector[76] +matrix[77][365] * vector[77] +matrix[78][365] * vector[78] +matrix[79][365] * vector[79] +matrix[80][365] * vector[80] +matrix[81][365] * vector[81] +matrix[82][365] * vector[82] +matrix[83][365] * vector[83] +matrix[84][365] * vector[84] +matrix[85][365] * vector[85] +matrix[86][365] * vector[86] +matrix[87][365] * vector[87] +matrix[88][365] * vector[88] +matrix[89][365] * vector[89] +matrix[90][365] * vector[90] +matrix[91][365] * vector[91] +matrix[92][365] * vector[92] +matrix[93][365] * vector[93] +matrix[94][365] * vector[94] +matrix[95][365] * vector[95] +matrix[96][365] * vector[96] +matrix[97][365] * vector[97] +matrix[98][365] * vector[98] +matrix[99][365] * vector[99] +b[365];
assign result[366] = matrix[0][366] * vector[0] +matrix[1][366] * vector[1] +matrix[2][366] * vector[2] +matrix[3][366] * vector[3] +matrix[4][366] * vector[4] +matrix[5][366] * vector[5] +matrix[6][366] * vector[6] +matrix[7][366] * vector[7] +matrix[8][366] * vector[8] +matrix[9][366] * vector[9] +matrix[10][366] * vector[10] +matrix[11][366] * vector[11] +matrix[12][366] * vector[12] +matrix[13][366] * vector[13] +matrix[14][366] * vector[14] +matrix[15][366] * vector[15] +matrix[16][366] * vector[16] +matrix[17][366] * vector[17] +matrix[18][366] * vector[18] +matrix[19][366] * vector[19] +matrix[20][366] * vector[20] +matrix[21][366] * vector[21] +matrix[22][366] * vector[22] +matrix[23][366] * vector[23] +matrix[24][366] * vector[24] +matrix[25][366] * vector[25] +matrix[26][366] * vector[26] +matrix[27][366] * vector[27] +matrix[28][366] * vector[28] +matrix[29][366] * vector[29] +matrix[30][366] * vector[30] +matrix[31][366] * vector[31] +matrix[32][366] * vector[32] +matrix[33][366] * vector[33] +matrix[34][366] * vector[34] +matrix[35][366] * vector[35] +matrix[36][366] * vector[36] +matrix[37][366] * vector[37] +matrix[38][366] * vector[38] +matrix[39][366] * vector[39] +matrix[40][366] * vector[40] +matrix[41][366] * vector[41] +matrix[42][366] * vector[42] +matrix[43][366] * vector[43] +matrix[44][366] * vector[44] +matrix[45][366] * vector[45] +matrix[46][366] * vector[46] +matrix[47][366] * vector[47] +matrix[48][366] * vector[48] +matrix[49][366] * vector[49] +matrix[50][366] * vector[50] +matrix[51][366] * vector[51] +matrix[52][366] * vector[52] +matrix[53][366] * vector[53] +matrix[54][366] * vector[54] +matrix[55][366] * vector[55] +matrix[56][366] * vector[56] +matrix[57][366] * vector[57] +matrix[58][366] * vector[58] +matrix[59][366] * vector[59] +matrix[60][366] * vector[60] +matrix[61][366] * vector[61] +matrix[62][366] * vector[62] +matrix[63][366] * vector[63] +matrix[64][366] * vector[64] +matrix[65][366] * vector[65] +matrix[66][366] * vector[66] +matrix[67][366] * vector[67] +matrix[68][366] * vector[68] +matrix[69][366] * vector[69] +matrix[70][366] * vector[70] +matrix[71][366] * vector[71] +matrix[72][366] * vector[72] +matrix[73][366] * vector[73] +matrix[74][366] * vector[74] +matrix[75][366] * vector[75] +matrix[76][366] * vector[76] +matrix[77][366] * vector[77] +matrix[78][366] * vector[78] +matrix[79][366] * vector[79] +matrix[80][366] * vector[80] +matrix[81][366] * vector[81] +matrix[82][366] * vector[82] +matrix[83][366] * vector[83] +matrix[84][366] * vector[84] +matrix[85][366] * vector[85] +matrix[86][366] * vector[86] +matrix[87][366] * vector[87] +matrix[88][366] * vector[88] +matrix[89][366] * vector[89] +matrix[90][366] * vector[90] +matrix[91][366] * vector[91] +matrix[92][366] * vector[92] +matrix[93][366] * vector[93] +matrix[94][366] * vector[94] +matrix[95][366] * vector[95] +matrix[96][366] * vector[96] +matrix[97][366] * vector[97] +matrix[98][366] * vector[98] +matrix[99][366] * vector[99] +b[366];
assign result[367] = matrix[0][367] * vector[0] +matrix[1][367] * vector[1] +matrix[2][367] * vector[2] +matrix[3][367] * vector[3] +matrix[4][367] * vector[4] +matrix[5][367] * vector[5] +matrix[6][367] * vector[6] +matrix[7][367] * vector[7] +matrix[8][367] * vector[8] +matrix[9][367] * vector[9] +matrix[10][367] * vector[10] +matrix[11][367] * vector[11] +matrix[12][367] * vector[12] +matrix[13][367] * vector[13] +matrix[14][367] * vector[14] +matrix[15][367] * vector[15] +matrix[16][367] * vector[16] +matrix[17][367] * vector[17] +matrix[18][367] * vector[18] +matrix[19][367] * vector[19] +matrix[20][367] * vector[20] +matrix[21][367] * vector[21] +matrix[22][367] * vector[22] +matrix[23][367] * vector[23] +matrix[24][367] * vector[24] +matrix[25][367] * vector[25] +matrix[26][367] * vector[26] +matrix[27][367] * vector[27] +matrix[28][367] * vector[28] +matrix[29][367] * vector[29] +matrix[30][367] * vector[30] +matrix[31][367] * vector[31] +matrix[32][367] * vector[32] +matrix[33][367] * vector[33] +matrix[34][367] * vector[34] +matrix[35][367] * vector[35] +matrix[36][367] * vector[36] +matrix[37][367] * vector[37] +matrix[38][367] * vector[38] +matrix[39][367] * vector[39] +matrix[40][367] * vector[40] +matrix[41][367] * vector[41] +matrix[42][367] * vector[42] +matrix[43][367] * vector[43] +matrix[44][367] * vector[44] +matrix[45][367] * vector[45] +matrix[46][367] * vector[46] +matrix[47][367] * vector[47] +matrix[48][367] * vector[48] +matrix[49][367] * vector[49] +matrix[50][367] * vector[50] +matrix[51][367] * vector[51] +matrix[52][367] * vector[52] +matrix[53][367] * vector[53] +matrix[54][367] * vector[54] +matrix[55][367] * vector[55] +matrix[56][367] * vector[56] +matrix[57][367] * vector[57] +matrix[58][367] * vector[58] +matrix[59][367] * vector[59] +matrix[60][367] * vector[60] +matrix[61][367] * vector[61] +matrix[62][367] * vector[62] +matrix[63][367] * vector[63] +matrix[64][367] * vector[64] +matrix[65][367] * vector[65] +matrix[66][367] * vector[66] +matrix[67][367] * vector[67] +matrix[68][367] * vector[68] +matrix[69][367] * vector[69] +matrix[70][367] * vector[70] +matrix[71][367] * vector[71] +matrix[72][367] * vector[72] +matrix[73][367] * vector[73] +matrix[74][367] * vector[74] +matrix[75][367] * vector[75] +matrix[76][367] * vector[76] +matrix[77][367] * vector[77] +matrix[78][367] * vector[78] +matrix[79][367] * vector[79] +matrix[80][367] * vector[80] +matrix[81][367] * vector[81] +matrix[82][367] * vector[82] +matrix[83][367] * vector[83] +matrix[84][367] * vector[84] +matrix[85][367] * vector[85] +matrix[86][367] * vector[86] +matrix[87][367] * vector[87] +matrix[88][367] * vector[88] +matrix[89][367] * vector[89] +matrix[90][367] * vector[90] +matrix[91][367] * vector[91] +matrix[92][367] * vector[92] +matrix[93][367] * vector[93] +matrix[94][367] * vector[94] +matrix[95][367] * vector[95] +matrix[96][367] * vector[96] +matrix[97][367] * vector[97] +matrix[98][367] * vector[98] +matrix[99][367] * vector[99] +b[367];
assign result[368] = matrix[0][368] * vector[0] +matrix[1][368] * vector[1] +matrix[2][368] * vector[2] +matrix[3][368] * vector[3] +matrix[4][368] * vector[4] +matrix[5][368] * vector[5] +matrix[6][368] * vector[6] +matrix[7][368] * vector[7] +matrix[8][368] * vector[8] +matrix[9][368] * vector[9] +matrix[10][368] * vector[10] +matrix[11][368] * vector[11] +matrix[12][368] * vector[12] +matrix[13][368] * vector[13] +matrix[14][368] * vector[14] +matrix[15][368] * vector[15] +matrix[16][368] * vector[16] +matrix[17][368] * vector[17] +matrix[18][368] * vector[18] +matrix[19][368] * vector[19] +matrix[20][368] * vector[20] +matrix[21][368] * vector[21] +matrix[22][368] * vector[22] +matrix[23][368] * vector[23] +matrix[24][368] * vector[24] +matrix[25][368] * vector[25] +matrix[26][368] * vector[26] +matrix[27][368] * vector[27] +matrix[28][368] * vector[28] +matrix[29][368] * vector[29] +matrix[30][368] * vector[30] +matrix[31][368] * vector[31] +matrix[32][368] * vector[32] +matrix[33][368] * vector[33] +matrix[34][368] * vector[34] +matrix[35][368] * vector[35] +matrix[36][368] * vector[36] +matrix[37][368] * vector[37] +matrix[38][368] * vector[38] +matrix[39][368] * vector[39] +matrix[40][368] * vector[40] +matrix[41][368] * vector[41] +matrix[42][368] * vector[42] +matrix[43][368] * vector[43] +matrix[44][368] * vector[44] +matrix[45][368] * vector[45] +matrix[46][368] * vector[46] +matrix[47][368] * vector[47] +matrix[48][368] * vector[48] +matrix[49][368] * vector[49] +matrix[50][368] * vector[50] +matrix[51][368] * vector[51] +matrix[52][368] * vector[52] +matrix[53][368] * vector[53] +matrix[54][368] * vector[54] +matrix[55][368] * vector[55] +matrix[56][368] * vector[56] +matrix[57][368] * vector[57] +matrix[58][368] * vector[58] +matrix[59][368] * vector[59] +matrix[60][368] * vector[60] +matrix[61][368] * vector[61] +matrix[62][368] * vector[62] +matrix[63][368] * vector[63] +matrix[64][368] * vector[64] +matrix[65][368] * vector[65] +matrix[66][368] * vector[66] +matrix[67][368] * vector[67] +matrix[68][368] * vector[68] +matrix[69][368] * vector[69] +matrix[70][368] * vector[70] +matrix[71][368] * vector[71] +matrix[72][368] * vector[72] +matrix[73][368] * vector[73] +matrix[74][368] * vector[74] +matrix[75][368] * vector[75] +matrix[76][368] * vector[76] +matrix[77][368] * vector[77] +matrix[78][368] * vector[78] +matrix[79][368] * vector[79] +matrix[80][368] * vector[80] +matrix[81][368] * vector[81] +matrix[82][368] * vector[82] +matrix[83][368] * vector[83] +matrix[84][368] * vector[84] +matrix[85][368] * vector[85] +matrix[86][368] * vector[86] +matrix[87][368] * vector[87] +matrix[88][368] * vector[88] +matrix[89][368] * vector[89] +matrix[90][368] * vector[90] +matrix[91][368] * vector[91] +matrix[92][368] * vector[92] +matrix[93][368] * vector[93] +matrix[94][368] * vector[94] +matrix[95][368] * vector[95] +matrix[96][368] * vector[96] +matrix[97][368] * vector[97] +matrix[98][368] * vector[98] +matrix[99][368] * vector[99] +b[368];
assign result[369] = matrix[0][369] * vector[0] +matrix[1][369] * vector[1] +matrix[2][369] * vector[2] +matrix[3][369] * vector[3] +matrix[4][369] * vector[4] +matrix[5][369] * vector[5] +matrix[6][369] * vector[6] +matrix[7][369] * vector[7] +matrix[8][369] * vector[8] +matrix[9][369] * vector[9] +matrix[10][369] * vector[10] +matrix[11][369] * vector[11] +matrix[12][369] * vector[12] +matrix[13][369] * vector[13] +matrix[14][369] * vector[14] +matrix[15][369] * vector[15] +matrix[16][369] * vector[16] +matrix[17][369] * vector[17] +matrix[18][369] * vector[18] +matrix[19][369] * vector[19] +matrix[20][369] * vector[20] +matrix[21][369] * vector[21] +matrix[22][369] * vector[22] +matrix[23][369] * vector[23] +matrix[24][369] * vector[24] +matrix[25][369] * vector[25] +matrix[26][369] * vector[26] +matrix[27][369] * vector[27] +matrix[28][369] * vector[28] +matrix[29][369] * vector[29] +matrix[30][369] * vector[30] +matrix[31][369] * vector[31] +matrix[32][369] * vector[32] +matrix[33][369] * vector[33] +matrix[34][369] * vector[34] +matrix[35][369] * vector[35] +matrix[36][369] * vector[36] +matrix[37][369] * vector[37] +matrix[38][369] * vector[38] +matrix[39][369] * vector[39] +matrix[40][369] * vector[40] +matrix[41][369] * vector[41] +matrix[42][369] * vector[42] +matrix[43][369] * vector[43] +matrix[44][369] * vector[44] +matrix[45][369] * vector[45] +matrix[46][369] * vector[46] +matrix[47][369] * vector[47] +matrix[48][369] * vector[48] +matrix[49][369] * vector[49] +matrix[50][369] * vector[50] +matrix[51][369] * vector[51] +matrix[52][369] * vector[52] +matrix[53][369] * vector[53] +matrix[54][369] * vector[54] +matrix[55][369] * vector[55] +matrix[56][369] * vector[56] +matrix[57][369] * vector[57] +matrix[58][369] * vector[58] +matrix[59][369] * vector[59] +matrix[60][369] * vector[60] +matrix[61][369] * vector[61] +matrix[62][369] * vector[62] +matrix[63][369] * vector[63] +matrix[64][369] * vector[64] +matrix[65][369] * vector[65] +matrix[66][369] * vector[66] +matrix[67][369] * vector[67] +matrix[68][369] * vector[68] +matrix[69][369] * vector[69] +matrix[70][369] * vector[70] +matrix[71][369] * vector[71] +matrix[72][369] * vector[72] +matrix[73][369] * vector[73] +matrix[74][369] * vector[74] +matrix[75][369] * vector[75] +matrix[76][369] * vector[76] +matrix[77][369] * vector[77] +matrix[78][369] * vector[78] +matrix[79][369] * vector[79] +matrix[80][369] * vector[80] +matrix[81][369] * vector[81] +matrix[82][369] * vector[82] +matrix[83][369] * vector[83] +matrix[84][369] * vector[84] +matrix[85][369] * vector[85] +matrix[86][369] * vector[86] +matrix[87][369] * vector[87] +matrix[88][369] * vector[88] +matrix[89][369] * vector[89] +matrix[90][369] * vector[90] +matrix[91][369] * vector[91] +matrix[92][369] * vector[92] +matrix[93][369] * vector[93] +matrix[94][369] * vector[94] +matrix[95][369] * vector[95] +matrix[96][369] * vector[96] +matrix[97][369] * vector[97] +matrix[98][369] * vector[98] +matrix[99][369] * vector[99] +b[369];
assign result[370] = matrix[0][370] * vector[0] +matrix[1][370] * vector[1] +matrix[2][370] * vector[2] +matrix[3][370] * vector[3] +matrix[4][370] * vector[4] +matrix[5][370] * vector[5] +matrix[6][370] * vector[6] +matrix[7][370] * vector[7] +matrix[8][370] * vector[8] +matrix[9][370] * vector[9] +matrix[10][370] * vector[10] +matrix[11][370] * vector[11] +matrix[12][370] * vector[12] +matrix[13][370] * vector[13] +matrix[14][370] * vector[14] +matrix[15][370] * vector[15] +matrix[16][370] * vector[16] +matrix[17][370] * vector[17] +matrix[18][370] * vector[18] +matrix[19][370] * vector[19] +matrix[20][370] * vector[20] +matrix[21][370] * vector[21] +matrix[22][370] * vector[22] +matrix[23][370] * vector[23] +matrix[24][370] * vector[24] +matrix[25][370] * vector[25] +matrix[26][370] * vector[26] +matrix[27][370] * vector[27] +matrix[28][370] * vector[28] +matrix[29][370] * vector[29] +matrix[30][370] * vector[30] +matrix[31][370] * vector[31] +matrix[32][370] * vector[32] +matrix[33][370] * vector[33] +matrix[34][370] * vector[34] +matrix[35][370] * vector[35] +matrix[36][370] * vector[36] +matrix[37][370] * vector[37] +matrix[38][370] * vector[38] +matrix[39][370] * vector[39] +matrix[40][370] * vector[40] +matrix[41][370] * vector[41] +matrix[42][370] * vector[42] +matrix[43][370] * vector[43] +matrix[44][370] * vector[44] +matrix[45][370] * vector[45] +matrix[46][370] * vector[46] +matrix[47][370] * vector[47] +matrix[48][370] * vector[48] +matrix[49][370] * vector[49] +matrix[50][370] * vector[50] +matrix[51][370] * vector[51] +matrix[52][370] * vector[52] +matrix[53][370] * vector[53] +matrix[54][370] * vector[54] +matrix[55][370] * vector[55] +matrix[56][370] * vector[56] +matrix[57][370] * vector[57] +matrix[58][370] * vector[58] +matrix[59][370] * vector[59] +matrix[60][370] * vector[60] +matrix[61][370] * vector[61] +matrix[62][370] * vector[62] +matrix[63][370] * vector[63] +matrix[64][370] * vector[64] +matrix[65][370] * vector[65] +matrix[66][370] * vector[66] +matrix[67][370] * vector[67] +matrix[68][370] * vector[68] +matrix[69][370] * vector[69] +matrix[70][370] * vector[70] +matrix[71][370] * vector[71] +matrix[72][370] * vector[72] +matrix[73][370] * vector[73] +matrix[74][370] * vector[74] +matrix[75][370] * vector[75] +matrix[76][370] * vector[76] +matrix[77][370] * vector[77] +matrix[78][370] * vector[78] +matrix[79][370] * vector[79] +matrix[80][370] * vector[80] +matrix[81][370] * vector[81] +matrix[82][370] * vector[82] +matrix[83][370] * vector[83] +matrix[84][370] * vector[84] +matrix[85][370] * vector[85] +matrix[86][370] * vector[86] +matrix[87][370] * vector[87] +matrix[88][370] * vector[88] +matrix[89][370] * vector[89] +matrix[90][370] * vector[90] +matrix[91][370] * vector[91] +matrix[92][370] * vector[92] +matrix[93][370] * vector[93] +matrix[94][370] * vector[94] +matrix[95][370] * vector[95] +matrix[96][370] * vector[96] +matrix[97][370] * vector[97] +matrix[98][370] * vector[98] +matrix[99][370] * vector[99] +b[370];
assign result[371] = matrix[0][371] * vector[0] +matrix[1][371] * vector[1] +matrix[2][371] * vector[2] +matrix[3][371] * vector[3] +matrix[4][371] * vector[4] +matrix[5][371] * vector[5] +matrix[6][371] * vector[6] +matrix[7][371] * vector[7] +matrix[8][371] * vector[8] +matrix[9][371] * vector[9] +matrix[10][371] * vector[10] +matrix[11][371] * vector[11] +matrix[12][371] * vector[12] +matrix[13][371] * vector[13] +matrix[14][371] * vector[14] +matrix[15][371] * vector[15] +matrix[16][371] * vector[16] +matrix[17][371] * vector[17] +matrix[18][371] * vector[18] +matrix[19][371] * vector[19] +matrix[20][371] * vector[20] +matrix[21][371] * vector[21] +matrix[22][371] * vector[22] +matrix[23][371] * vector[23] +matrix[24][371] * vector[24] +matrix[25][371] * vector[25] +matrix[26][371] * vector[26] +matrix[27][371] * vector[27] +matrix[28][371] * vector[28] +matrix[29][371] * vector[29] +matrix[30][371] * vector[30] +matrix[31][371] * vector[31] +matrix[32][371] * vector[32] +matrix[33][371] * vector[33] +matrix[34][371] * vector[34] +matrix[35][371] * vector[35] +matrix[36][371] * vector[36] +matrix[37][371] * vector[37] +matrix[38][371] * vector[38] +matrix[39][371] * vector[39] +matrix[40][371] * vector[40] +matrix[41][371] * vector[41] +matrix[42][371] * vector[42] +matrix[43][371] * vector[43] +matrix[44][371] * vector[44] +matrix[45][371] * vector[45] +matrix[46][371] * vector[46] +matrix[47][371] * vector[47] +matrix[48][371] * vector[48] +matrix[49][371] * vector[49] +matrix[50][371] * vector[50] +matrix[51][371] * vector[51] +matrix[52][371] * vector[52] +matrix[53][371] * vector[53] +matrix[54][371] * vector[54] +matrix[55][371] * vector[55] +matrix[56][371] * vector[56] +matrix[57][371] * vector[57] +matrix[58][371] * vector[58] +matrix[59][371] * vector[59] +matrix[60][371] * vector[60] +matrix[61][371] * vector[61] +matrix[62][371] * vector[62] +matrix[63][371] * vector[63] +matrix[64][371] * vector[64] +matrix[65][371] * vector[65] +matrix[66][371] * vector[66] +matrix[67][371] * vector[67] +matrix[68][371] * vector[68] +matrix[69][371] * vector[69] +matrix[70][371] * vector[70] +matrix[71][371] * vector[71] +matrix[72][371] * vector[72] +matrix[73][371] * vector[73] +matrix[74][371] * vector[74] +matrix[75][371] * vector[75] +matrix[76][371] * vector[76] +matrix[77][371] * vector[77] +matrix[78][371] * vector[78] +matrix[79][371] * vector[79] +matrix[80][371] * vector[80] +matrix[81][371] * vector[81] +matrix[82][371] * vector[82] +matrix[83][371] * vector[83] +matrix[84][371] * vector[84] +matrix[85][371] * vector[85] +matrix[86][371] * vector[86] +matrix[87][371] * vector[87] +matrix[88][371] * vector[88] +matrix[89][371] * vector[89] +matrix[90][371] * vector[90] +matrix[91][371] * vector[91] +matrix[92][371] * vector[92] +matrix[93][371] * vector[93] +matrix[94][371] * vector[94] +matrix[95][371] * vector[95] +matrix[96][371] * vector[96] +matrix[97][371] * vector[97] +matrix[98][371] * vector[98] +matrix[99][371] * vector[99] +b[371];
assign result[372] = matrix[0][372] * vector[0] +matrix[1][372] * vector[1] +matrix[2][372] * vector[2] +matrix[3][372] * vector[3] +matrix[4][372] * vector[4] +matrix[5][372] * vector[5] +matrix[6][372] * vector[6] +matrix[7][372] * vector[7] +matrix[8][372] * vector[8] +matrix[9][372] * vector[9] +matrix[10][372] * vector[10] +matrix[11][372] * vector[11] +matrix[12][372] * vector[12] +matrix[13][372] * vector[13] +matrix[14][372] * vector[14] +matrix[15][372] * vector[15] +matrix[16][372] * vector[16] +matrix[17][372] * vector[17] +matrix[18][372] * vector[18] +matrix[19][372] * vector[19] +matrix[20][372] * vector[20] +matrix[21][372] * vector[21] +matrix[22][372] * vector[22] +matrix[23][372] * vector[23] +matrix[24][372] * vector[24] +matrix[25][372] * vector[25] +matrix[26][372] * vector[26] +matrix[27][372] * vector[27] +matrix[28][372] * vector[28] +matrix[29][372] * vector[29] +matrix[30][372] * vector[30] +matrix[31][372] * vector[31] +matrix[32][372] * vector[32] +matrix[33][372] * vector[33] +matrix[34][372] * vector[34] +matrix[35][372] * vector[35] +matrix[36][372] * vector[36] +matrix[37][372] * vector[37] +matrix[38][372] * vector[38] +matrix[39][372] * vector[39] +matrix[40][372] * vector[40] +matrix[41][372] * vector[41] +matrix[42][372] * vector[42] +matrix[43][372] * vector[43] +matrix[44][372] * vector[44] +matrix[45][372] * vector[45] +matrix[46][372] * vector[46] +matrix[47][372] * vector[47] +matrix[48][372] * vector[48] +matrix[49][372] * vector[49] +matrix[50][372] * vector[50] +matrix[51][372] * vector[51] +matrix[52][372] * vector[52] +matrix[53][372] * vector[53] +matrix[54][372] * vector[54] +matrix[55][372] * vector[55] +matrix[56][372] * vector[56] +matrix[57][372] * vector[57] +matrix[58][372] * vector[58] +matrix[59][372] * vector[59] +matrix[60][372] * vector[60] +matrix[61][372] * vector[61] +matrix[62][372] * vector[62] +matrix[63][372] * vector[63] +matrix[64][372] * vector[64] +matrix[65][372] * vector[65] +matrix[66][372] * vector[66] +matrix[67][372] * vector[67] +matrix[68][372] * vector[68] +matrix[69][372] * vector[69] +matrix[70][372] * vector[70] +matrix[71][372] * vector[71] +matrix[72][372] * vector[72] +matrix[73][372] * vector[73] +matrix[74][372] * vector[74] +matrix[75][372] * vector[75] +matrix[76][372] * vector[76] +matrix[77][372] * vector[77] +matrix[78][372] * vector[78] +matrix[79][372] * vector[79] +matrix[80][372] * vector[80] +matrix[81][372] * vector[81] +matrix[82][372] * vector[82] +matrix[83][372] * vector[83] +matrix[84][372] * vector[84] +matrix[85][372] * vector[85] +matrix[86][372] * vector[86] +matrix[87][372] * vector[87] +matrix[88][372] * vector[88] +matrix[89][372] * vector[89] +matrix[90][372] * vector[90] +matrix[91][372] * vector[91] +matrix[92][372] * vector[92] +matrix[93][372] * vector[93] +matrix[94][372] * vector[94] +matrix[95][372] * vector[95] +matrix[96][372] * vector[96] +matrix[97][372] * vector[97] +matrix[98][372] * vector[98] +matrix[99][372] * vector[99] +b[372];
assign result[373] = matrix[0][373] * vector[0] +matrix[1][373] * vector[1] +matrix[2][373] * vector[2] +matrix[3][373] * vector[3] +matrix[4][373] * vector[4] +matrix[5][373] * vector[5] +matrix[6][373] * vector[6] +matrix[7][373] * vector[7] +matrix[8][373] * vector[8] +matrix[9][373] * vector[9] +matrix[10][373] * vector[10] +matrix[11][373] * vector[11] +matrix[12][373] * vector[12] +matrix[13][373] * vector[13] +matrix[14][373] * vector[14] +matrix[15][373] * vector[15] +matrix[16][373] * vector[16] +matrix[17][373] * vector[17] +matrix[18][373] * vector[18] +matrix[19][373] * vector[19] +matrix[20][373] * vector[20] +matrix[21][373] * vector[21] +matrix[22][373] * vector[22] +matrix[23][373] * vector[23] +matrix[24][373] * vector[24] +matrix[25][373] * vector[25] +matrix[26][373] * vector[26] +matrix[27][373] * vector[27] +matrix[28][373] * vector[28] +matrix[29][373] * vector[29] +matrix[30][373] * vector[30] +matrix[31][373] * vector[31] +matrix[32][373] * vector[32] +matrix[33][373] * vector[33] +matrix[34][373] * vector[34] +matrix[35][373] * vector[35] +matrix[36][373] * vector[36] +matrix[37][373] * vector[37] +matrix[38][373] * vector[38] +matrix[39][373] * vector[39] +matrix[40][373] * vector[40] +matrix[41][373] * vector[41] +matrix[42][373] * vector[42] +matrix[43][373] * vector[43] +matrix[44][373] * vector[44] +matrix[45][373] * vector[45] +matrix[46][373] * vector[46] +matrix[47][373] * vector[47] +matrix[48][373] * vector[48] +matrix[49][373] * vector[49] +matrix[50][373] * vector[50] +matrix[51][373] * vector[51] +matrix[52][373] * vector[52] +matrix[53][373] * vector[53] +matrix[54][373] * vector[54] +matrix[55][373] * vector[55] +matrix[56][373] * vector[56] +matrix[57][373] * vector[57] +matrix[58][373] * vector[58] +matrix[59][373] * vector[59] +matrix[60][373] * vector[60] +matrix[61][373] * vector[61] +matrix[62][373] * vector[62] +matrix[63][373] * vector[63] +matrix[64][373] * vector[64] +matrix[65][373] * vector[65] +matrix[66][373] * vector[66] +matrix[67][373] * vector[67] +matrix[68][373] * vector[68] +matrix[69][373] * vector[69] +matrix[70][373] * vector[70] +matrix[71][373] * vector[71] +matrix[72][373] * vector[72] +matrix[73][373] * vector[73] +matrix[74][373] * vector[74] +matrix[75][373] * vector[75] +matrix[76][373] * vector[76] +matrix[77][373] * vector[77] +matrix[78][373] * vector[78] +matrix[79][373] * vector[79] +matrix[80][373] * vector[80] +matrix[81][373] * vector[81] +matrix[82][373] * vector[82] +matrix[83][373] * vector[83] +matrix[84][373] * vector[84] +matrix[85][373] * vector[85] +matrix[86][373] * vector[86] +matrix[87][373] * vector[87] +matrix[88][373] * vector[88] +matrix[89][373] * vector[89] +matrix[90][373] * vector[90] +matrix[91][373] * vector[91] +matrix[92][373] * vector[92] +matrix[93][373] * vector[93] +matrix[94][373] * vector[94] +matrix[95][373] * vector[95] +matrix[96][373] * vector[96] +matrix[97][373] * vector[97] +matrix[98][373] * vector[98] +matrix[99][373] * vector[99] +b[373];
assign result[374] = matrix[0][374] * vector[0] +matrix[1][374] * vector[1] +matrix[2][374] * vector[2] +matrix[3][374] * vector[3] +matrix[4][374] * vector[4] +matrix[5][374] * vector[5] +matrix[6][374] * vector[6] +matrix[7][374] * vector[7] +matrix[8][374] * vector[8] +matrix[9][374] * vector[9] +matrix[10][374] * vector[10] +matrix[11][374] * vector[11] +matrix[12][374] * vector[12] +matrix[13][374] * vector[13] +matrix[14][374] * vector[14] +matrix[15][374] * vector[15] +matrix[16][374] * vector[16] +matrix[17][374] * vector[17] +matrix[18][374] * vector[18] +matrix[19][374] * vector[19] +matrix[20][374] * vector[20] +matrix[21][374] * vector[21] +matrix[22][374] * vector[22] +matrix[23][374] * vector[23] +matrix[24][374] * vector[24] +matrix[25][374] * vector[25] +matrix[26][374] * vector[26] +matrix[27][374] * vector[27] +matrix[28][374] * vector[28] +matrix[29][374] * vector[29] +matrix[30][374] * vector[30] +matrix[31][374] * vector[31] +matrix[32][374] * vector[32] +matrix[33][374] * vector[33] +matrix[34][374] * vector[34] +matrix[35][374] * vector[35] +matrix[36][374] * vector[36] +matrix[37][374] * vector[37] +matrix[38][374] * vector[38] +matrix[39][374] * vector[39] +matrix[40][374] * vector[40] +matrix[41][374] * vector[41] +matrix[42][374] * vector[42] +matrix[43][374] * vector[43] +matrix[44][374] * vector[44] +matrix[45][374] * vector[45] +matrix[46][374] * vector[46] +matrix[47][374] * vector[47] +matrix[48][374] * vector[48] +matrix[49][374] * vector[49] +matrix[50][374] * vector[50] +matrix[51][374] * vector[51] +matrix[52][374] * vector[52] +matrix[53][374] * vector[53] +matrix[54][374] * vector[54] +matrix[55][374] * vector[55] +matrix[56][374] * vector[56] +matrix[57][374] * vector[57] +matrix[58][374] * vector[58] +matrix[59][374] * vector[59] +matrix[60][374] * vector[60] +matrix[61][374] * vector[61] +matrix[62][374] * vector[62] +matrix[63][374] * vector[63] +matrix[64][374] * vector[64] +matrix[65][374] * vector[65] +matrix[66][374] * vector[66] +matrix[67][374] * vector[67] +matrix[68][374] * vector[68] +matrix[69][374] * vector[69] +matrix[70][374] * vector[70] +matrix[71][374] * vector[71] +matrix[72][374] * vector[72] +matrix[73][374] * vector[73] +matrix[74][374] * vector[74] +matrix[75][374] * vector[75] +matrix[76][374] * vector[76] +matrix[77][374] * vector[77] +matrix[78][374] * vector[78] +matrix[79][374] * vector[79] +matrix[80][374] * vector[80] +matrix[81][374] * vector[81] +matrix[82][374] * vector[82] +matrix[83][374] * vector[83] +matrix[84][374] * vector[84] +matrix[85][374] * vector[85] +matrix[86][374] * vector[86] +matrix[87][374] * vector[87] +matrix[88][374] * vector[88] +matrix[89][374] * vector[89] +matrix[90][374] * vector[90] +matrix[91][374] * vector[91] +matrix[92][374] * vector[92] +matrix[93][374] * vector[93] +matrix[94][374] * vector[94] +matrix[95][374] * vector[95] +matrix[96][374] * vector[96] +matrix[97][374] * vector[97] +matrix[98][374] * vector[98] +matrix[99][374] * vector[99] +b[374];
assign result[375] = matrix[0][375] * vector[0] +matrix[1][375] * vector[1] +matrix[2][375] * vector[2] +matrix[3][375] * vector[3] +matrix[4][375] * vector[4] +matrix[5][375] * vector[5] +matrix[6][375] * vector[6] +matrix[7][375] * vector[7] +matrix[8][375] * vector[8] +matrix[9][375] * vector[9] +matrix[10][375] * vector[10] +matrix[11][375] * vector[11] +matrix[12][375] * vector[12] +matrix[13][375] * vector[13] +matrix[14][375] * vector[14] +matrix[15][375] * vector[15] +matrix[16][375] * vector[16] +matrix[17][375] * vector[17] +matrix[18][375] * vector[18] +matrix[19][375] * vector[19] +matrix[20][375] * vector[20] +matrix[21][375] * vector[21] +matrix[22][375] * vector[22] +matrix[23][375] * vector[23] +matrix[24][375] * vector[24] +matrix[25][375] * vector[25] +matrix[26][375] * vector[26] +matrix[27][375] * vector[27] +matrix[28][375] * vector[28] +matrix[29][375] * vector[29] +matrix[30][375] * vector[30] +matrix[31][375] * vector[31] +matrix[32][375] * vector[32] +matrix[33][375] * vector[33] +matrix[34][375] * vector[34] +matrix[35][375] * vector[35] +matrix[36][375] * vector[36] +matrix[37][375] * vector[37] +matrix[38][375] * vector[38] +matrix[39][375] * vector[39] +matrix[40][375] * vector[40] +matrix[41][375] * vector[41] +matrix[42][375] * vector[42] +matrix[43][375] * vector[43] +matrix[44][375] * vector[44] +matrix[45][375] * vector[45] +matrix[46][375] * vector[46] +matrix[47][375] * vector[47] +matrix[48][375] * vector[48] +matrix[49][375] * vector[49] +matrix[50][375] * vector[50] +matrix[51][375] * vector[51] +matrix[52][375] * vector[52] +matrix[53][375] * vector[53] +matrix[54][375] * vector[54] +matrix[55][375] * vector[55] +matrix[56][375] * vector[56] +matrix[57][375] * vector[57] +matrix[58][375] * vector[58] +matrix[59][375] * vector[59] +matrix[60][375] * vector[60] +matrix[61][375] * vector[61] +matrix[62][375] * vector[62] +matrix[63][375] * vector[63] +matrix[64][375] * vector[64] +matrix[65][375] * vector[65] +matrix[66][375] * vector[66] +matrix[67][375] * vector[67] +matrix[68][375] * vector[68] +matrix[69][375] * vector[69] +matrix[70][375] * vector[70] +matrix[71][375] * vector[71] +matrix[72][375] * vector[72] +matrix[73][375] * vector[73] +matrix[74][375] * vector[74] +matrix[75][375] * vector[75] +matrix[76][375] * vector[76] +matrix[77][375] * vector[77] +matrix[78][375] * vector[78] +matrix[79][375] * vector[79] +matrix[80][375] * vector[80] +matrix[81][375] * vector[81] +matrix[82][375] * vector[82] +matrix[83][375] * vector[83] +matrix[84][375] * vector[84] +matrix[85][375] * vector[85] +matrix[86][375] * vector[86] +matrix[87][375] * vector[87] +matrix[88][375] * vector[88] +matrix[89][375] * vector[89] +matrix[90][375] * vector[90] +matrix[91][375] * vector[91] +matrix[92][375] * vector[92] +matrix[93][375] * vector[93] +matrix[94][375] * vector[94] +matrix[95][375] * vector[95] +matrix[96][375] * vector[96] +matrix[97][375] * vector[97] +matrix[98][375] * vector[98] +matrix[99][375] * vector[99] +b[375];
assign result[376] = matrix[0][376] * vector[0] +matrix[1][376] * vector[1] +matrix[2][376] * vector[2] +matrix[3][376] * vector[3] +matrix[4][376] * vector[4] +matrix[5][376] * vector[5] +matrix[6][376] * vector[6] +matrix[7][376] * vector[7] +matrix[8][376] * vector[8] +matrix[9][376] * vector[9] +matrix[10][376] * vector[10] +matrix[11][376] * vector[11] +matrix[12][376] * vector[12] +matrix[13][376] * vector[13] +matrix[14][376] * vector[14] +matrix[15][376] * vector[15] +matrix[16][376] * vector[16] +matrix[17][376] * vector[17] +matrix[18][376] * vector[18] +matrix[19][376] * vector[19] +matrix[20][376] * vector[20] +matrix[21][376] * vector[21] +matrix[22][376] * vector[22] +matrix[23][376] * vector[23] +matrix[24][376] * vector[24] +matrix[25][376] * vector[25] +matrix[26][376] * vector[26] +matrix[27][376] * vector[27] +matrix[28][376] * vector[28] +matrix[29][376] * vector[29] +matrix[30][376] * vector[30] +matrix[31][376] * vector[31] +matrix[32][376] * vector[32] +matrix[33][376] * vector[33] +matrix[34][376] * vector[34] +matrix[35][376] * vector[35] +matrix[36][376] * vector[36] +matrix[37][376] * vector[37] +matrix[38][376] * vector[38] +matrix[39][376] * vector[39] +matrix[40][376] * vector[40] +matrix[41][376] * vector[41] +matrix[42][376] * vector[42] +matrix[43][376] * vector[43] +matrix[44][376] * vector[44] +matrix[45][376] * vector[45] +matrix[46][376] * vector[46] +matrix[47][376] * vector[47] +matrix[48][376] * vector[48] +matrix[49][376] * vector[49] +matrix[50][376] * vector[50] +matrix[51][376] * vector[51] +matrix[52][376] * vector[52] +matrix[53][376] * vector[53] +matrix[54][376] * vector[54] +matrix[55][376] * vector[55] +matrix[56][376] * vector[56] +matrix[57][376] * vector[57] +matrix[58][376] * vector[58] +matrix[59][376] * vector[59] +matrix[60][376] * vector[60] +matrix[61][376] * vector[61] +matrix[62][376] * vector[62] +matrix[63][376] * vector[63] +matrix[64][376] * vector[64] +matrix[65][376] * vector[65] +matrix[66][376] * vector[66] +matrix[67][376] * vector[67] +matrix[68][376] * vector[68] +matrix[69][376] * vector[69] +matrix[70][376] * vector[70] +matrix[71][376] * vector[71] +matrix[72][376] * vector[72] +matrix[73][376] * vector[73] +matrix[74][376] * vector[74] +matrix[75][376] * vector[75] +matrix[76][376] * vector[76] +matrix[77][376] * vector[77] +matrix[78][376] * vector[78] +matrix[79][376] * vector[79] +matrix[80][376] * vector[80] +matrix[81][376] * vector[81] +matrix[82][376] * vector[82] +matrix[83][376] * vector[83] +matrix[84][376] * vector[84] +matrix[85][376] * vector[85] +matrix[86][376] * vector[86] +matrix[87][376] * vector[87] +matrix[88][376] * vector[88] +matrix[89][376] * vector[89] +matrix[90][376] * vector[90] +matrix[91][376] * vector[91] +matrix[92][376] * vector[92] +matrix[93][376] * vector[93] +matrix[94][376] * vector[94] +matrix[95][376] * vector[95] +matrix[96][376] * vector[96] +matrix[97][376] * vector[97] +matrix[98][376] * vector[98] +matrix[99][376] * vector[99] +b[376];
assign result[377] = matrix[0][377] * vector[0] +matrix[1][377] * vector[1] +matrix[2][377] * vector[2] +matrix[3][377] * vector[3] +matrix[4][377] * vector[4] +matrix[5][377] * vector[5] +matrix[6][377] * vector[6] +matrix[7][377] * vector[7] +matrix[8][377] * vector[8] +matrix[9][377] * vector[9] +matrix[10][377] * vector[10] +matrix[11][377] * vector[11] +matrix[12][377] * vector[12] +matrix[13][377] * vector[13] +matrix[14][377] * vector[14] +matrix[15][377] * vector[15] +matrix[16][377] * vector[16] +matrix[17][377] * vector[17] +matrix[18][377] * vector[18] +matrix[19][377] * vector[19] +matrix[20][377] * vector[20] +matrix[21][377] * vector[21] +matrix[22][377] * vector[22] +matrix[23][377] * vector[23] +matrix[24][377] * vector[24] +matrix[25][377] * vector[25] +matrix[26][377] * vector[26] +matrix[27][377] * vector[27] +matrix[28][377] * vector[28] +matrix[29][377] * vector[29] +matrix[30][377] * vector[30] +matrix[31][377] * vector[31] +matrix[32][377] * vector[32] +matrix[33][377] * vector[33] +matrix[34][377] * vector[34] +matrix[35][377] * vector[35] +matrix[36][377] * vector[36] +matrix[37][377] * vector[37] +matrix[38][377] * vector[38] +matrix[39][377] * vector[39] +matrix[40][377] * vector[40] +matrix[41][377] * vector[41] +matrix[42][377] * vector[42] +matrix[43][377] * vector[43] +matrix[44][377] * vector[44] +matrix[45][377] * vector[45] +matrix[46][377] * vector[46] +matrix[47][377] * vector[47] +matrix[48][377] * vector[48] +matrix[49][377] * vector[49] +matrix[50][377] * vector[50] +matrix[51][377] * vector[51] +matrix[52][377] * vector[52] +matrix[53][377] * vector[53] +matrix[54][377] * vector[54] +matrix[55][377] * vector[55] +matrix[56][377] * vector[56] +matrix[57][377] * vector[57] +matrix[58][377] * vector[58] +matrix[59][377] * vector[59] +matrix[60][377] * vector[60] +matrix[61][377] * vector[61] +matrix[62][377] * vector[62] +matrix[63][377] * vector[63] +matrix[64][377] * vector[64] +matrix[65][377] * vector[65] +matrix[66][377] * vector[66] +matrix[67][377] * vector[67] +matrix[68][377] * vector[68] +matrix[69][377] * vector[69] +matrix[70][377] * vector[70] +matrix[71][377] * vector[71] +matrix[72][377] * vector[72] +matrix[73][377] * vector[73] +matrix[74][377] * vector[74] +matrix[75][377] * vector[75] +matrix[76][377] * vector[76] +matrix[77][377] * vector[77] +matrix[78][377] * vector[78] +matrix[79][377] * vector[79] +matrix[80][377] * vector[80] +matrix[81][377] * vector[81] +matrix[82][377] * vector[82] +matrix[83][377] * vector[83] +matrix[84][377] * vector[84] +matrix[85][377] * vector[85] +matrix[86][377] * vector[86] +matrix[87][377] * vector[87] +matrix[88][377] * vector[88] +matrix[89][377] * vector[89] +matrix[90][377] * vector[90] +matrix[91][377] * vector[91] +matrix[92][377] * vector[92] +matrix[93][377] * vector[93] +matrix[94][377] * vector[94] +matrix[95][377] * vector[95] +matrix[96][377] * vector[96] +matrix[97][377] * vector[97] +matrix[98][377] * vector[98] +matrix[99][377] * vector[99] +b[377];
assign result[378] = matrix[0][378] * vector[0] +matrix[1][378] * vector[1] +matrix[2][378] * vector[2] +matrix[3][378] * vector[3] +matrix[4][378] * vector[4] +matrix[5][378] * vector[5] +matrix[6][378] * vector[6] +matrix[7][378] * vector[7] +matrix[8][378] * vector[8] +matrix[9][378] * vector[9] +matrix[10][378] * vector[10] +matrix[11][378] * vector[11] +matrix[12][378] * vector[12] +matrix[13][378] * vector[13] +matrix[14][378] * vector[14] +matrix[15][378] * vector[15] +matrix[16][378] * vector[16] +matrix[17][378] * vector[17] +matrix[18][378] * vector[18] +matrix[19][378] * vector[19] +matrix[20][378] * vector[20] +matrix[21][378] * vector[21] +matrix[22][378] * vector[22] +matrix[23][378] * vector[23] +matrix[24][378] * vector[24] +matrix[25][378] * vector[25] +matrix[26][378] * vector[26] +matrix[27][378] * vector[27] +matrix[28][378] * vector[28] +matrix[29][378] * vector[29] +matrix[30][378] * vector[30] +matrix[31][378] * vector[31] +matrix[32][378] * vector[32] +matrix[33][378] * vector[33] +matrix[34][378] * vector[34] +matrix[35][378] * vector[35] +matrix[36][378] * vector[36] +matrix[37][378] * vector[37] +matrix[38][378] * vector[38] +matrix[39][378] * vector[39] +matrix[40][378] * vector[40] +matrix[41][378] * vector[41] +matrix[42][378] * vector[42] +matrix[43][378] * vector[43] +matrix[44][378] * vector[44] +matrix[45][378] * vector[45] +matrix[46][378] * vector[46] +matrix[47][378] * vector[47] +matrix[48][378] * vector[48] +matrix[49][378] * vector[49] +matrix[50][378] * vector[50] +matrix[51][378] * vector[51] +matrix[52][378] * vector[52] +matrix[53][378] * vector[53] +matrix[54][378] * vector[54] +matrix[55][378] * vector[55] +matrix[56][378] * vector[56] +matrix[57][378] * vector[57] +matrix[58][378] * vector[58] +matrix[59][378] * vector[59] +matrix[60][378] * vector[60] +matrix[61][378] * vector[61] +matrix[62][378] * vector[62] +matrix[63][378] * vector[63] +matrix[64][378] * vector[64] +matrix[65][378] * vector[65] +matrix[66][378] * vector[66] +matrix[67][378] * vector[67] +matrix[68][378] * vector[68] +matrix[69][378] * vector[69] +matrix[70][378] * vector[70] +matrix[71][378] * vector[71] +matrix[72][378] * vector[72] +matrix[73][378] * vector[73] +matrix[74][378] * vector[74] +matrix[75][378] * vector[75] +matrix[76][378] * vector[76] +matrix[77][378] * vector[77] +matrix[78][378] * vector[78] +matrix[79][378] * vector[79] +matrix[80][378] * vector[80] +matrix[81][378] * vector[81] +matrix[82][378] * vector[82] +matrix[83][378] * vector[83] +matrix[84][378] * vector[84] +matrix[85][378] * vector[85] +matrix[86][378] * vector[86] +matrix[87][378] * vector[87] +matrix[88][378] * vector[88] +matrix[89][378] * vector[89] +matrix[90][378] * vector[90] +matrix[91][378] * vector[91] +matrix[92][378] * vector[92] +matrix[93][378] * vector[93] +matrix[94][378] * vector[94] +matrix[95][378] * vector[95] +matrix[96][378] * vector[96] +matrix[97][378] * vector[97] +matrix[98][378] * vector[98] +matrix[99][378] * vector[99] +b[378];
assign result[379] = matrix[0][379] * vector[0] +matrix[1][379] * vector[1] +matrix[2][379] * vector[2] +matrix[3][379] * vector[3] +matrix[4][379] * vector[4] +matrix[5][379] * vector[5] +matrix[6][379] * vector[6] +matrix[7][379] * vector[7] +matrix[8][379] * vector[8] +matrix[9][379] * vector[9] +matrix[10][379] * vector[10] +matrix[11][379] * vector[11] +matrix[12][379] * vector[12] +matrix[13][379] * vector[13] +matrix[14][379] * vector[14] +matrix[15][379] * vector[15] +matrix[16][379] * vector[16] +matrix[17][379] * vector[17] +matrix[18][379] * vector[18] +matrix[19][379] * vector[19] +matrix[20][379] * vector[20] +matrix[21][379] * vector[21] +matrix[22][379] * vector[22] +matrix[23][379] * vector[23] +matrix[24][379] * vector[24] +matrix[25][379] * vector[25] +matrix[26][379] * vector[26] +matrix[27][379] * vector[27] +matrix[28][379] * vector[28] +matrix[29][379] * vector[29] +matrix[30][379] * vector[30] +matrix[31][379] * vector[31] +matrix[32][379] * vector[32] +matrix[33][379] * vector[33] +matrix[34][379] * vector[34] +matrix[35][379] * vector[35] +matrix[36][379] * vector[36] +matrix[37][379] * vector[37] +matrix[38][379] * vector[38] +matrix[39][379] * vector[39] +matrix[40][379] * vector[40] +matrix[41][379] * vector[41] +matrix[42][379] * vector[42] +matrix[43][379] * vector[43] +matrix[44][379] * vector[44] +matrix[45][379] * vector[45] +matrix[46][379] * vector[46] +matrix[47][379] * vector[47] +matrix[48][379] * vector[48] +matrix[49][379] * vector[49] +matrix[50][379] * vector[50] +matrix[51][379] * vector[51] +matrix[52][379] * vector[52] +matrix[53][379] * vector[53] +matrix[54][379] * vector[54] +matrix[55][379] * vector[55] +matrix[56][379] * vector[56] +matrix[57][379] * vector[57] +matrix[58][379] * vector[58] +matrix[59][379] * vector[59] +matrix[60][379] * vector[60] +matrix[61][379] * vector[61] +matrix[62][379] * vector[62] +matrix[63][379] * vector[63] +matrix[64][379] * vector[64] +matrix[65][379] * vector[65] +matrix[66][379] * vector[66] +matrix[67][379] * vector[67] +matrix[68][379] * vector[68] +matrix[69][379] * vector[69] +matrix[70][379] * vector[70] +matrix[71][379] * vector[71] +matrix[72][379] * vector[72] +matrix[73][379] * vector[73] +matrix[74][379] * vector[74] +matrix[75][379] * vector[75] +matrix[76][379] * vector[76] +matrix[77][379] * vector[77] +matrix[78][379] * vector[78] +matrix[79][379] * vector[79] +matrix[80][379] * vector[80] +matrix[81][379] * vector[81] +matrix[82][379] * vector[82] +matrix[83][379] * vector[83] +matrix[84][379] * vector[84] +matrix[85][379] * vector[85] +matrix[86][379] * vector[86] +matrix[87][379] * vector[87] +matrix[88][379] * vector[88] +matrix[89][379] * vector[89] +matrix[90][379] * vector[90] +matrix[91][379] * vector[91] +matrix[92][379] * vector[92] +matrix[93][379] * vector[93] +matrix[94][379] * vector[94] +matrix[95][379] * vector[95] +matrix[96][379] * vector[96] +matrix[97][379] * vector[97] +matrix[98][379] * vector[98] +matrix[99][379] * vector[99] +b[379];
assign result[380] = matrix[0][380] * vector[0] +matrix[1][380] * vector[1] +matrix[2][380] * vector[2] +matrix[3][380] * vector[3] +matrix[4][380] * vector[4] +matrix[5][380] * vector[5] +matrix[6][380] * vector[6] +matrix[7][380] * vector[7] +matrix[8][380] * vector[8] +matrix[9][380] * vector[9] +matrix[10][380] * vector[10] +matrix[11][380] * vector[11] +matrix[12][380] * vector[12] +matrix[13][380] * vector[13] +matrix[14][380] * vector[14] +matrix[15][380] * vector[15] +matrix[16][380] * vector[16] +matrix[17][380] * vector[17] +matrix[18][380] * vector[18] +matrix[19][380] * vector[19] +matrix[20][380] * vector[20] +matrix[21][380] * vector[21] +matrix[22][380] * vector[22] +matrix[23][380] * vector[23] +matrix[24][380] * vector[24] +matrix[25][380] * vector[25] +matrix[26][380] * vector[26] +matrix[27][380] * vector[27] +matrix[28][380] * vector[28] +matrix[29][380] * vector[29] +matrix[30][380] * vector[30] +matrix[31][380] * vector[31] +matrix[32][380] * vector[32] +matrix[33][380] * vector[33] +matrix[34][380] * vector[34] +matrix[35][380] * vector[35] +matrix[36][380] * vector[36] +matrix[37][380] * vector[37] +matrix[38][380] * vector[38] +matrix[39][380] * vector[39] +matrix[40][380] * vector[40] +matrix[41][380] * vector[41] +matrix[42][380] * vector[42] +matrix[43][380] * vector[43] +matrix[44][380] * vector[44] +matrix[45][380] * vector[45] +matrix[46][380] * vector[46] +matrix[47][380] * vector[47] +matrix[48][380] * vector[48] +matrix[49][380] * vector[49] +matrix[50][380] * vector[50] +matrix[51][380] * vector[51] +matrix[52][380] * vector[52] +matrix[53][380] * vector[53] +matrix[54][380] * vector[54] +matrix[55][380] * vector[55] +matrix[56][380] * vector[56] +matrix[57][380] * vector[57] +matrix[58][380] * vector[58] +matrix[59][380] * vector[59] +matrix[60][380] * vector[60] +matrix[61][380] * vector[61] +matrix[62][380] * vector[62] +matrix[63][380] * vector[63] +matrix[64][380] * vector[64] +matrix[65][380] * vector[65] +matrix[66][380] * vector[66] +matrix[67][380] * vector[67] +matrix[68][380] * vector[68] +matrix[69][380] * vector[69] +matrix[70][380] * vector[70] +matrix[71][380] * vector[71] +matrix[72][380] * vector[72] +matrix[73][380] * vector[73] +matrix[74][380] * vector[74] +matrix[75][380] * vector[75] +matrix[76][380] * vector[76] +matrix[77][380] * vector[77] +matrix[78][380] * vector[78] +matrix[79][380] * vector[79] +matrix[80][380] * vector[80] +matrix[81][380] * vector[81] +matrix[82][380] * vector[82] +matrix[83][380] * vector[83] +matrix[84][380] * vector[84] +matrix[85][380] * vector[85] +matrix[86][380] * vector[86] +matrix[87][380] * vector[87] +matrix[88][380] * vector[88] +matrix[89][380] * vector[89] +matrix[90][380] * vector[90] +matrix[91][380] * vector[91] +matrix[92][380] * vector[92] +matrix[93][380] * vector[93] +matrix[94][380] * vector[94] +matrix[95][380] * vector[95] +matrix[96][380] * vector[96] +matrix[97][380] * vector[97] +matrix[98][380] * vector[98] +matrix[99][380] * vector[99] +b[380];
assign result[381] = matrix[0][381] * vector[0] +matrix[1][381] * vector[1] +matrix[2][381] * vector[2] +matrix[3][381] * vector[3] +matrix[4][381] * vector[4] +matrix[5][381] * vector[5] +matrix[6][381] * vector[6] +matrix[7][381] * vector[7] +matrix[8][381] * vector[8] +matrix[9][381] * vector[9] +matrix[10][381] * vector[10] +matrix[11][381] * vector[11] +matrix[12][381] * vector[12] +matrix[13][381] * vector[13] +matrix[14][381] * vector[14] +matrix[15][381] * vector[15] +matrix[16][381] * vector[16] +matrix[17][381] * vector[17] +matrix[18][381] * vector[18] +matrix[19][381] * vector[19] +matrix[20][381] * vector[20] +matrix[21][381] * vector[21] +matrix[22][381] * vector[22] +matrix[23][381] * vector[23] +matrix[24][381] * vector[24] +matrix[25][381] * vector[25] +matrix[26][381] * vector[26] +matrix[27][381] * vector[27] +matrix[28][381] * vector[28] +matrix[29][381] * vector[29] +matrix[30][381] * vector[30] +matrix[31][381] * vector[31] +matrix[32][381] * vector[32] +matrix[33][381] * vector[33] +matrix[34][381] * vector[34] +matrix[35][381] * vector[35] +matrix[36][381] * vector[36] +matrix[37][381] * vector[37] +matrix[38][381] * vector[38] +matrix[39][381] * vector[39] +matrix[40][381] * vector[40] +matrix[41][381] * vector[41] +matrix[42][381] * vector[42] +matrix[43][381] * vector[43] +matrix[44][381] * vector[44] +matrix[45][381] * vector[45] +matrix[46][381] * vector[46] +matrix[47][381] * vector[47] +matrix[48][381] * vector[48] +matrix[49][381] * vector[49] +matrix[50][381] * vector[50] +matrix[51][381] * vector[51] +matrix[52][381] * vector[52] +matrix[53][381] * vector[53] +matrix[54][381] * vector[54] +matrix[55][381] * vector[55] +matrix[56][381] * vector[56] +matrix[57][381] * vector[57] +matrix[58][381] * vector[58] +matrix[59][381] * vector[59] +matrix[60][381] * vector[60] +matrix[61][381] * vector[61] +matrix[62][381] * vector[62] +matrix[63][381] * vector[63] +matrix[64][381] * vector[64] +matrix[65][381] * vector[65] +matrix[66][381] * vector[66] +matrix[67][381] * vector[67] +matrix[68][381] * vector[68] +matrix[69][381] * vector[69] +matrix[70][381] * vector[70] +matrix[71][381] * vector[71] +matrix[72][381] * vector[72] +matrix[73][381] * vector[73] +matrix[74][381] * vector[74] +matrix[75][381] * vector[75] +matrix[76][381] * vector[76] +matrix[77][381] * vector[77] +matrix[78][381] * vector[78] +matrix[79][381] * vector[79] +matrix[80][381] * vector[80] +matrix[81][381] * vector[81] +matrix[82][381] * vector[82] +matrix[83][381] * vector[83] +matrix[84][381] * vector[84] +matrix[85][381] * vector[85] +matrix[86][381] * vector[86] +matrix[87][381] * vector[87] +matrix[88][381] * vector[88] +matrix[89][381] * vector[89] +matrix[90][381] * vector[90] +matrix[91][381] * vector[91] +matrix[92][381] * vector[92] +matrix[93][381] * vector[93] +matrix[94][381] * vector[94] +matrix[95][381] * vector[95] +matrix[96][381] * vector[96] +matrix[97][381] * vector[97] +matrix[98][381] * vector[98] +matrix[99][381] * vector[99] +b[381];
assign result[382] = matrix[0][382] * vector[0] +matrix[1][382] * vector[1] +matrix[2][382] * vector[2] +matrix[3][382] * vector[3] +matrix[4][382] * vector[4] +matrix[5][382] * vector[5] +matrix[6][382] * vector[6] +matrix[7][382] * vector[7] +matrix[8][382] * vector[8] +matrix[9][382] * vector[9] +matrix[10][382] * vector[10] +matrix[11][382] * vector[11] +matrix[12][382] * vector[12] +matrix[13][382] * vector[13] +matrix[14][382] * vector[14] +matrix[15][382] * vector[15] +matrix[16][382] * vector[16] +matrix[17][382] * vector[17] +matrix[18][382] * vector[18] +matrix[19][382] * vector[19] +matrix[20][382] * vector[20] +matrix[21][382] * vector[21] +matrix[22][382] * vector[22] +matrix[23][382] * vector[23] +matrix[24][382] * vector[24] +matrix[25][382] * vector[25] +matrix[26][382] * vector[26] +matrix[27][382] * vector[27] +matrix[28][382] * vector[28] +matrix[29][382] * vector[29] +matrix[30][382] * vector[30] +matrix[31][382] * vector[31] +matrix[32][382] * vector[32] +matrix[33][382] * vector[33] +matrix[34][382] * vector[34] +matrix[35][382] * vector[35] +matrix[36][382] * vector[36] +matrix[37][382] * vector[37] +matrix[38][382] * vector[38] +matrix[39][382] * vector[39] +matrix[40][382] * vector[40] +matrix[41][382] * vector[41] +matrix[42][382] * vector[42] +matrix[43][382] * vector[43] +matrix[44][382] * vector[44] +matrix[45][382] * vector[45] +matrix[46][382] * vector[46] +matrix[47][382] * vector[47] +matrix[48][382] * vector[48] +matrix[49][382] * vector[49] +matrix[50][382] * vector[50] +matrix[51][382] * vector[51] +matrix[52][382] * vector[52] +matrix[53][382] * vector[53] +matrix[54][382] * vector[54] +matrix[55][382] * vector[55] +matrix[56][382] * vector[56] +matrix[57][382] * vector[57] +matrix[58][382] * vector[58] +matrix[59][382] * vector[59] +matrix[60][382] * vector[60] +matrix[61][382] * vector[61] +matrix[62][382] * vector[62] +matrix[63][382] * vector[63] +matrix[64][382] * vector[64] +matrix[65][382] * vector[65] +matrix[66][382] * vector[66] +matrix[67][382] * vector[67] +matrix[68][382] * vector[68] +matrix[69][382] * vector[69] +matrix[70][382] * vector[70] +matrix[71][382] * vector[71] +matrix[72][382] * vector[72] +matrix[73][382] * vector[73] +matrix[74][382] * vector[74] +matrix[75][382] * vector[75] +matrix[76][382] * vector[76] +matrix[77][382] * vector[77] +matrix[78][382] * vector[78] +matrix[79][382] * vector[79] +matrix[80][382] * vector[80] +matrix[81][382] * vector[81] +matrix[82][382] * vector[82] +matrix[83][382] * vector[83] +matrix[84][382] * vector[84] +matrix[85][382] * vector[85] +matrix[86][382] * vector[86] +matrix[87][382] * vector[87] +matrix[88][382] * vector[88] +matrix[89][382] * vector[89] +matrix[90][382] * vector[90] +matrix[91][382] * vector[91] +matrix[92][382] * vector[92] +matrix[93][382] * vector[93] +matrix[94][382] * vector[94] +matrix[95][382] * vector[95] +matrix[96][382] * vector[96] +matrix[97][382] * vector[97] +matrix[98][382] * vector[98] +matrix[99][382] * vector[99] +b[382];
assign result[383] = matrix[0][383] * vector[0] +matrix[1][383] * vector[1] +matrix[2][383] * vector[2] +matrix[3][383] * vector[3] +matrix[4][383] * vector[4] +matrix[5][383] * vector[5] +matrix[6][383] * vector[6] +matrix[7][383] * vector[7] +matrix[8][383] * vector[8] +matrix[9][383] * vector[9] +matrix[10][383] * vector[10] +matrix[11][383] * vector[11] +matrix[12][383] * vector[12] +matrix[13][383] * vector[13] +matrix[14][383] * vector[14] +matrix[15][383] * vector[15] +matrix[16][383] * vector[16] +matrix[17][383] * vector[17] +matrix[18][383] * vector[18] +matrix[19][383] * vector[19] +matrix[20][383] * vector[20] +matrix[21][383] * vector[21] +matrix[22][383] * vector[22] +matrix[23][383] * vector[23] +matrix[24][383] * vector[24] +matrix[25][383] * vector[25] +matrix[26][383] * vector[26] +matrix[27][383] * vector[27] +matrix[28][383] * vector[28] +matrix[29][383] * vector[29] +matrix[30][383] * vector[30] +matrix[31][383] * vector[31] +matrix[32][383] * vector[32] +matrix[33][383] * vector[33] +matrix[34][383] * vector[34] +matrix[35][383] * vector[35] +matrix[36][383] * vector[36] +matrix[37][383] * vector[37] +matrix[38][383] * vector[38] +matrix[39][383] * vector[39] +matrix[40][383] * vector[40] +matrix[41][383] * vector[41] +matrix[42][383] * vector[42] +matrix[43][383] * vector[43] +matrix[44][383] * vector[44] +matrix[45][383] * vector[45] +matrix[46][383] * vector[46] +matrix[47][383] * vector[47] +matrix[48][383] * vector[48] +matrix[49][383] * vector[49] +matrix[50][383] * vector[50] +matrix[51][383] * vector[51] +matrix[52][383] * vector[52] +matrix[53][383] * vector[53] +matrix[54][383] * vector[54] +matrix[55][383] * vector[55] +matrix[56][383] * vector[56] +matrix[57][383] * vector[57] +matrix[58][383] * vector[58] +matrix[59][383] * vector[59] +matrix[60][383] * vector[60] +matrix[61][383] * vector[61] +matrix[62][383] * vector[62] +matrix[63][383] * vector[63] +matrix[64][383] * vector[64] +matrix[65][383] * vector[65] +matrix[66][383] * vector[66] +matrix[67][383] * vector[67] +matrix[68][383] * vector[68] +matrix[69][383] * vector[69] +matrix[70][383] * vector[70] +matrix[71][383] * vector[71] +matrix[72][383] * vector[72] +matrix[73][383] * vector[73] +matrix[74][383] * vector[74] +matrix[75][383] * vector[75] +matrix[76][383] * vector[76] +matrix[77][383] * vector[77] +matrix[78][383] * vector[78] +matrix[79][383] * vector[79] +matrix[80][383] * vector[80] +matrix[81][383] * vector[81] +matrix[82][383] * vector[82] +matrix[83][383] * vector[83] +matrix[84][383] * vector[84] +matrix[85][383] * vector[85] +matrix[86][383] * vector[86] +matrix[87][383] * vector[87] +matrix[88][383] * vector[88] +matrix[89][383] * vector[89] +matrix[90][383] * vector[90] +matrix[91][383] * vector[91] +matrix[92][383] * vector[92] +matrix[93][383] * vector[93] +matrix[94][383] * vector[94] +matrix[95][383] * vector[95] +matrix[96][383] * vector[96] +matrix[97][383] * vector[97] +matrix[98][383] * vector[98] +matrix[99][383] * vector[99] +b[383];
assign result[384] = matrix[0][384] * vector[0] +matrix[1][384] * vector[1] +matrix[2][384] * vector[2] +matrix[3][384] * vector[3] +matrix[4][384] * vector[4] +matrix[5][384] * vector[5] +matrix[6][384] * vector[6] +matrix[7][384] * vector[7] +matrix[8][384] * vector[8] +matrix[9][384] * vector[9] +matrix[10][384] * vector[10] +matrix[11][384] * vector[11] +matrix[12][384] * vector[12] +matrix[13][384] * vector[13] +matrix[14][384] * vector[14] +matrix[15][384] * vector[15] +matrix[16][384] * vector[16] +matrix[17][384] * vector[17] +matrix[18][384] * vector[18] +matrix[19][384] * vector[19] +matrix[20][384] * vector[20] +matrix[21][384] * vector[21] +matrix[22][384] * vector[22] +matrix[23][384] * vector[23] +matrix[24][384] * vector[24] +matrix[25][384] * vector[25] +matrix[26][384] * vector[26] +matrix[27][384] * vector[27] +matrix[28][384] * vector[28] +matrix[29][384] * vector[29] +matrix[30][384] * vector[30] +matrix[31][384] * vector[31] +matrix[32][384] * vector[32] +matrix[33][384] * vector[33] +matrix[34][384] * vector[34] +matrix[35][384] * vector[35] +matrix[36][384] * vector[36] +matrix[37][384] * vector[37] +matrix[38][384] * vector[38] +matrix[39][384] * vector[39] +matrix[40][384] * vector[40] +matrix[41][384] * vector[41] +matrix[42][384] * vector[42] +matrix[43][384] * vector[43] +matrix[44][384] * vector[44] +matrix[45][384] * vector[45] +matrix[46][384] * vector[46] +matrix[47][384] * vector[47] +matrix[48][384] * vector[48] +matrix[49][384] * vector[49] +matrix[50][384] * vector[50] +matrix[51][384] * vector[51] +matrix[52][384] * vector[52] +matrix[53][384] * vector[53] +matrix[54][384] * vector[54] +matrix[55][384] * vector[55] +matrix[56][384] * vector[56] +matrix[57][384] * vector[57] +matrix[58][384] * vector[58] +matrix[59][384] * vector[59] +matrix[60][384] * vector[60] +matrix[61][384] * vector[61] +matrix[62][384] * vector[62] +matrix[63][384] * vector[63] +matrix[64][384] * vector[64] +matrix[65][384] * vector[65] +matrix[66][384] * vector[66] +matrix[67][384] * vector[67] +matrix[68][384] * vector[68] +matrix[69][384] * vector[69] +matrix[70][384] * vector[70] +matrix[71][384] * vector[71] +matrix[72][384] * vector[72] +matrix[73][384] * vector[73] +matrix[74][384] * vector[74] +matrix[75][384] * vector[75] +matrix[76][384] * vector[76] +matrix[77][384] * vector[77] +matrix[78][384] * vector[78] +matrix[79][384] * vector[79] +matrix[80][384] * vector[80] +matrix[81][384] * vector[81] +matrix[82][384] * vector[82] +matrix[83][384] * vector[83] +matrix[84][384] * vector[84] +matrix[85][384] * vector[85] +matrix[86][384] * vector[86] +matrix[87][384] * vector[87] +matrix[88][384] * vector[88] +matrix[89][384] * vector[89] +matrix[90][384] * vector[90] +matrix[91][384] * vector[91] +matrix[92][384] * vector[92] +matrix[93][384] * vector[93] +matrix[94][384] * vector[94] +matrix[95][384] * vector[95] +matrix[96][384] * vector[96] +matrix[97][384] * vector[97] +matrix[98][384] * vector[98] +matrix[99][384] * vector[99] +b[384];
assign result[385] = matrix[0][385] * vector[0] +matrix[1][385] * vector[1] +matrix[2][385] * vector[2] +matrix[3][385] * vector[3] +matrix[4][385] * vector[4] +matrix[5][385] * vector[5] +matrix[6][385] * vector[6] +matrix[7][385] * vector[7] +matrix[8][385] * vector[8] +matrix[9][385] * vector[9] +matrix[10][385] * vector[10] +matrix[11][385] * vector[11] +matrix[12][385] * vector[12] +matrix[13][385] * vector[13] +matrix[14][385] * vector[14] +matrix[15][385] * vector[15] +matrix[16][385] * vector[16] +matrix[17][385] * vector[17] +matrix[18][385] * vector[18] +matrix[19][385] * vector[19] +matrix[20][385] * vector[20] +matrix[21][385] * vector[21] +matrix[22][385] * vector[22] +matrix[23][385] * vector[23] +matrix[24][385] * vector[24] +matrix[25][385] * vector[25] +matrix[26][385] * vector[26] +matrix[27][385] * vector[27] +matrix[28][385] * vector[28] +matrix[29][385] * vector[29] +matrix[30][385] * vector[30] +matrix[31][385] * vector[31] +matrix[32][385] * vector[32] +matrix[33][385] * vector[33] +matrix[34][385] * vector[34] +matrix[35][385] * vector[35] +matrix[36][385] * vector[36] +matrix[37][385] * vector[37] +matrix[38][385] * vector[38] +matrix[39][385] * vector[39] +matrix[40][385] * vector[40] +matrix[41][385] * vector[41] +matrix[42][385] * vector[42] +matrix[43][385] * vector[43] +matrix[44][385] * vector[44] +matrix[45][385] * vector[45] +matrix[46][385] * vector[46] +matrix[47][385] * vector[47] +matrix[48][385] * vector[48] +matrix[49][385] * vector[49] +matrix[50][385] * vector[50] +matrix[51][385] * vector[51] +matrix[52][385] * vector[52] +matrix[53][385] * vector[53] +matrix[54][385] * vector[54] +matrix[55][385] * vector[55] +matrix[56][385] * vector[56] +matrix[57][385] * vector[57] +matrix[58][385] * vector[58] +matrix[59][385] * vector[59] +matrix[60][385] * vector[60] +matrix[61][385] * vector[61] +matrix[62][385] * vector[62] +matrix[63][385] * vector[63] +matrix[64][385] * vector[64] +matrix[65][385] * vector[65] +matrix[66][385] * vector[66] +matrix[67][385] * vector[67] +matrix[68][385] * vector[68] +matrix[69][385] * vector[69] +matrix[70][385] * vector[70] +matrix[71][385] * vector[71] +matrix[72][385] * vector[72] +matrix[73][385] * vector[73] +matrix[74][385] * vector[74] +matrix[75][385] * vector[75] +matrix[76][385] * vector[76] +matrix[77][385] * vector[77] +matrix[78][385] * vector[78] +matrix[79][385] * vector[79] +matrix[80][385] * vector[80] +matrix[81][385] * vector[81] +matrix[82][385] * vector[82] +matrix[83][385] * vector[83] +matrix[84][385] * vector[84] +matrix[85][385] * vector[85] +matrix[86][385] * vector[86] +matrix[87][385] * vector[87] +matrix[88][385] * vector[88] +matrix[89][385] * vector[89] +matrix[90][385] * vector[90] +matrix[91][385] * vector[91] +matrix[92][385] * vector[92] +matrix[93][385] * vector[93] +matrix[94][385] * vector[94] +matrix[95][385] * vector[95] +matrix[96][385] * vector[96] +matrix[97][385] * vector[97] +matrix[98][385] * vector[98] +matrix[99][385] * vector[99] +b[385];
assign result[386] = matrix[0][386] * vector[0] +matrix[1][386] * vector[1] +matrix[2][386] * vector[2] +matrix[3][386] * vector[3] +matrix[4][386] * vector[4] +matrix[5][386] * vector[5] +matrix[6][386] * vector[6] +matrix[7][386] * vector[7] +matrix[8][386] * vector[8] +matrix[9][386] * vector[9] +matrix[10][386] * vector[10] +matrix[11][386] * vector[11] +matrix[12][386] * vector[12] +matrix[13][386] * vector[13] +matrix[14][386] * vector[14] +matrix[15][386] * vector[15] +matrix[16][386] * vector[16] +matrix[17][386] * vector[17] +matrix[18][386] * vector[18] +matrix[19][386] * vector[19] +matrix[20][386] * vector[20] +matrix[21][386] * vector[21] +matrix[22][386] * vector[22] +matrix[23][386] * vector[23] +matrix[24][386] * vector[24] +matrix[25][386] * vector[25] +matrix[26][386] * vector[26] +matrix[27][386] * vector[27] +matrix[28][386] * vector[28] +matrix[29][386] * vector[29] +matrix[30][386] * vector[30] +matrix[31][386] * vector[31] +matrix[32][386] * vector[32] +matrix[33][386] * vector[33] +matrix[34][386] * vector[34] +matrix[35][386] * vector[35] +matrix[36][386] * vector[36] +matrix[37][386] * vector[37] +matrix[38][386] * vector[38] +matrix[39][386] * vector[39] +matrix[40][386] * vector[40] +matrix[41][386] * vector[41] +matrix[42][386] * vector[42] +matrix[43][386] * vector[43] +matrix[44][386] * vector[44] +matrix[45][386] * vector[45] +matrix[46][386] * vector[46] +matrix[47][386] * vector[47] +matrix[48][386] * vector[48] +matrix[49][386] * vector[49] +matrix[50][386] * vector[50] +matrix[51][386] * vector[51] +matrix[52][386] * vector[52] +matrix[53][386] * vector[53] +matrix[54][386] * vector[54] +matrix[55][386] * vector[55] +matrix[56][386] * vector[56] +matrix[57][386] * vector[57] +matrix[58][386] * vector[58] +matrix[59][386] * vector[59] +matrix[60][386] * vector[60] +matrix[61][386] * vector[61] +matrix[62][386] * vector[62] +matrix[63][386] * vector[63] +matrix[64][386] * vector[64] +matrix[65][386] * vector[65] +matrix[66][386] * vector[66] +matrix[67][386] * vector[67] +matrix[68][386] * vector[68] +matrix[69][386] * vector[69] +matrix[70][386] * vector[70] +matrix[71][386] * vector[71] +matrix[72][386] * vector[72] +matrix[73][386] * vector[73] +matrix[74][386] * vector[74] +matrix[75][386] * vector[75] +matrix[76][386] * vector[76] +matrix[77][386] * vector[77] +matrix[78][386] * vector[78] +matrix[79][386] * vector[79] +matrix[80][386] * vector[80] +matrix[81][386] * vector[81] +matrix[82][386] * vector[82] +matrix[83][386] * vector[83] +matrix[84][386] * vector[84] +matrix[85][386] * vector[85] +matrix[86][386] * vector[86] +matrix[87][386] * vector[87] +matrix[88][386] * vector[88] +matrix[89][386] * vector[89] +matrix[90][386] * vector[90] +matrix[91][386] * vector[91] +matrix[92][386] * vector[92] +matrix[93][386] * vector[93] +matrix[94][386] * vector[94] +matrix[95][386] * vector[95] +matrix[96][386] * vector[96] +matrix[97][386] * vector[97] +matrix[98][386] * vector[98] +matrix[99][386] * vector[99] +b[386];
assign result[387] = matrix[0][387] * vector[0] +matrix[1][387] * vector[1] +matrix[2][387] * vector[2] +matrix[3][387] * vector[3] +matrix[4][387] * vector[4] +matrix[5][387] * vector[5] +matrix[6][387] * vector[6] +matrix[7][387] * vector[7] +matrix[8][387] * vector[8] +matrix[9][387] * vector[9] +matrix[10][387] * vector[10] +matrix[11][387] * vector[11] +matrix[12][387] * vector[12] +matrix[13][387] * vector[13] +matrix[14][387] * vector[14] +matrix[15][387] * vector[15] +matrix[16][387] * vector[16] +matrix[17][387] * vector[17] +matrix[18][387] * vector[18] +matrix[19][387] * vector[19] +matrix[20][387] * vector[20] +matrix[21][387] * vector[21] +matrix[22][387] * vector[22] +matrix[23][387] * vector[23] +matrix[24][387] * vector[24] +matrix[25][387] * vector[25] +matrix[26][387] * vector[26] +matrix[27][387] * vector[27] +matrix[28][387] * vector[28] +matrix[29][387] * vector[29] +matrix[30][387] * vector[30] +matrix[31][387] * vector[31] +matrix[32][387] * vector[32] +matrix[33][387] * vector[33] +matrix[34][387] * vector[34] +matrix[35][387] * vector[35] +matrix[36][387] * vector[36] +matrix[37][387] * vector[37] +matrix[38][387] * vector[38] +matrix[39][387] * vector[39] +matrix[40][387] * vector[40] +matrix[41][387] * vector[41] +matrix[42][387] * vector[42] +matrix[43][387] * vector[43] +matrix[44][387] * vector[44] +matrix[45][387] * vector[45] +matrix[46][387] * vector[46] +matrix[47][387] * vector[47] +matrix[48][387] * vector[48] +matrix[49][387] * vector[49] +matrix[50][387] * vector[50] +matrix[51][387] * vector[51] +matrix[52][387] * vector[52] +matrix[53][387] * vector[53] +matrix[54][387] * vector[54] +matrix[55][387] * vector[55] +matrix[56][387] * vector[56] +matrix[57][387] * vector[57] +matrix[58][387] * vector[58] +matrix[59][387] * vector[59] +matrix[60][387] * vector[60] +matrix[61][387] * vector[61] +matrix[62][387] * vector[62] +matrix[63][387] * vector[63] +matrix[64][387] * vector[64] +matrix[65][387] * vector[65] +matrix[66][387] * vector[66] +matrix[67][387] * vector[67] +matrix[68][387] * vector[68] +matrix[69][387] * vector[69] +matrix[70][387] * vector[70] +matrix[71][387] * vector[71] +matrix[72][387] * vector[72] +matrix[73][387] * vector[73] +matrix[74][387] * vector[74] +matrix[75][387] * vector[75] +matrix[76][387] * vector[76] +matrix[77][387] * vector[77] +matrix[78][387] * vector[78] +matrix[79][387] * vector[79] +matrix[80][387] * vector[80] +matrix[81][387] * vector[81] +matrix[82][387] * vector[82] +matrix[83][387] * vector[83] +matrix[84][387] * vector[84] +matrix[85][387] * vector[85] +matrix[86][387] * vector[86] +matrix[87][387] * vector[87] +matrix[88][387] * vector[88] +matrix[89][387] * vector[89] +matrix[90][387] * vector[90] +matrix[91][387] * vector[91] +matrix[92][387] * vector[92] +matrix[93][387] * vector[93] +matrix[94][387] * vector[94] +matrix[95][387] * vector[95] +matrix[96][387] * vector[96] +matrix[97][387] * vector[97] +matrix[98][387] * vector[98] +matrix[99][387] * vector[99] +b[387];
assign result[388] = matrix[0][388] * vector[0] +matrix[1][388] * vector[1] +matrix[2][388] * vector[2] +matrix[3][388] * vector[3] +matrix[4][388] * vector[4] +matrix[5][388] * vector[5] +matrix[6][388] * vector[6] +matrix[7][388] * vector[7] +matrix[8][388] * vector[8] +matrix[9][388] * vector[9] +matrix[10][388] * vector[10] +matrix[11][388] * vector[11] +matrix[12][388] * vector[12] +matrix[13][388] * vector[13] +matrix[14][388] * vector[14] +matrix[15][388] * vector[15] +matrix[16][388] * vector[16] +matrix[17][388] * vector[17] +matrix[18][388] * vector[18] +matrix[19][388] * vector[19] +matrix[20][388] * vector[20] +matrix[21][388] * vector[21] +matrix[22][388] * vector[22] +matrix[23][388] * vector[23] +matrix[24][388] * vector[24] +matrix[25][388] * vector[25] +matrix[26][388] * vector[26] +matrix[27][388] * vector[27] +matrix[28][388] * vector[28] +matrix[29][388] * vector[29] +matrix[30][388] * vector[30] +matrix[31][388] * vector[31] +matrix[32][388] * vector[32] +matrix[33][388] * vector[33] +matrix[34][388] * vector[34] +matrix[35][388] * vector[35] +matrix[36][388] * vector[36] +matrix[37][388] * vector[37] +matrix[38][388] * vector[38] +matrix[39][388] * vector[39] +matrix[40][388] * vector[40] +matrix[41][388] * vector[41] +matrix[42][388] * vector[42] +matrix[43][388] * vector[43] +matrix[44][388] * vector[44] +matrix[45][388] * vector[45] +matrix[46][388] * vector[46] +matrix[47][388] * vector[47] +matrix[48][388] * vector[48] +matrix[49][388] * vector[49] +matrix[50][388] * vector[50] +matrix[51][388] * vector[51] +matrix[52][388] * vector[52] +matrix[53][388] * vector[53] +matrix[54][388] * vector[54] +matrix[55][388] * vector[55] +matrix[56][388] * vector[56] +matrix[57][388] * vector[57] +matrix[58][388] * vector[58] +matrix[59][388] * vector[59] +matrix[60][388] * vector[60] +matrix[61][388] * vector[61] +matrix[62][388] * vector[62] +matrix[63][388] * vector[63] +matrix[64][388] * vector[64] +matrix[65][388] * vector[65] +matrix[66][388] * vector[66] +matrix[67][388] * vector[67] +matrix[68][388] * vector[68] +matrix[69][388] * vector[69] +matrix[70][388] * vector[70] +matrix[71][388] * vector[71] +matrix[72][388] * vector[72] +matrix[73][388] * vector[73] +matrix[74][388] * vector[74] +matrix[75][388] * vector[75] +matrix[76][388] * vector[76] +matrix[77][388] * vector[77] +matrix[78][388] * vector[78] +matrix[79][388] * vector[79] +matrix[80][388] * vector[80] +matrix[81][388] * vector[81] +matrix[82][388] * vector[82] +matrix[83][388] * vector[83] +matrix[84][388] * vector[84] +matrix[85][388] * vector[85] +matrix[86][388] * vector[86] +matrix[87][388] * vector[87] +matrix[88][388] * vector[88] +matrix[89][388] * vector[89] +matrix[90][388] * vector[90] +matrix[91][388] * vector[91] +matrix[92][388] * vector[92] +matrix[93][388] * vector[93] +matrix[94][388] * vector[94] +matrix[95][388] * vector[95] +matrix[96][388] * vector[96] +matrix[97][388] * vector[97] +matrix[98][388] * vector[98] +matrix[99][388] * vector[99] +b[388];
assign result[389] = matrix[0][389] * vector[0] +matrix[1][389] * vector[1] +matrix[2][389] * vector[2] +matrix[3][389] * vector[3] +matrix[4][389] * vector[4] +matrix[5][389] * vector[5] +matrix[6][389] * vector[6] +matrix[7][389] * vector[7] +matrix[8][389] * vector[8] +matrix[9][389] * vector[9] +matrix[10][389] * vector[10] +matrix[11][389] * vector[11] +matrix[12][389] * vector[12] +matrix[13][389] * vector[13] +matrix[14][389] * vector[14] +matrix[15][389] * vector[15] +matrix[16][389] * vector[16] +matrix[17][389] * vector[17] +matrix[18][389] * vector[18] +matrix[19][389] * vector[19] +matrix[20][389] * vector[20] +matrix[21][389] * vector[21] +matrix[22][389] * vector[22] +matrix[23][389] * vector[23] +matrix[24][389] * vector[24] +matrix[25][389] * vector[25] +matrix[26][389] * vector[26] +matrix[27][389] * vector[27] +matrix[28][389] * vector[28] +matrix[29][389] * vector[29] +matrix[30][389] * vector[30] +matrix[31][389] * vector[31] +matrix[32][389] * vector[32] +matrix[33][389] * vector[33] +matrix[34][389] * vector[34] +matrix[35][389] * vector[35] +matrix[36][389] * vector[36] +matrix[37][389] * vector[37] +matrix[38][389] * vector[38] +matrix[39][389] * vector[39] +matrix[40][389] * vector[40] +matrix[41][389] * vector[41] +matrix[42][389] * vector[42] +matrix[43][389] * vector[43] +matrix[44][389] * vector[44] +matrix[45][389] * vector[45] +matrix[46][389] * vector[46] +matrix[47][389] * vector[47] +matrix[48][389] * vector[48] +matrix[49][389] * vector[49] +matrix[50][389] * vector[50] +matrix[51][389] * vector[51] +matrix[52][389] * vector[52] +matrix[53][389] * vector[53] +matrix[54][389] * vector[54] +matrix[55][389] * vector[55] +matrix[56][389] * vector[56] +matrix[57][389] * vector[57] +matrix[58][389] * vector[58] +matrix[59][389] * vector[59] +matrix[60][389] * vector[60] +matrix[61][389] * vector[61] +matrix[62][389] * vector[62] +matrix[63][389] * vector[63] +matrix[64][389] * vector[64] +matrix[65][389] * vector[65] +matrix[66][389] * vector[66] +matrix[67][389] * vector[67] +matrix[68][389] * vector[68] +matrix[69][389] * vector[69] +matrix[70][389] * vector[70] +matrix[71][389] * vector[71] +matrix[72][389] * vector[72] +matrix[73][389] * vector[73] +matrix[74][389] * vector[74] +matrix[75][389] * vector[75] +matrix[76][389] * vector[76] +matrix[77][389] * vector[77] +matrix[78][389] * vector[78] +matrix[79][389] * vector[79] +matrix[80][389] * vector[80] +matrix[81][389] * vector[81] +matrix[82][389] * vector[82] +matrix[83][389] * vector[83] +matrix[84][389] * vector[84] +matrix[85][389] * vector[85] +matrix[86][389] * vector[86] +matrix[87][389] * vector[87] +matrix[88][389] * vector[88] +matrix[89][389] * vector[89] +matrix[90][389] * vector[90] +matrix[91][389] * vector[91] +matrix[92][389] * vector[92] +matrix[93][389] * vector[93] +matrix[94][389] * vector[94] +matrix[95][389] * vector[95] +matrix[96][389] * vector[96] +matrix[97][389] * vector[97] +matrix[98][389] * vector[98] +matrix[99][389] * vector[99] +b[389];
assign result[390] = matrix[0][390] * vector[0] +matrix[1][390] * vector[1] +matrix[2][390] * vector[2] +matrix[3][390] * vector[3] +matrix[4][390] * vector[4] +matrix[5][390] * vector[5] +matrix[6][390] * vector[6] +matrix[7][390] * vector[7] +matrix[8][390] * vector[8] +matrix[9][390] * vector[9] +matrix[10][390] * vector[10] +matrix[11][390] * vector[11] +matrix[12][390] * vector[12] +matrix[13][390] * vector[13] +matrix[14][390] * vector[14] +matrix[15][390] * vector[15] +matrix[16][390] * vector[16] +matrix[17][390] * vector[17] +matrix[18][390] * vector[18] +matrix[19][390] * vector[19] +matrix[20][390] * vector[20] +matrix[21][390] * vector[21] +matrix[22][390] * vector[22] +matrix[23][390] * vector[23] +matrix[24][390] * vector[24] +matrix[25][390] * vector[25] +matrix[26][390] * vector[26] +matrix[27][390] * vector[27] +matrix[28][390] * vector[28] +matrix[29][390] * vector[29] +matrix[30][390] * vector[30] +matrix[31][390] * vector[31] +matrix[32][390] * vector[32] +matrix[33][390] * vector[33] +matrix[34][390] * vector[34] +matrix[35][390] * vector[35] +matrix[36][390] * vector[36] +matrix[37][390] * vector[37] +matrix[38][390] * vector[38] +matrix[39][390] * vector[39] +matrix[40][390] * vector[40] +matrix[41][390] * vector[41] +matrix[42][390] * vector[42] +matrix[43][390] * vector[43] +matrix[44][390] * vector[44] +matrix[45][390] * vector[45] +matrix[46][390] * vector[46] +matrix[47][390] * vector[47] +matrix[48][390] * vector[48] +matrix[49][390] * vector[49] +matrix[50][390] * vector[50] +matrix[51][390] * vector[51] +matrix[52][390] * vector[52] +matrix[53][390] * vector[53] +matrix[54][390] * vector[54] +matrix[55][390] * vector[55] +matrix[56][390] * vector[56] +matrix[57][390] * vector[57] +matrix[58][390] * vector[58] +matrix[59][390] * vector[59] +matrix[60][390] * vector[60] +matrix[61][390] * vector[61] +matrix[62][390] * vector[62] +matrix[63][390] * vector[63] +matrix[64][390] * vector[64] +matrix[65][390] * vector[65] +matrix[66][390] * vector[66] +matrix[67][390] * vector[67] +matrix[68][390] * vector[68] +matrix[69][390] * vector[69] +matrix[70][390] * vector[70] +matrix[71][390] * vector[71] +matrix[72][390] * vector[72] +matrix[73][390] * vector[73] +matrix[74][390] * vector[74] +matrix[75][390] * vector[75] +matrix[76][390] * vector[76] +matrix[77][390] * vector[77] +matrix[78][390] * vector[78] +matrix[79][390] * vector[79] +matrix[80][390] * vector[80] +matrix[81][390] * vector[81] +matrix[82][390] * vector[82] +matrix[83][390] * vector[83] +matrix[84][390] * vector[84] +matrix[85][390] * vector[85] +matrix[86][390] * vector[86] +matrix[87][390] * vector[87] +matrix[88][390] * vector[88] +matrix[89][390] * vector[89] +matrix[90][390] * vector[90] +matrix[91][390] * vector[91] +matrix[92][390] * vector[92] +matrix[93][390] * vector[93] +matrix[94][390] * vector[94] +matrix[95][390] * vector[95] +matrix[96][390] * vector[96] +matrix[97][390] * vector[97] +matrix[98][390] * vector[98] +matrix[99][390] * vector[99] +b[390];
assign result[391] = matrix[0][391] * vector[0] +matrix[1][391] * vector[1] +matrix[2][391] * vector[2] +matrix[3][391] * vector[3] +matrix[4][391] * vector[4] +matrix[5][391] * vector[5] +matrix[6][391] * vector[6] +matrix[7][391] * vector[7] +matrix[8][391] * vector[8] +matrix[9][391] * vector[9] +matrix[10][391] * vector[10] +matrix[11][391] * vector[11] +matrix[12][391] * vector[12] +matrix[13][391] * vector[13] +matrix[14][391] * vector[14] +matrix[15][391] * vector[15] +matrix[16][391] * vector[16] +matrix[17][391] * vector[17] +matrix[18][391] * vector[18] +matrix[19][391] * vector[19] +matrix[20][391] * vector[20] +matrix[21][391] * vector[21] +matrix[22][391] * vector[22] +matrix[23][391] * vector[23] +matrix[24][391] * vector[24] +matrix[25][391] * vector[25] +matrix[26][391] * vector[26] +matrix[27][391] * vector[27] +matrix[28][391] * vector[28] +matrix[29][391] * vector[29] +matrix[30][391] * vector[30] +matrix[31][391] * vector[31] +matrix[32][391] * vector[32] +matrix[33][391] * vector[33] +matrix[34][391] * vector[34] +matrix[35][391] * vector[35] +matrix[36][391] * vector[36] +matrix[37][391] * vector[37] +matrix[38][391] * vector[38] +matrix[39][391] * vector[39] +matrix[40][391] * vector[40] +matrix[41][391] * vector[41] +matrix[42][391] * vector[42] +matrix[43][391] * vector[43] +matrix[44][391] * vector[44] +matrix[45][391] * vector[45] +matrix[46][391] * vector[46] +matrix[47][391] * vector[47] +matrix[48][391] * vector[48] +matrix[49][391] * vector[49] +matrix[50][391] * vector[50] +matrix[51][391] * vector[51] +matrix[52][391] * vector[52] +matrix[53][391] * vector[53] +matrix[54][391] * vector[54] +matrix[55][391] * vector[55] +matrix[56][391] * vector[56] +matrix[57][391] * vector[57] +matrix[58][391] * vector[58] +matrix[59][391] * vector[59] +matrix[60][391] * vector[60] +matrix[61][391] * vector[61] +matrix[62][391] * vector[62] +matrix[63][391] * vector[63] +matrix[64][391] * vector[64] +matrix[65][391] * vector[65] +matrix[66][391] * vector[66] +matrix[67][391] * vector[67] +matrix[68][391] * vector[68] +matrix[69][391] * vector[69] +matrix[70][391] * vector[70] +matrix[71][391] * vector[71] +matrix[72][391] * vector[72] +matrix[73][391] * vector[73] +matrix[74][391] * vector[74] +matrix[75][391] * vector[75] +matrix[76][391] * vector[76] +matrix[77][391] * vector[77] +matrix[78][391] * vector[78] +matrix[79][391] * vector[79] +matrix[80][391] * vector[80] +matrix[81][391] * vector[81] +matrix[82][391] * vector[82] +matrix[83][391] * vector[83] +matrix[84][391] * vector[84] +matrix[85][391] * vector[85] +matrix[86][391] * vector[86] +matrix[87][391] * vector[87] +matrix[88][391] * vector[88] +matrix[89][391] * vector[89] +matrix[90][391] * vector[90] +matrix[91][391] * vector[91] +matrix[92][391] * vector[92] +matrix[93][391] * vector[93] +matrix[94][391] * vector[94] +matrix[95][391] * vector[95] +matrix[96][391] * vector[96] +matrix[97][391] * vector[97] +matrix[98][391] * vector[98] +matrix[99][391] * vector[99] +b[391];
assign result[392] = matrix[0][392] * vector[0] +matrix[1][392] * vector[1] +matrix[2][392] * vector[2] +matrix[3][392] * vector[3] +matrix[4][392] * vector[4] +matrix[5][392] * vector[5] +matrix[6][392] * vector[6] +matrix[7][392] * vector[7] +matrix[8][392] * vector[8] +matrix[9][392] * vector[9] +matrix[10][392] * vector[10] +matrix[11][392] * vector[11] +matrix[12][392] * vector[12] +matrix[13][392] * vector[13] +matrix[14][392] * vector[14] +matrix[15][392] * vector[15] +matrix[16][392] * vector[16] +matrix[17][392] * vector[17] +matrix[18][392] * vector[18] +matrix[19][392] * vector[19] +matrix[20][392] * vector[20] +matrix[21][392] * vector[21] +matrix[22][392] * vector[22] +matrix[23][392] * vector[23] +matrix[24][392] * vector[24] +matrix[25][392] * vector[25] +matrix[26][392] * vector[26] +matrix[27][392] * vector[27] +matrix[28][392] * vector[28] +matrix[29][392] * vector[29] +matrix[30][392] * vector[30] +matrix[31][392] * vector[31] +matrix[32][392] * vector[32] +matrix[33][392] * vector[33] +matrix[34][392] * vector[34] +matrix[35][392] * vector[35] +matrix[36][392] * vector[36] +matrix[37][392] * vector[37] +matrix[38][392] * vector[38] +matrix[39][392] * vector[39] +matrix[40][392] * vector[40] +matrix[41][392] * vector[41] +matrix[42][392] * vector[42] +matrix[43][392] * vector[43] +matrix[44][392] * vector[44] +matrix[45][392] * vector[45] +matrix[46][392] * vector[46] +matrix[47][392] * vector[47] +matrix[48][392] * vector[48] +matrix[49][392] * vector[49] +matrix[50][392] * vector[50] +matrix[51][392] * vector[51] +matrix[52][392] * vector[52] +matrix[53][392] * vector[53] +matrix[54][392] * vector[54] +matrix[55][392] * vector[55] +matrix[56][392] * vector[56] +matrix[57][392] * vector[57] +matrix[58][392] * vector[58] +matrix[59][392] * vector[59] +matrix[60][392] * vector[60] +matrix[61][392] * vector[61] +matrix[62][392] * vector[62] +matrix[63][392] * vector[63] +matrix[64][392] * vector[64] +matrix[65][392] * vector[65] +matrix[66][392] * vector[66] +matrix[67][392] * vector[67] +matrix[68][392] * vector[68] +matrix[69][392] * vector[69] +matrix[70][392] * vector[70] +matrix[71][392] * vector[71] +matrix[72][392] * vector[72] +matrix[73][392] * vector[73] +matrix[74][392] * vector[74] +matrix[75][392] * vector[75] +matrix[76][392] * vector[76] +matrix[77][392] * vector[77] +matrix[78][392] * vector[78] +matrix[79][392] * vector[79] +matrix[80][392] * vector[80] +matrix[81][392] * vector[81] +matrix[82][392] * vector[82] +matrix[83][392] * vector[83] +matrix[84][392] * vector[84] +matrix[85][392] * vector[85] +matrix[86][392] * vector[86] +matrix[87][392] * vector[87] +matrix[88][392] * vector[88] +matrix[89][392] * vector[89] +matrix[90][392] * vector[90] +matrix[91][392] * vector[91] +matrix[92][392] * vector[92] +matrix[93][392] * vector[93] +matrix[94][392] * vector[94] +matrix[95][392] * vector[95] +matrix[96][392] * vector[96] +matrix[97][392] * vector[97] +matrix[98][392] * vector[98] +matrix[99][392] * vector[99] +b[392];
assign result[393] = matrix[0][393] * vector[0] +matrix[1][393] * vector[1] +matrix[2][393] * vector[2] +matrix[3][393] * vector[3] +matrix[4][393] * vector[4] +matrix[5][393] * vector[5] +matrix[6][393] * vector[6] +matrix[7][393] * vector[7] +matrix[8][393] * vector[8] +matrix[9][393] * vector[9] +matrix[10][393] * vector[10] +matrix[11][393] * vector[11] +matrix[12][393] * vector[12] +matrix[13][393] * vector[13] +matrix[14][393] * vector[14] +matrix[15][393] * vector[15] +matrix[16][393] * vector[16] +matrix[17][393] * vector[17] +matrix[18][393] * vector[18] +matrix[19][393] * vector[19] +matrix[20][393] * vector[20] +matrix[21][393] * vector[21] +matrix[22][393] * vector[22] +matrix[23][393] * vector[23] +matrix[24][393] * vector[24] +matrix[25][393] * vector[25] +matrix[26][393] * vector[26] +matrix[27][393] * vector[27] +matrix[28][393] * vector[28] +matrix[29][393] * vector[29] +matrix[30][393] * vector[30] +matrix[31][393] * vector[31] +matrix[32][393] * vector[32] +matrix[33][393] * vector[33] +matrix[34][393] * vector[34] +matrix[35][393] * vector[35] +matrix[36][393] * vector[36] +matrix[37][393] * vector[37] +matrix[38][393] * vector[38] +matrix[39][393] * vector[39] +matrix[40][393] * vector[40] +matrix[41][393] * vector[41] +matrix[42][393] * vector[42] +matrix[43][393] * vector[43] +matrix[44][393] * vector[44] +matrix[45][393] * vector[45] +matrix[46][393] * vector[46] +matrix[47][393] * vector[47] +matrix[48][393] * vector[48] +matrix[49][393] * vector[49] +matrix[50][393] * vector[50] +matrix[51][393] * vector[51] +matrix[52][393] * vector[52] +matrix[53][393] * vector[53] +matrix[54][393] * vector[54] +matrix[55][393] * vector[55] +matrix[56][393] * vector[56] +matrix[57][393] * vector[57] +matrix[58][393] * vector[58] +matrix[59][393] * vector[59] +matrix[60][393] * vector[60] +matrix[61][393] * vector[61] +matrix[62][393] * vector[62] +matrix[63][393] * vector[63] +matrix[64][393] * vector[64] +matrix[65][393] * vector[65] +matrix[66][393] * vector[66] +matrix[67][393] * vector[67] +matrix[68][393] * vector[68] +matrix[69][393] * vector[69] +matrix[70][393] * vector[70] +matrix[71][393] * vector[71] +matrix[72][393] * vector[72] +matrix[73][393] * vector[73] +matrix[74][393] * vector[74] +matrix[75][393] * vector[75] +matrix[76][393] * vector[76] +matrix[77][393] * vector[77] +matrix[78][393] * vector[78] +matrix[79][393] * vector[79] +matrix[80][393] * vector[80] +matrix[81][393] * vector[81] +matrix[82][393] * vector[82] +matrix[83][393] * vector[83] +matrix[84][393] * vector[84] +matrix[85][393] * vector[85] +matrix[86][393] * vector[86] +matrix[87][393] * vector[87] +matrix[88][393] * vector[88] +matrix[89][393] * vector[89] +matrix[90][393] * vector[90] +matrix[91][393] * vector[91] +matrix[92][393] * vector[92] +matrix[93][393] * vector[93] +matrix[94][393] * vector[94] +matrix[95][393] * vector[95] +matrix[96][393] * vector[96] +matrix[97][393] * vector[97] +matrix[98][393] * vector[98] +matrix[99][393] * vector[99] +b[393];
assign result[394] = matrix[0][394] * vector[0] +matrix[1][394] * vector[1] +matrix[2][394] * vector[2] +matrix[3][394] * vector[3] +matrix[4][394] * vector[4] +matrix[5][394] * vector[5] +matrix[6][394] * vector[6] +matrix[7][394] * vector[7] +matrix[8][394] * vector[8] +matrix[9][394] * vector[9] +matrix[10][394] * vector[10] +matrix[11][394] * vector[11] +matrix[12][394] * vector[12] +matrix[13][394] * vector[13] +matrix[14][394] * vector[14] +matrix[15][394] * vector[15] +matrix[16][394] * vector[16] +matrix[17][394] * vector[17] +matrix[18][394] * vector[18] +matrix[19][394] * vector[19] +matrix[20][394] * vector[20] +matrix[21][394] * vector[21] +matrix[22][394] * vector[22] +matrix[23][394] * vector[23] +matrix[24][394] * vector[24] +matrix[25][394] * vector[25] +matrix[26][394] * vector[26] +matrix[27][394] * vector[27] +matrix[28][394] * vector[28] +matrix[29][394] * vector[29] +matrix[30][394] * vector[30] +matrix[31][394] * vector[31] +matrix[32][394] * vector[32] +matrix[33][394] * vector[33] +matrix[34][394] * vector[34] +matrix[35][394] * vector[35] +matrix[36][394] * vector[36] +matrix[37][394] * vector[37] +matrix[38][394] * vector[38] +matrix[39][394] * vector[39] +matrix[40][394] * vector[40] +matrix[41][394] * vector[41] +matrix[42][394] * vector[42] +matrix[43][394] * vector[43] +matrix[44][394] * vector[44] +matrix[45][394] * vector[45] +matrix[46][394] * vector[46] +matrix[47][394] * vector[47] +matrix[48][394] * vector[48] +matrix[49][394] * vector[49] +matrix[50][394] * vector[50] +matrix[51][394] * vector[51] +matrix[52][394] * vector[52] +matrix[53][394] * vector[53] +matrix[54][394] * vector[54] +matrix[55][394] * vector[55] +matrix[56][394] * vector[56] +matrix[57][394] * vector[57] +matrix[58][394] * vector[58] +matrix[59][394] * vector[59] +matrix[60][394] * vector[60] +matrix[61][394] * vector[61] +matrix[62][394] * vector[62] +matrix[63][394] * vector[63] +matrix[64][394] * vector[64] +matrix[65][394] * vector[65] +matrix[66][394] * vector[66] +matrix[67][394] * vector[67] +matrix[68][394] * vector[68] +matrix[69][394] * vector[69] +matrix[70][394] * vector[70] +matrix[71][394] * vector[71] +matrix[72][394] * vector[72] +matrix[73][394] * vector[73] +matrix[74][394] * vector[74] +matrix[75][394] * vector[75] +matrix[76][394] * vector[76] +matrix[77][394] * vector[77] +matrix[78][394] * vector[78] +matrix[79][394] * vector[79] +matrix[80][394] * vector[80] +matrix[81][394] * vector[81] +matrix[82][394] * vector[82] +matrix[83][394] * vector[83] +matrix[84][394] * vector[84] +matrix[85][394] * vector[85] +matrix[86][394] * vector[86] +matrix[87][394] * vector[87] +matrix[88][394] * vector[88] +matrix[89][394] * vector[89] +matrix[90][394] * vector[90] +matrix[91][394] * vector[91] +matrix[92][394] * vector[92] +matrix[93][394] * vector[93] +matrix[94][394] * vector[94] +matrix[95][394] * vector[95] +matrix[96][394] * vector[96] +matrix[97][394] * vector[97] +matrix[98][394] * vector[98] +matrix[99][394] * vector[99] +b[394];
assign result[395] = matrix[0][395] * vector[0] +matrix[1][395] * vector[1] +matrix[2][395] * vector[2] +matrix[3][395] * vector[3] +matrix[4][395] * vector[4] +matrix[5][395] * vector[5] +matrix[6][395] * vector[6] +matrix[7][395] * vector[7] +matrix[8][395] * vector[8] +matrix[9][395] * vector[9] +matrix[10][395] * vector[10] +matrix[11][395] * vector[11] +matrix[12][395] * vector[12] +matrix[13][395] * vector[13] +matrix[14][395] * vector[14] +matrix[15][395] * vector[15] +matrix[16][395] * vector[16] +matrix[17][395] * vector[17] +matrix[18][395] * vector[18] +matrix[19][395] * vector[19] +matrix[20][395] * vector[20] +matrix[21][395] * vector[21] +matrix[22][395] * vector[22] +matrix[23][395] * vector[23] +matrix[24][395] * vector[24] +matrix[25][395] * vector[25] +matrix[26][395] * vector[26] +matrix[27][395] * vector[27] +matrix[28][395] * vector[28] +matrix[29][395] * vector[29] +matrix[30][395] * vector[30] +matrix[31][395] * vector[31] +matrix[32][395] * vector[32] +matrix[33][395] * vector[33] +matrix[34][395] * vector[34] +matrix[35][395] * vector[35] +matrix[36][395] * vector[36] +matrix[37][395] * vector[37] +matrix[38][395] * vector[38] +matrix[39][395] * vector[39] +matrix[40][395] * vector[40] +matrix[41][395] * vector[41] +matrix[42][395] * vector[42] +matrix[43][395] * vector[43] +matrix[44][395] * vector[44] +matrix[45][395] * vector[45] +matrix[46][395] * vector[46] +matrix[47][395] * vector[47] +matrix[48][395] * vector[48] +matrix[49][395] * vector[49] +matrix[50][395] * vector[50] +matrix[51][395] * vector[51] +matrix[52][395] * vector[52] +matrix[53][395] * vector[53] +matrix[54][395] * vector[54] +matrix[55][395] * vector[55] +matrix[56][395] * vector[56] +matrix[57][395] * vector[57] +matrix[58][395] * vector[58] +matrix[59][395] * vector[59] +matrix[60][395] * vector[60] +matrix[61][395] * vector[61] +matrix[62][395] * vector[62] +matrix[63][395] * vector[63] +matrix[64][395] * vector[64] +matrix[65][395] * vector[65] +matrix[66][395] * vector[66] +matrix[67][395] * vector[67] +matrix[68][395] * vector[68] +matrix[69][395] * vector[69] +matrix[70][395] * vector[70] +matrix[71][395] * vector[71] +matrix[72][395] * vector[72] +matrix[73][395] * vector[73] +matrix[74][395] * vector[74] +matrix[75][395] * vector[75] +matrix[76][395] * vector[76] +matrix[77][395] * vector[77] +matrix[78][395] * vector[78] +matrix[79][395] * vector[79] +matrix[80][395] * vector[80] +matrix[81][395] * vector[81] +matrix[82][395] * vector[82] +matrix[83][395] * vector[83] +matrix[84][395] * vector[84] +matrix[85][395] * vector[85] +matrix[86][395] * vector[86] +matrix[87][395] * vector[87] +matrix[88][395] * vector[88] +matrix[89][395] * vector[89] +matrix[90][395] * vector[90] +matrix[91][395] * vector[91] +matrix[92][395] * vector[92] +matrix[93][395] * vector[93] +matrix[94][395] * vector[94] +matrix[95][395] * vector[95] +matrix[96][395] * vector[96] +matrix[97][395] * vector[97] +matrix[98][395] * vector[98] +matrix[99][395] * vector[99] +b[395];
assign result[396] = matrix[0][396] * vector[0] +matrix[1][396] * vector[1] +matrix[2][396] * vector[2] +matrix[3][396] * vector[3] +matrix[4][396] * vector[4] +matrix[5][396] * vector[5] +matrix[6][396] * vector[6] +matrix[7][396] * vector[7] +matrix[8][396] * vector[8] +matrix[9][396] * vector[9] +matrix[10][396] * vector[10] +matrix[11][396] * vector[11] +matrix[12][396] * vector[12] +matrix[13][396] * vector[13] +matrix[14][396] * vector[14] +matrix[15][396] * vector[15] +matrix[16][396] * vector[16] +matrix[17][396] * vector[17] +matrix[18][396] * vector[18] +matrix[19][396] * vector[19] +matrix[20][396] * vector[20] +matrix[21][396] * vector[21] +matrix[22][396] * vector[22] +matrix[23][396] * vector[23] +matrix[24][396] * vector[24] +matrix[25][396] * vector[25] +matrix[26][396] * vector[26] +matrix[27][396] * vector[27] +matrix[28][396] * vector[28] +matrix[29][396] * vector[29] +matrix[30][396] * vector[30] +matrix[31][396] * vector[31] +matrix[32][396] * vector[32] +matrix[33][396] * vector[33] +matrix[34][396] * vector[34] +matrix[35][396] * vector[35] +matrix[36][396] * vector[36] +matrix[37][396] * vector[37] +matrix[38][396] * vector[38] +matrix[39][396] * vector[39] +matrix[40][396] * vector[40] +matrix[41][396] * vector[41] +matrix[42][396] * vector[42] +matrix[43][396] * vector[43] +matrix[44][396] * vector[44] +matrix[45][396] * vector[45] +matrix[46][396] * vector[46] +matrix[47][396] * vector[47] +matrix[48][396] * vector[48] +matrix[49][396] * vector[49] +matrix[50][396] * vector[50] +matrix[51][396] * vector[51] +matrix[52][396] * vector[52] +matrix[53][396] * vector[53] +matrix[54][396] * vector[54] +matrix[55][396] * vector[55] +matrix[56][396] * vector[56] +matrix[57][396] * vector[57] +matrix[58][396] * vector[58] +matrix[59][396] * vector[59] +matrix[60][396] * vector[60] +matrix[61][396] * vector[61] +matrix[62][396] * vector[62] +matrix[63][396] * vector[63] +matrix[64][396] * vector[64] +matrix[65][396] * vector[65] +matrix[66][396] * vector[66] +matrix[67][396] * vector[67] +matrix[68][396] * vector[68] +matrix[69][396] * vector[69] +matrix[70][396] * vector[70] +matrix[71][396] * vector[71] +matrix[72][396] * vector[72] +matrix[73][396] * vector[73] +matrix[74][396] * vector[74] +matrix[75][396] * vector[75] +matrix[76][396] * vector[76] +matrix[77][396] * vector[77] +matrix[78][396] * vector[78] +matrix[79][396] * vector[79] +matrix[80][396] * vector[80] +matrix[81][396] * vector[81] +matrix[82][396] * vector[82] +matrix[83][396] * vector[83] +matrix[84][396] * vector[84] +matrix[85][396] * vector[85] +matrix[86][396] * vector[86] +matrix[87][396] * vector[87] +matrix[88][396] * vector[88] +matrix[89][396] * vector[89] +matrix[90][396] * vector[90] +matrix[91][396] * vector[91] +matrix[92][396] * vector[92] +matrix[93][396] * vector[93] +matrix[94][396] * vector[94] +matrix[95][396] * vector[95] +matrix[96][396] * vector[96] +matrix[97][396] * vector[97] +matrix[98][396] * vector[98] +matrix[99][396] * vector[99] +b[396];
assign result[397] = matrix[0][397] * vector[0] +matrix[1][397] * vector[1] +matrix[2][397] * vector[2] +matrix[3][397] * vector[3] +matrix[4][397] * vector[4] +matrix[5][397] * vector[5] +matrix[6][397] * vector[6] +matrix[7][397] * vector[7] +matrix[8][397] * vector[8] +matrix[9][397] * vector[9] +matrix[10][397] * vector[10] +matrix[11][397] * vector[11] +matrix[12][397] * vector[12] +matrix[13][397] * vector[13] +matrix[14][397] * vector[14] +matrix[15][397] * vector[15] +matrix[16][397] * vector[16] +matrix[17][397] * vector[17] +matrix[18][397] * vector[18] +matrix[19][397] * vector[19] +matrix[20][397] * vector[20] +matrix[21][397] * vector[21] +matrix[22][397] * vector[22] +matrix[23][397] * vector[23] +matrix[24][397] * vector[24] +matrix[25][397] * vector[25] +matrix[26][397] * vector[26] +matrix[27][397] * vector[27] +matrix[28][397] * vector[28] +matrix[29][397] * vector[29] +matrix[30][397] * vector[30] +matrix[31][397] * vector[31] +matrix[32][397] * vector[32] +matrix[33][397] * vector[33] +matrix[34][397] * vector[34] +matrix[35][397] * vector[35] +matrix[36][397] * vector[36] +matrix[37][397] * vector[37] +matrix[38][397] * vector[38] +matrix[39][397] * vector[39] +matrix[40][397] * vector[40] +matrix[41][397] * vector[41] +matrix[42][397] * vector[42] +matrix[43][397] * vector[43] +matrix[44][397] * vector[44] +matrix[45][397] * vector[45] +matrix[46][397] * vector[46] +matrix[47][397] * vector[47] +matrix[48][397] * vector[48] +matrix[49][397] * vector[49] +matrix[50][397] * vector[50] +matrix[51][397] * vector[51] +matrix[52][397] * vector[52] +matrix[53][397] * vector[53] +matrix[54][397] * vector[54] +matrix[55][397] * vector[55] +matrix[56][397] * vector[56] +matrix[57][397] * vector[57] +matrix[58][397] * vector[58] +matrix[59][397] * vector[59] +matrix[60][397] * vector[60] +matrix[61][397] * vector[61] +matrix[62][397] * vector[62] +matrix[63][397] * vector[63] +matrix[64][397] * vector[64] +matrix[65][397] * vector[65] +matrix[66][397] * vector[66] +matrix[67][397] * vector[67] +matrix[68][397] * vector[68] +matrix[69][397] * vector[69] +matrix[70][397] * vector[70] +matrix[71][397] * vector[71] +matrix[72][397] * vector[72] +matrix[73][397] * vector[73] +matrix[74][397] * vector[74] +matrix[75][397] * vector[75] +matrix[76][397] * vector[76] +matrix[77][397] * vector[77] +matrix[78][397] * vector[78] +matrix[79][397] * vector[79] +matrix[80][397] * vector[80] +matrix[81][397] * vector[81] +matrix[82][397] * vector[82] +matrix[83][397] * vector[83] +matrix[84][397] * vector[84] +matrix[85][397] * vector[85] +matrix[86][397] * vector[86] +matrix[87][397] * vector[87] +matrix[88][397] * vector[88] +matrix[89][397] * vector[89] +matrix[90][397] * vector[90] +matrix[91][397] * vector[91] +matrix[92][397] * vector[92] +matrix[93][397] * vector[93] +matrix[94][397] * vector[94] +matrix[95][397] * vector[95] +matrix[96][397] * vector[96] +matrix[97][397] * vector[97] +matrix[98][397] * vector[98] +matrix[99][397] * vector[99] +b[397];
assign result[398] = matrix[0][398] * vector[0] +matrix[1][398] * vector[1] +matrix[2][398] * vector[2] +matrix[3][398] * vector[3] +matrix[4][398] * vector[4] +matrix[5][398] * vector[5] +matrix[6][398] * vector[6] +matrix[7][398] * vector[7] +matrix[8][398] * vector[8] +matrix[9][398] * vector[9] +matrix[10][398] * vector[10] +matrix[11][398] * vector[11] +matrix[12][398] * vector[12] +matrix[13][398] * vector[13] +matrix[14][398] * vector[14] +matrix[15][398] * vector[15] +matrix[16][398] * vector[16] +matrix[17][398] * vector[17] +matrix[18][398] * vector[18] +matrix[19][398] * vector[19] +matrix[20][398] * vector[20] +matrix[21][398] * vector[21] +matrix[22][398] * vector[22] +matrix[23][398] * vector[23] +matrix[24][398] * vector[24] +matrix[25][398] * vector[25] +matrix[26][398] * vector[26] +matrix[27][398] * vector[27] +matrix[28][398] * vector[28] +matrix[29][398] * vector[29] +matrix[30][398] * vector[30] +matrix[31][398] * vector[31] +matrix[32][398] * vector[32] +matrix[33][398] * vector[33] +matrix[34][398] * vector[34] +matrix[35][398] * vector[35] +matrix[36][398] * vector[36] +matrix[37][398] * vector[37] +matrix[38][398] * vector[38] +matrix[39][398] * vector[39] +matrix[40][398] * vector[40] +matrix[41][398] * vector[41] +matrix[42][398] * vector[42] +matrix[43][398] * vector[43] +matrix[44][398] * vector[44] +matrix[45][398] * vector[45] +matrix[46][398] * vector[46] +matrix[47][398] * vector[47] +matrix[48][398] * vector[48] +matrix[49][398] * vector[49] +matrix[50][398] * vector[50] +matrix[51][398] * vector[51] +matrix[52][398] * vector[52] +matrix[53][398] * vector[53] +matrix[54][398] * vector[54] +matrix[55][398] * vector[55] +matrix[56][398] * vector[56] +matrix[57][398] * vector[57] +matrix[58][398] * vector[58] +matrix[59][398] * vector[59] +matrix[60][398] * vector[60] +matrix[61][398] * vector[61] +matrix[62][398] * vector[62] +matrix[63][398] * vector[63] +matrix[64][398] * vector[64] +matrix[65][398] * vector[65] +matrix[66][398] * vector[66] +matrix[67][398] * vector[67] +matrix[68][398] * vector[68] +matrix[69][398] * vector[69] +matrix[70][398] * vector[70] +matrix[71][398] * vector[71] +matrix[72][398] * vector[72] +matrix[73][398] * vector[73] +matrix[74][398] * vector[74] +matrix[75][398] * vector[75] +matrix[76][398] * vector[76] +matrix[77][398] * vector[77] +matrix[78][398] * vector[78] +matrix[79][398] * vector[79] +matrix[80][398] * vector[80] +matrix[81][398] * vector[81] +matrix[82][398] * vector[82] +matrix[83][398] * vector[83] +matrix[84][398] * vector[84] +matrix[85][398] * vector[85] +matrix[86][398] * vector[86] +matrix[87][398] * vector[87] +matrix[88][398] * vector[88] +matrix[89][398] * vector[89] +matrix[90][398] * vector[90] +matrix[91][398] * vector[91] +matrix[92][398] * vector[92] +matrix[93][398] * vector[93] +matrix[94][398] * vector[94] +matrix[95][398] * vector[95] +matrix[96][398] * vector[96] +matrix[97][398] * vector[97] +matrix[98][398] * vector[98] +matrix[99][398] * vector[99] +b[398];
assign result[399] = matrix[0][399] * vector[0] +matrix[1][399] * vector[1] +matrix[2][399] * vector[2] +matrix[3][399] * vector[3] +matrix[4][399] * vector[4] +matrix[5][399] * vector[5] +matrix[6][399] * vector[6] +matrix[7][399] * vector[7] +matrix[8][399] * vector[8] +matrix[9][399] * vector[9] +matrix[10][399] * vector[10] +matrix[11][399] * vector[11] +matrix[12][399] * vector[12] +matrix[13][399] * vector[13] +matrix[14][399] * vector[14] +matrix[15][399] * vector[15] +matrix[16][399] * vector[16] +matrix[17][399] * vector[17] +matrix[18][399] * vector[18] +matrix[19][399] * vector[19] +matrix[20][399] * vector[20] +matrix[21][399] * vector[21] +matrix[22][399] * vector[22] +matrix[23][399] * vector[23] +matrix[24][399] * vector[24] +matrix[25][399] * vector[25] +matrix[26][399] * vector[26] +matrix[27][399] * vector[27] +matrix[28][399] * vector[28] +matrix[29][399] * vector[29] +matrix[30][399] * vector[30] +matrix[31][399] * vector[31] +matrix[32][399] * vector[32] +matrix[33][399] * vector[33] +matrix[34][399] * vector[34] +matrix[35][399] * vector[35] +matrix[36][399] * vector[36] +matrix[37][399] * vector[37] +matrix[38][399] * vector[38] +matrix[39][399] * vector[39] +matrix[40][399] * vector[40] +matrix[41][399] * vector[41] +matrix[42][399] * vector[42] +matrix[43][399] * vector[43] +matrix[44][399] * vector[44] +matrix[45][399] * vector[45] +matrix[46][399] * vector[46] +matrix[47][399] * vector[47] +matrix[48][399] * vector[48] +matrix[49][399] * vector[49] +matrix[50][399] * vector[50] +matrix[51][399] * vector[51] +matrix[52][399] * vector[52] +matrix[53][399] * vector[53] +matrix[54][399] * vector[54] +matrix[55][399] * vector[55] +matrix[56][399] * vector[56] +matrix[57][399] * vector[57] +matrix[58][399] * vector[58] +matrix[59][399] * vector[59] +matrix[60][399] * vector[60] +matrix[61][399] * vector[61] +matrix[62][399] * vector[62] +matrix[63][399] * vector[63] +matrix[64][399] * vector[64] +matrix[65][399] * vector[65] +matrix[66][399] * vector[66] +matrix[67][399] * vector[67] +matrix[68][399] * vector[68] +matrix[69][399] * vector[69] +matrix[70][399] * vector[70] +matrix[71][399] * vector[71] +matrix[72][399] * vector[72] +matrix[73][399] * vector[73] +matrix[74][399] * vector[74] +matrix[75][399] * vector[75] +matrix[76][399] * vector[76] +matrix[77][399] * vector[77] +matrix[78][399] * vector[78] +matrix[79][399] * vector[79] +matrix[80][399] * vector[80] +matrix[81][399] * vector[81] +matrix[82][399] * vector[82] +matrix[83][399] * vector[83] +matrix[84][399] * vector[84] +matrix[85][399] * vector[85] +matrix[86][399] * vector[86] +matrix[87][399] * vector[87] +matrix[88][399] * vector[88] +matrix[89][399] * vector[89] +matrix[90][399] * vector[90] +matrix[91][399] * vector[91] +matrix[92][399] * vector[92] +matrix[93][399] * vector[93] +matrix[94][399] * vector[94] +matrix[95][399] * vector[95] +matrix[96][399] * vector[96] +matrix[97][399] * vector[97] +matrix[98][399] * vector[98] +matrix[99][399] * vector[99] +b[399];

endmodule
