`include "tanh.sv"
module tanh_tb; reg signed [31:0] x; wire signed [31:0] y; tanh dut (.x(x),
                                                                     .y(y));
    
    // Clock
    reg clk;
    
    // Initialize clock
    initial begin
        clk            = 0;
        forever #5 clk = ~clk;
    end
    
    // Stimulus
    initial begin
        
#10;x=-240000000;
#10;x=-239990000;
#10;x=-239980000;
#10;x=-239970000;
#10;x=-239960000;
#10;x=-239950000;
#10;x=-239940000;
#10;x=-239930000;
#10;x=-239920000;
#10;x=-239910000;
#10;x=-239900000;
#10;x=-239890000;
#10;x=-239880000;
#10;x=-239870000;
#10;x=-239860000;
#10;x=-239850000;
#10;x=-239840000;
#10;x=-239830000;
#10;x=-239820000;
#10;x=-239810000;
#10;x=-239800000;
#10;x=-239790000;
#10;x=-239780000;
#10;x=-239770000;
#10;x=-239760000;
#10;x=-239750000;
#10;x=-239740000;
#10;x=-239730000;
#10;x=-239720000;
#10;x=-239710000;
#10;x=-239700000;
#10;x=-239690000;
#10;x=-239680000;
#10;x=-239670000;
#10;x=-239660000;
#10;x=-239650000;
#10;x=-239640000;
#10;x=-239630000;
#10;x=-239620000;
#10;x=-239610000;
#10;x=-239600000;
#10;x=-239590000;
#10;x=-239580000;
#10;x=-239570000;
#10;x=-239560000;
#10;x=-239550000;
#10;x=-239540000;
#10;x=-239530000;
#10;x=-239520000;
#10;x=-239510000;
#10;x=-239500000;
#10;x=-239490000;
#10;x=-239480000;
#10;x=-239470000;
#10;x=-239460000;
#10;x=-239450000;
#10;x=-239440000;
#10;x=-239430000;
#10;x=-239420000;
#10;x=-239410000;
#10;x=-239400000;
#10;x=-239390000;
#10;x=-239380000;
#10;x=-239370000;
#10;x=-239360000;
#10;x=-239350000;
#10;x=-239340000;
#10;x=-239330000;
#10;x=-239320000;
#10;x=-239310000;
#10;x=-239300000;
#10;x=-239290000;
#10;x=-239280000;
#10;x=-239270000;
#10;x=-239260000;
#10;x=-239250000;
#10;x=-239240000;
#10;x=-239230000;
#10;x=-239220000;
#10;x=-239210000;
#10;x=-239200000;
#10;x=-239190000;
#10;x=-239180000;
#10;x=-239170000;
#10;x=-239160000;
#10;x=-239150000;
#10;x=-239140000;
#10;x=-239130000;
#10;x=-239120000;
#10;x=-239110000;
#10;x=-239100000;
#10;x=-239090000;
#10;x=-239080000;
#10;x=-239070000;
#10;x=-239060000;
#10;x=-239050000;
#10;x=-239040000;
#10;x=-239030000;
#10;x=-239020000;
#10;x=-239010000;
#10;x=-239000000;
#10;x=-238990000;
#10;x=-238980000;
#10;x=-238970000;
#10;x=-238960000;
#10;x=-238950000;
#10;x=-238940000;
#10;x=-238930000;
#10;x=-238920000;
#10;x=-238910000;
#10;x=-238900000;
#10;x=-238890000;
#10;x=-238880000;
#10;x=-238870000;
#10;x=-238860000;
#10;x=-238850000;
#10;x=-238840000;
#10;x=-238830000;
#10;x=-238820000;
#10;x=-238810000;
#10;x=-238800000;
#10;x=-238790000;
#10;x=-238780000;
#10;x=-238770000;
#10;x=-238760000;
#10;x=-238750000;
#10;x=-238740000;
#10;x=-238730000;
#10;x=-238720000;
#10;x=-238710000;
#10;x=-238700000;
#10;x=-238690000;
#10;x=-238680000;
#10;x=-238670000;
#10;x=-238660000;
#10;x=-238650000;
#10;x=-238640000;
#10;x=-238630000;
#10;x=-238620000;
#10;x=-238610000;
#10;x=-238600000;
#10;x=-238590000;
#10;x=-238580000;
#10;x=-238570000;
#10;x=-238560000;
#10;x=-238550000;
#10;x=-238540000;
#10;x=-238530000;
#10;x=-238520000;
#10;x=-238510000;
#10;x=-238500000;
#10;x=-238490000;
#10;x=-238480000;
#10;x=-238470000;
#10;x=-238460000;
#10;x=-238450000;
#10;x=-238440000;
#10;x=-238430000;
#10;x=-238420000;
#10;x=-238410000;
#10;x=-238400000;
#10;x=-238390000;
#10;x=-238380000;
#10;x=-238370000;
#10;x=-238360000;
#10;x=-238350000;
#10;x=-238340000;
#10;x=-238330000;
#10;x=-238320000;
#10;x=-238310000;
#10;x=-238300000;
#10;x=-238290000;
#10;x=-238280000;
#10;x=-238270000;
#10;x=-238260000;
#10;x=-238250000;
#10;x=-238240000;
#10;x=-238230000;
#10;x=-238220000;
#10;x=-238210000;
#10;x=-238200000;
#10;x=-238190000;
#10;x=-238180000;
#10;x=-238170000;
#10;x=-238160000;
#10;x=-238150000;
#10;x=-238140000;
#10;x=-238130000;
#10;x=-238120000;
#10;x=-238110000;
#10;x=-238100000;
#10;x=-238090000;
#10;x=-238080000;
#10;x=-238070000;
#10;x=-238060000;
#10;x=-238050000;
#10;x=-238040000;
#10;x=-238030000;
#10;x=-238020000;
#10;x=-238010000;
#10;x=-238000000;
#10;x=-237990000;
#10;x=-237980000;
#10;x=-237970000;
#10;x=-237960000;
#10;x=-237950000;
#10;x=-237940000;
#10;x=-237930000;
#10;x=-237920000;
#10;x=-237910000;
#10;x=-237900000;
#10;x=-237890000;
#10;x=-237880000;
#10;x=-237870000;
#10;x=-237860000;
#10;x=-237850000;
#10;x=-237840000;
#10;x=-237830000;
#10;x=-237820000;
#10;x=-237810000;
#10;x=-237800000;
#10;x=-237790000;
#10;x=-237780000;
#10;x=-237770000;
#10;x=-237760000;
#10;x=-237750000;
#10;x=-237740000;
#10;x=-237730000;
#10;x=-237720000;
#10;x=-237710000;
#10;x=-237700000;
#10;x=-237690000;
#10;x=-237680000;
#10;x=-237670000;
#10;x=-237660000;
#10;x=-237650000;
#10;x=-237640000;
#10;x=-237630000;
#10;x=-237620000;
#10;x=-237610000;
#10;x=-237600000;
#10;x=-237590000;
#10;x=-237580000;
#10;x=-237570000;
#10;x=-237560000;
#10;x=-237550000;
#10;x=-237540000;
#10;x=-237530000;
#10;x=-237520000;
#10;x=-237510000;
#10;x=-237500000;
#10;x=-237490000;
#10;x=-237480000;
#10;x=-237470000;
#10;x=-237460000;
#10;x=-237450000;
#10;x=-237440000;
#10;x=-237430000;
#10;x=-237420000;
#10;x=-237410000;
#10;x=-237400000;
#10;x=-237390000;
#10;x=-237380000;
#10;x=-237370000;
#10;x=-237360000;
#10;x=-237350000;
#10;x=-237340000;
#10;x=-237330000;
#10;x=-237320000;
#10;x=-237310000;
#10;x=-237300000;
#10;x=-237290000;
#10;x=-237280000;
#10;x=-237270000;
#10;x=-237260000;
#10;x=-237250000;
#10;x=-237240000;
#10;x=-237230000;
#10;x=-237220000;
#10;x=-237210000;
#10;x=-237200000;
#10;x=-237190000;
#10;x=-237180000;
#10;x=-237170000;
#10;x=-237160000;
#10;x=-237150000;
#10;x=-237140000;
#10;x=-237130000;
#10;x=-237120000;
#10;x=-237110000;
#10;x=-237100000;
#10;x=-237090000;
#10;x=-237080000;
#10;x=-237070000;
#10;x=-237060000;
#10;x=-237050000;
#10;x=-237040000;
#10;x=-237030000;
#10;x=-237020000;
#10;x=-237010000;
#10;x=-237000000;
#10;x=-236990000;
#10;x=-236980000;
#10;x=-236970000;
#10;x=-236960000;
#10;x=-236950000;
#10;x=-236940000;
#10;x=-236930000;
#10;x=-236920000;
#10;x=-236910000;
#10;x=-236900000;
#10;x=-236890000;
#10;x=-236880000;
#10;x=-236870000;
#10;x=-236860000;
#10;x=-236850000;
#10;x=-236840000;
#10;x=-236830000;
#10;x=-236820000;
#10;x=-236810000;
#10;x=-236800000;
#10;x=-236790000;
#10;x=-236780000;
#10;x=-236770000;
#10;x=-236760000;
#10;x=-236750000;
#10;x=-236740000;
#10;x=-236730000;
#10;x=-236720000;
#10;x=-236710000;
#10;x=-236700000;
#10;x=-236690000;
#10;x=-236680000;
#10;x=-236670000;
#10;x=-236660000;
#10;x=-236650000;
#10;x=-236640000;
#10;x=-236630000;
#10;x=-236620000;
#10;x=-236610000;
#10;x=-236600000;
#10;x=-236590000;
#10;x=-236580000;
#10;x=-236570000;
#10;x=-236560000;
#10;x=-236550000;
#10;x=-236540000;
#10;x=-236530000;
#10;x=-236520000;
#10;x=-236510000;
#10;x=-236500000;
#10;x=-236490000;
#10;x=-236480000;
#10;x=-236470000;
#10;x=-236460000;
#10;x=-236450000;
#10;x=-236440000;
#10;x=-236430000;
#10;x=-236420000;
#10;x=-236410000;
#10;x=-236400000;
#10;x=-236390000;
#10;x=-236380000;
#10;x=-236370000;
#10;x=-236360000;
#10;x=-236350000;
#10;x=-236340000;
#10;x=-236330000;
#10;x=-236320000;
#10;x=-236310000;
#10;x=-236300000;
#10;x=-236290000;
#10;x=-236280000;
#10;x=-236270000;
#10;x=-236260000;
#10;x=-236250000;
#10;x=-236240000;
#10;x=-236230000;
#10;x=-236220000;
#10;x=-236210000;
#10;x=-236200000;
#10;x=-236190000;
#10;x=-236180000;
#10;x=-236170000;
#10;x=-236160000;
#10;x=-236150000;
#10;x=-236140000;
#10;x=-236130000;
#10;x=-236120000;
#10;x=-236110000;
#10;x=-236100000;
#10;x=-236090000;
#10;x=-236080000;
#10;x=-236070000;
#10;x=-236060000;
#10;x=-236050000;
#10;x=-236040000;
#10;x=-236030000;
#10;x=-236020000;
#10;x=-236010000;
#10;x=-236000000;
#10;x=-235990000;
#10;x=-235980000;
#10;x=-235970000;
#10;x=-235960000;
#10;x=-235950000;
#10;x=-235940000;
#10;x=-235930000;
#10;x=-235920000;
#10;x=-235910000;
#10;x=-235900000;
#10;x=-235890000;
#10;x=-235880000;
#10;x=-235870000;
#10;x=-235860000;
#10;x=-235850000;
#10;x=-235840000;
#10;x=-235830000;
#10;x=-235820000;
#10;x=-235810000;
#10;x=-235800000;
#10;x=-235790000;
#10;x=-235780000;
#10;x=-235770000;
#10;x=-235760000;
#10;x=-235750000;
#10;x=-235740000;
#10;x=-235730000;
#10;x=-235720000;
#10;x=-235710000;
#10;x=-235700000;
#10;x=-235690000;
#10;x=-235680000;
#10;x=-235670000;
#10;x=-235660000;
#10;x=-235650000;
#10;x=-235640000;
#10;x=-235630000;
#10;x=-235620000;
#10;x=-235610000;
#10;x=-235600000;
#10;x=-235590000;
#10;x=-235580000;
#10;x=-235570000;
#10;x=-235560000;
#10;x=-235550000;
#10;x=-235540000;
#10;x=-235530000;
#10;x=-235520000;
#10;x=-235510000;
#10;x=-235500000;
#10;x=-235490000;
#10;x=-235480000;
#10;x=-235470000;
#10;x=-235460000;
#10;x=-235450000;
#10;x=-235440000;
#10;x=-235430000;
#10;x=-235420000;
#10;x=-235410000;
#10;x=-235400000;
#10;x=-235390000;
#10;x=-235380000;
#10;x=-235370000;
#10;x=-235360000;
#10;x=-235350000;
#10;x=-235340000;
#10;x=-235330000;
#10;x=-235320000;
#10;x=-235310000;
#10;x=-235300000;
#10;x=-235290000;
#10;x=-235280000;
#10;x=-235270000;
#10;x=-235260000;
#10;x=-235250000;
#10;x=-235240000;
#10;x=-235230000;
#10;x=-235220000;
#10;x=-235210000;
#10;x=-235200000;
#10;x=-235190000;
#10;x=-235180000;
#10;x=-235170000;
#10;x=-235160000;
#10;x=-235150000;
#10;x=-235140000;
#10;x=-235130000;
#10;x=-235120000;
#10;x=-235110000;
#10;x=-235100000;
#10;x=-235090000;
#10;x=-235080000;
#10;x=-235070000;
#10;x=-235060000;
#10;x=-235050000;
#10;x=-235040000;
#10;x=-235030000;
#10;x=-235020000;
#10;x=-235010000;
#10;x=-235000000;
#10;x=-234990000;
#10;x=-234980000;
#10;x=-234970000;
#10;x=-234960000;
#10;x=-234950000;
#10;x=-234940000;
#10;x=-234930000;
#10;x=-234920000;
#10;x=-234910000;
#10;x=-234900000;
#10;x=-234890000;
#10;x=-234880000;
#10;x=-234870000;
#10;x=-234860000;
#10;x=-234850000;
#10;x=-234840000;
#10;x=-234830000;
#10;x=-234820000;
#10;x=-234810000;
#10;x=-234800000;
#10;x=-234790000;
#10;x=-234780000;
#10;x=-234770000;
#10;x=-234760000;
#10;x=-234750000;
#10;x=-234740000;
#10;x=-234730000;
#10;x=-234720000;
#10;x=-234710000;
#10;x=-234700000;
#10;x=-234690000;
#10;x=-234680000;
#10;x=-234670000;
#10;x=-234660000;
#10;x=-234650000;
#10;x=-234640000;
#10;x=-234630000;
#10;x=-234620000;
#10;x=-234610000;
#10;x=-234600000;
#10;x=-234590000;
#10;x=-234580000;
#10;x=-234570000;
#10;x=-234560000;
#10;x=-234550000;
#10;x=-234540000;
#10;x=-234530000;
#10;x=-234520000;
#10;x=-234510000;
#10;x=-234500000;
#10;x=-234490000;
#10;x=-234480000;
#10;x=-234470000;
#10;x=-234460000;
#10;x=-234450000;
#10;x=-234440000;
#10;x=-234430000;
#10;x=-234420000;
#10;x=-234410000;
#10;x=-234400000;
#10;x=-234390000;
#10;x=-234380000;
#10;x=-234370000;
#10;x=-234360000;
#10;x=-234350000;
#10;x=-234340000;
#10;x=-234330000;
#10;x=-234320000;
#10;x=-234310000;
#10;x=-234300000;
#10;x=-234290000;
#10;x=-234280000;
#10;x=-234270000;
#10;x=-234260000;
#10;x=-234250000;
#10;x=-234240000;
#10;x=-234230000;
#10;x=-234220000;
#10;x=-234210000;
#10;x=-234200000;
#10;x=-234190000;
#10;x=-234180000;
#10;x=-234170000;
#10;x=-234160000;
#10;x=-234150000;
#10;x=-234140000;
#10;x=-234130000;
#10;x=-234120000;
#10;x=-234110000;
#10;x=-234100000;
#10;x=-234090000;
#10;x=-234080000;
#10;x=-234070000;
#10;x=-234060000;
#10;x=-234050000;
#10;x=-234040000;
#10;x=-234030000;
#10;x=-234020000;
#10;x=-234010000;
#10;x=-234000000;
#10;x=-233990000;
#10;x=-233980000;
#10;x=-233970000;
#10;x=-233960000;
#10;x=-233950000;
#10;x=-233940000;
#10;x=-233930000;
#10;x=-233920000;
#10;x=-233910000;
#10;x=-233900000;
#10;x=-233890000;
#10;x=-233880000;
#10;x=-233870000;
#10;x=-233860000;
#10;x=-233850000;
#10;x=-233840000;
#10;x=-233830000;
#10;x=-233820000;
#10;x=-233810000;
#10;x=-233800000;
#10;x=-233790000;
#10;x=-233780000;
#10;x=-233770000;
#10;x=-233760000;
#10;x=-233750000;
#10;x=-233740000;
#10;x=-233730000;
#10;x=-233720000;
#10;x=-233710000;
#10;x=-233700000;
#10;x=-233690000;
#10;x=-233680000;
#10;x=-233670000;
#10;x=-233660000;
#10;x=-233650000;
#10;x=-233640000;
#10;x=-233630000;
#10;x=-233620000;
#10;x=-233610000;
#10;x=-233600000;
#10;x=-233590000;
#10;x=-233580000;
#10;x=-233570000;
#10;x=-233560000;
#10;x=-233550000;
#10;x=-233540000;
#10;x=-233530000;
#10;x=-233520000;
#10;x=-233510000;
#10;x=-233500000;
#10;x=-233490000;
#10;x=-233480000;
#10;x=-233470000;
#10;x=-233460000;
#10;x=-233450000;
#10;x=-233440000;
#10;x=-233430000;
#10;x=-233420000;
#10;x=-233410000;
#10;x=-233400000;
#10;x=-233390000;
#10;x=-233380000;
#10;x=-233370000;
#10;x=-233360000;
#10;x=-233350000;
#10;x=-233340000;
#10;x=-233330000;
#10;x=-233320000;
#10;x=-233310000;
#10;x=-233300000;
#10;x=-233290000;
#10;x=-233280000;
#10;x=-233270000;
#10;x=-233260000;
#10;x=-233250000;
#10;x=-233240000;
#10;x=-233230000;
#10;x=-233220000;
#10;x=-233210000;
#10;x=-233200000;
#10;x=-233190000;
#10;x=-233180000;
#10;x=-233170000;
#10;x=-233160000;
#10;x=-233150000;
#10;x=-233140000;
#10;x=-233130000;
#10;x=-233120000;
#10;x=-233110000;
#10;x=-233100000;
#10;x=-233090000;
#10;x=-233080000;
#10;x=-233070000;
#10;x=-233060000;
#10;x=-233050000;
#10;x=-233040000;
#10;x=-233030000;
#10;x=-233020000;
#10;x=-233010000;
#10;x=-233000000;
#10;x=-232990000;
#10;x=-232980000;
#10;x=-232970000;
#10;x=-232960000;
#10;x=-232950000;
#10;x=-232940000;
#10;x=-232930000;
#10;x=-232920000;
#10;x=-232910000;
#10;x=-232900000;
#10;x=-232890000;
#10;x=-232880000;
#10;x=-232870000;
#10;x=-232860000;
#10;x=-232850000;
#10;x=-232840000;
#10;x=-232830000;
#10;x=-232820000;
#10;x=-232810000;
#10;x=-232800000;
#10;x=-232790000;
#10;x=-232780000;
#10;x=-232770000;
#10;x=-232760000;
#10;x=-232750000;
#10;x=-232740000;
#10;x=-232730000;
#10;x=-232720000;
#10;x=-232710000;
#10;x=-232700000;
#10;x=-232690000;
#10;x=-232680000;
#10;x=-232670000;
#10;x=-232660000;
#10;x=-232650000;
#10;x=-232640000;
#10;x=-232630000;
#10;x=-232620000;
#10;x=-232610000;
#10;x=-232600000;
#10;x=-232590000;
#10;x=-232580000;
#10;x=-232570000;
#10;x=-232560000;
#10;x=-232550000;
#10;x=-232540000;
#10;x=-232530000;
#10;x=-232520000;
#10;x=-232510000;
#10;x=-232500000;
#10;x=-232490000;
#10;x=-232480000;
#10;x=-232470000;
#10;x=-232460000;
#10;x=-232450000;
#10;x=-232440000;
#10;x=-232430000;
#10;x=-232420000;
#10;x=-232410000;
#10;x=-232400000;
#10;x=-232390000;
#10;x=-232380000;
#10;x=-232370000;
#10;x=-232360000;
#10;x=-232350000;
#10;x=-232340000;
#10;x=-232330000;
#10;x=-232320000;
#10;x=-232310000;
#10;x=-232300000;
#10;x=-232290000;
#10;x=-232280000;
#10;x=-232270000;
#10;x=-232260000;
#10;x=-232250000;
#10;x=-232240000;
#10;x=-232230000;
#10;x=-232220000;
#10;x=-232210000;
#10;x=-232200000;
#10;x=-232190000;
#10;x=-232180000;
#10;x=-232170000;
#10;x=-232160000;
#10;x=-232150000;
#10;x=-232140000;
#10;x=-232130000;
#10;x=-232120000;
#10;x=-232110000;
#10;x=-232100000;
#10;x=-232090000;
#10;x=-232080000;
#10;x=-232070000;
#10;x=-232060000;
#10;x=-232050000;
#10;x=-232040000;
#10;x=-232030000;
#10;x=-232020000;
#10;x=-232010000;
#10;x=-232000000;
#10;x=-231990000;
#10;x=-231980000;
#10;x=-231970000;
#10;x=-231960000;
#10;x=-231950000;
#10;x=-231940000;
#10;x=-231930000;
#10;x=-231920000;
#10;x=-231910000;
#10;x=-231900000;
#10;x=-231890000;
#10;x=-231880000;
#10;x=-231870000;
#10;x=-231860000;
#10;x=-231850000;
#10;x=-231840000;
#10;x=-231830000;
#10;x=-231820000;
#10;x=-231810000;
#10;x=-231800000;
#10;x=-231790000;
#10;x=-231780000;
#10;x=-231770000;
#10;x=-231760000;
#10;x=-231750000;
#10;x=-231740000;
#10;x=-231730000;
#10;x=-231720000;
#10;x=-231710000;
#10;x=-231700000;
#10;x=-231690000;
#10;x=-231680000;
#10;x=-231670000;
#10;x=-231660000;
#10;x=-231650000;
#10;x=-231640000;
#10;x=-231630000;
#10;x=-231620000;
#10;x=-231610000;
#10;x=-231600000;
#10;x=-231590000;
#10;x=-231580000;
#10;x=-231570000;
#10;x=-231560000;
#10;x=-231550000;
#10;x=-231540000;
#10;x=-231530000;
#10;x=-231520000;
#10;x=-231510000;
#10;x=-231500000;
#10;x=-231490000;
#10;x=-231480000;
#10;x=-231470000;
#10;x=-231460000;
#10;x=-231450000;
#10;x=-231440000;
#10;x=-231430000;
#10;x=-231420000;
#10;x=-231410000;
#10;x=-231400000;
#10;x=-231390000;
#10;x=-231380000;
#10;x=-231370000;
#10;x=-231360000;
#10;x=-231350000;
#10;x=-231340000;
#10;x=-231330000;
#10;x=-231320000;
#10;x=-231310000;
#10;x=-231300000;
#10;x=-231290000;
#10;x=-231280000;
#10;x=-231270000;
#10;x=-231260000;
#10;x=-231250000;
#10;x=-231240000;
#10;x=-231230000;
#10;x=-231220000;
#10;x=-231210000;
#10;x=-231200000;
#10;x=-231190000;
#10;x=-231180000;
#10;x=-231170000;
#10;x=-231160000;
#10;x=-231150000;
#10;x=-231140000;
#10;x=-231130000;
#10;x=-231120000;
#10;x=-231110000;
#10;x=-231100000;
#10;x=-231090000;
#10;x=-231080000;
#10;x=-231070000;
#10;x=-231060000;
#10;x=-231050000;
#10;x=-231040000;
#10;x=-231030000;
#10;x=-231020000;
#10;x=-231010000;
#10;x=-231000000;
#10;x=-230990000;
#10;x=-230980000;
#10;x=-230970000;
#10;x=-230960000;
#10;x=-230950000;
#10;x=-230940000;
#10;x=-230930000;
#10;x=-230920000;
#10;x=-230910000;
#10;x=-230900000;
#10;x=-230890000;
#10;x=-230880000;
#10;x=-230870000;
#10;x=-230860000;
#10;x=-230850000;
#10;x=-230840000;
#10;x=-230830000;
#10;x=-230820000;
#10;x=-230810000;
#10;x=-230800000;
#10;x=-230790000;
#10;x=-230780000;
#10;x=-230770000;
#10;x=-230760000;
#10;x=-230750000;
#10;x=-230740000;
#10;x=-230730000;
#10;x=-230720000;
#10;x=-230710000;
#10;x=-230700000;
#10;x=-230690000;
#10;x=-230680000;
#10;x=-230670000;
#10;x=-230660000;
#10;x=-230650000;
#10;x=-230640000;
#10;x=-230630000;
#10;x=-230620000;
#10;x=-230610000;
#10;x=-230600000;
#10;x=-230590000;
#10;x=-230580000;
#10;x=-230570000;
#10;x=-230560000;
#10;x=-230550000;
#10;x=-230540000;
#10;x=-230530000;
#10;x=-230520000;
#10;x=-230510000;
#10;x=-230500000;
#10;x=-230490000;
#10;x=-230480000;
#10;x=-230470000;
#10;x=-230460000;
#10;x=-230450000;
#10;x=-230440000;
#10;x=-230430000;
#10;x=-230420000;
#10;x=-230410000;
#10;x=-230400000;
#10;x=-230390000;
#10;x=-230380000;
#10;x=-230370000;
#10;x=-230360000;
#10;x=-230350000;
#10;x=-230340000;
#10;x=-230330000;
#10;x=-230320000;
#10;x=-230310000;
#10;x=-230300000;
#10;x=-230290000;
#10;x=-230280000;
#10;x=-230270000;
#10;x=-230260000;
#10;x=-230250000;
#10;x=-230240000;
#10;x=-230230000;
#10;x=-230220000;
#10;x=-230210000;
#10;x=-230200000;
#10;x=-230190000;
#10;x=-230180000;
#10;x=-230170000;
#10;x=-230160000;
#10;x=-230150000;
#10;x=-230140000;
#10;x=-230130000;
#10;x=-230120000;
#10;x=-230110000;
#10;x=-230100000;
#10;x=-230090000;
#10;x=-230080000;
#10;x=-230070000;
#10;x=-230060000;
#10;x=-230050000;
#10;x=-230040000;
#10;x=-230030000;
#10;x=-230020000;
#10;x=-230010000;
#10;x=-230000000;
#10;x=-229990000;
#10;x=-229980000;
#10;x=-229970000;
#10;x=-229960000;
#10;x=-229950000;
#10;x=-229940000;
#10;x=-229930000;
#10;x=-229920000;
#10;x=-229910000;
#10;x=-229900000;
#10;x=-229890000;
#10;x=-229880000;
#10;x=-229870000;
#10;x=-229860000;
#10;x=-229850000;
#10;x=-229840000;
#10;x=-229830000;
#10;x=-229820000;
#10;x=-229810000;
#10;x=-229800000;
#10;x=-229790000;
#10;x=-229780000;
#10;x=-229770000;
#10;x=-229760000;
#10;x=-229750000;
#10;x=-229740000;
#10;x=-229730000;
#10;x=-229720000;
#10;x=-229710000;
#10;x=-229700000;
#10;x=-229690000;
#10;x=-229680000;
#10;x=-229670000;
#10;x=-229660000;
#10;x=-229650000;
#10;x=-229640000;
#10;x=-229630000;
#10;x=-229620000;
#10;x=-229610000;
#10;x=-229600000;
#10;x=-229590000;
#10;x=-229580000;
#10;x=-229570000;
#10;x=-229560000;
#10;x=-229550000;
#10;x=-229540000;
#10;x=-229530000;
#10;x=-229520000;
#10;x=-229510000;
#10;x=-229500000;
#10;x=-229490000;
#10;x=-229480000;
#10;x=-229470000;
#10;x=-229460000;
#10;x=-229450000;
#10;x=-229440000;
#10;x=-229430000;
#10;x=-229420000;
#10;x=-229410000;
#10;x=-229400000;
#10;x=-229390000;
#10;x=-229380000;
#10;x=-229370000;
#10;x=-229360000;
#10;x=-229350000;
#10;x=-229340000;
#10;x=-229330000;
#10;x=-229320000;
#10;x=-229310000;
#10;x=-229300000;
#10;x=-229290000;
#10;x=-229280000;
#10;x=-229270000;
#10;x=-229260000;
#10;x=-229250000;
#10;x=-229240000;
#10;x=-229230000;
#10;x=-229220000;
#10;x=-229210000;
#10;x=-229200000;
#10;x=-229190000;
#10;x=-229180000;
#10;x=-229170000;
#10;x=-229160000;
#10;x=-229150000;
#10;x=-229140000;
#10;x=-229130000;
#10;x=-229120000;
#10;x=-229110000;
#10;x=-229100000;
#10;x=-229090000;
#10;x=-229080000;
#10;x=-229070000;
#10;x=-229060000;
#10;x=-229050000;
#10;x=-229040000;
#10;x=-229030000;
#10;x=-229020000;
#10;x=-229010000;
#10;x=-229000000;
#10;x=-228990000;
#10;x=-228980000;
#10;x=-228970000;
#10;x=-228960000;
#10;x=-228950000;
#10;x=-228940000;
#10;x=-228930000;
#10;x=-228920000;
#10;x=-228910000;
#10;x=-228900000;
#10;x=-228890000;
#10;x=-228880000;
#10;x=-228870000;
#10;x=-228860000;
#10;x=-228850000;
#10;x=-228840000;
#10;x=-228830000;
#10;x=-228820000;
#10;x=-228810000;
#10;x=-228800000;
#10;x=-228790000;
#10;x=-228780000;
#10;x=-228770000;
#10;x=-228760000;
#10;x=-228750000;
#10;x=-228740000;
#10;x=-228730000;
#10;x=-228720000;
#10;x=-228710000;
#10;x=-228700000;
#10;x=-228690000;
#10;x=-228680000;
#10;x=-228670000;
#10;x=-228660000;
#10;x=-228650000;
#10;x=-228640000;
#10;x=-228630000;
#10;x=-228620000;
#10;x=-228610000;
#10;x=-228600000;
#10;x=-228590000;
#10;x=-228580000;
#10;x=-228570000;
#10;x=-228560000;
#10;x=-228550000;
#10;x=-228540000;
#10;x=-228530000;
#10;x=-228520000;
#10;x=-228510000;
#10;x=-228500000;
#10;x=-228490000;
#10;x=-228480000;
#10;x=-228470000;
#10;x=-228460000;
#10;x=-228450000;
#10;x=-228440000;
#10;x=-228430000;
#10;x=-228420000;
#10;x=-228410000;
#10;x=-228400000;
#10;x=-228390000;
#10;x=-228380000;
#10;x=-228370000;
#10;x=-228360000;
#10;x=-228350000;
#10;x=-228340000;
#10;x=-228330000;
#10;x=-228320000;
#10;x=-228310000;
#10;x=-228300000;
#10;x=-228290000;
#10;x=-228280000;
#10;x=-228270000;
#10;x=-228260000;
#10;x=-228250000;
#10;x=-228240000;
#10;x=-228230000;
#10;x=-228220000;
#10;x=-228210000;
#10;x=-228200000;
#10;x=-228190000;
#10;x=-228180000;
#10;x=-228170000;
#10;x=-228160000;
#10;x=-228150000;
#10;x=-228140000;
#10;x=-228130000;
#10;x=-228120000;
#10;x=-228110000;
#10;x=-228100000;
#10;x=-228090000;
#10;x=-228080000;
#10;x=-228070000;
#10;x=-228060000;
#10;x=-228050000;
#10;x=-228040000;
#10;x=-228030000;
#10;x=-228020000;
#10;x=-228010000;
#10;x=-228000000;
#10;x=-227990000;
#10;x=-227980000;
#10;x=-227970000;
#10;x=-227960000;
#10;x=-227950000;
#10;x=-227940000;
#10;x=-227930000;
#10;x=-227920000;
#10;x=-227910000;
#10;x=-227900000;
#10;x=-227890000;
#10;x=-227880000;
#10;x=-227870000;
#10;x=-227860000;
#10;x=-227850000;
#10;x=-227840000;
#10;x=-227830000;
#10;x=-227820000;
#10;x=-227810000;
#10;x=-227800000;
#10;x=-227790000;
#10;x=-227780000;
#10;x=-227770000;
#10;x=-227760000;
#10;x=-227750000;
#10;x=-227740000;
#10;x=-227730000;
#10;x=-227720000;
#10;x=-227710000;
#10;x=-227700000;
#10;x=-227690000;
#10;x=-227680000;
#10;x=-227670000;
#10;x=-227660000;
#10;x=-227650000;
#10;x=-227640000;
#10;x=-227630000;
#10;x=-227620000;
#10;x=-227610000;
#10;x=-227600000;
#10;x=-227590000;
#10;x=-227580000;
#10;x=-227570000;
#10;x=-227560000;
#10;x=-227550000;
#10;x=-227540000;
#10;x=-227530000;
#10;x=-227520000;
#10;x=-227510000;
#10;x=-227500000;
#10;x=-227490000;
#10;x=-227480000;
#10;x=-227470000;
#10;x=-227460000;
#10;x=-227450000;
#10;x=-227440000;
#10;x=-227430000;
#10;x=-227420000;
#10;x=-227410000;
#10;x=-227400000;
#10;x=-227390000;
#10;x=-227380000;
#10;x=-227370000;
#10;x=-227360000;
#10;x=-227350000;
#10;x=-227340000;
#10;x=-227330000;
#10;x=-227320000;
#10;x=-227310000;
#10;x=-227300000;
#10;x=-227290000;
#10;x=-227280000;
#10;x=-227270000;
#10;x=-227260000;
#10;x=-227250000;
#10;x=-227240000;
#10;x=-227230000;
#10;x=-227220000;
#10;x=-227210000;
#10;x=-227200000;
#10;x=-227190000;
#10;x=-227180000;
#10;x=-227170000;
#10;x=-227160000;
#10;x=-227150000;
#10;x=-227140000;
#10;x=-227130000;
#10;x=-227120000;
#10;x=-227110000;
#10;x=-227100000;
#10;x=-227090000;
#10;x=-227080000;
#10;x=-227070000;
#10;x=-227060000;
#10;x=-227050000;
#10;x=-227040000;
#10;x=-227030000;
#10;x=-227020000;
#10;x=-227010000;
#10;x=-227000000;
#10;x=-226990000;
#10;x=-226980000;
#10;x=-226970000;
#10;x=-226960000;
#10;x=-226950000;
#10;x=-226940000;
#10;x=-226930000;
#10;x=-226920000;
#10;x=-226910000;
#10;x=-226900000;
#10;x=-226890000;
#10;x=-226880000;
#10;x=-226870000;
#10;x=-226860000;
#10;x=-226850000;
#10;x=-226840000;
#10;x=-226830000;
#10;x=-226820000;
#10;x=-226810000;
#10;x=-226800000;
#10;x=-226790000;
#10;x=-226780000;
#10;x=-226770000;
#10;x=-226760000;
#10;x=-226750000;
#10;x=-226740000;
#10;x=-226730000;
#10;x=-226720000;
#10;x=-226710000;
#10;x=-226700000;
#10;x=-226690000;
#10;x=-226680000;
#10;x=-226670000;
#10;x=-226660000;
#10;x=-226650000;
#10;x=-226640000;
#10;x=-226630000;
#10;x=-226620000;
#10;x=-226610000;
#10;x=-226600000;
#10;x=-226590000;
#10;x=-226580000;
#10;x=-226570000;
#10;x=-226560000;
#10;x=-226550000;
#10;x=-226540000;
#10;x=-226530000;
#10;x=-226520000;
#10;x=-226510000;
#10;x=-226500000;
#10;x=-226490000;
#10;x=-226480000;
#10;x=-226470000;
#10;x=-226460000;
#10;x=-226450000;
#10;x=-226440000;
#10;x=-226430000;
#10;x=-226420000;
#10;x=-226410000;
#10;x=-226400000;
#10;x=-226390000;
#10;x=-226380000;
#10;x=-226370000;
#10;x=-226360000;
#10;x=-226350000;
#10;x=-226340000;
#10;x=-226330000;
#10;x=-226320000;
#10;x=-226310000;
#10;x=-226300000;
#10;x=-226290000;
#10;x=-226280000;
#10;x=-226270000;
#10;x=-226260000;
#10;x=-226250000;
#10;x=-226240000;
#10;x=-226230000;
#10;x=-226220000;
#10;x=-226210000;
#10;x=-226200000;
#10;x=-226190000;
#10;x=-226180000;
#10;x=-226170000;
#10;x=-226160000;
#10;x=-226150000;
#10;x=-226140000;
#10;x=-226130000;
#10;x=-226120000;
#10;x=-226110000;
#10;x=-226100000;
#10;x=-226090000;
#10;x=-226080000;
#10;x=-226070000;
#10;x=-226060000;
#10;x=-226050000;
#10;x=-226040000;
#10;x=-226030000;
#10;x=-226020000;
#10;x=-226010000;
#10;x=-226000000;
#10;x=-225990000;
#10;x=-225980000;
#10;x=-225970000;
#10;x=-225960000;
#10;x=-225950000;
#10;x=-225940000;
#10;x=-225930000;
#10;x=-225920000;
#10;x=-225910000;
#10;x=-225900000;
#10;x=-225890000;
#10;x=-225880000;
#10;x=-225870000;
#10;x=-225860000;
#10;x=-225850000;
#10;x=-225840000;
#10;x=-225830000;
#10;x=-225820000;
#10;x=-225810000;
#10;x=-225800000;
#10;x=-225790000;
#10;x=-225780000;
#10;x=-225770000;
#10;x=-225760000;
#10;x=-225750000;
#10;x=-225740000;
#10;x=-225730000;
#10;x=-225720000;
#10;x=-225710000;
#10;x=-225700000;
#10;x=-225690000;
#10;x=-225680000;
#10;x=-225670000;
#10;x=-225660000;
#10;x=-225650000;
#10;x=-225640000;
#10;x=-225630000;
#10;x=-225620000;
#10;x=-225610000;
#10;x=-225600000;
#10;x=-225590000;
#10;x=-225580000;
#10;x=-225570000;
#10;x=-225560000;
#10;x=-225550000;
#10;x=-225540000;
#10;x=-225530000;
#10;x=-225520000;
#10;x=-225510000;
#10;x=-225500000;
#10;x=-225490000;
#10;x=-225480000;
#10;x=-225470000;
#10;x=-225460000;
#10;x=-225450000;
#10;x=-225440000;
#10;x=-225430000;
#10;x=-225420000;
#10;x=-225410000;
#10;x=-225400000;
#10;x=-225390000;
#10;x=-225380000;
#10;x=-225370000;
#10;x=-225360000;
#10;x=-225350000;
#10;x=-225340000;
#10;x=-225330000;
#10;x=-225320000;
#10;x=-225310000;
#10;x=-225300000;
#10;x=-225290000;
#10;x=-225280000;
#10;x=-225270000;
#10;x=-225260000;
#10;x=-225250000;
#10;x=-225240000;
#10;x=-225230000;
#10;x=-225220000;
#10;x=-225210000;
#10;x=-225200000;
#10;x=-225190000;
#10;x=-225180000;
#10;x=-225170000;
#10;x=-225160000;
#10;x=-225150000;
#10;x=-225140000;
#10;x=-225130000;
#10;x=-225120000;
#10;x=-225110000;
#10;x=-225100000;
#10;x=-225090000;
#10;x=-225080000;
#10;x=-225070000;
#10;x=-225060000;
#10;x=-225050000;
#10;x=-225040000;
#10;x=-225030000;
#10;x=-225020000;
#10;x=-225010000;
#10;x=-225000000;
#10;x=-224990000;
#10;x=-224980000;
#10;x=-224970000;
#10;x=-224960000;
#10;x=-224950000;
#10;x=-224940000;
#10;x=-224930000;
#10;x=-224920000;
#10;x=-224910000;
#10;x=-224900000;
#10;x=-224890000;
#10;x=-224880000;
#10;x=-224870000;
#10;x=-224860000;
#10;x=-224850000;
#10;x=-224840000;
#10;x=-224830000;
#10;x=-224820000;
#10;x=-224810000;
#10;x=-224800000;
#10;x=-224790000;
#10;x=-224780000;
#10;x=-224770000;
#10;x=-224760000;
#10;x=-224750000;
#10;x=-224740000;
#10;x=-224730000;
#10;x=-224720000;
#10;x=-224710000;
#10;x=-224700000;
#10;x=-224690000;
#10;x=-224680000;
#10;x=-224670000;
#10;x=-224660000;
#10;x=-224650000;
#10;x=-224640000;
#10;x=-224630000;
#10;x=-224620000;
#10;x=-224610000;
#10;x=-224600000;
#10;x=-224590000;
#10;x=-224580000;
#10;x=-224570000;
#10;x=-224560000;
#10;x=-224550000;
#10;x=-224540000;
#10;x=-224530000;
#10;x=-224520000;
#10;x=-224510000;
#10;x=-224500000;
#10;x=-224490000;
#10;x=-224480000;
#10;x=-224470000;
#10;x=-224460000;
#10;x=-224450000;
#10;x=-224440000;
#10;x=-224430000;
#10;x=-224420000;
#10;x=-224410000;
#10;x=-224400000;
#10;x=-224390000;
#10;x=-224380000;
#10;x=-224370000;
#10;x=-224360000;
#10;x=-224350000;
#10;x=-224340000;
#10;x=-224330000;
#10;x=-224320000;
#10;x=-224310000;
#10;x=-224300000;
#10;x=-224290000;
#10;x=-224280000;
#10;x=-224270000;
#10;x=-224260000;
#10;x=-224250000;
#10;x=-224240000;
#10;x=-224230000;
#10;x=-224220000;
#10;x=-224210000;
#10;x=-224200000;
#10;x=-224190000;
#10;x=-224180000;
#10;x=-224170000;
#10;x=-224160000;
#10;x=-224150000;
#10;x=-224140000;
#10;x=-224130000;
#10;x=-224120000;
#10;x=-224110000;
#10;x=-224100000;
#10;x=-224090000;
#10;x=-224080000;
#10;x=-224070000;
#10;x=-224060000;
#10;x=-224050000;
#10;x=-224040000;
#10;x=-224030000;
#10;x=-224020000;
#10;x=-224010000;
#10;x=-224000000;
#10;x=-223990000;
#10;x=-223980000;
#10;x=-223970000;
#10;x=-223960000;
#10;x=-223950000;
#10;x=-223940000;
#10;x=-223930000;
#10;x=-223920000;
#10;x=-223910000;
#10;x=-223900000;
#10;x=-223890000;
#10;x=-223880000;
#10;x=-223870000;
#10;x=-223860000;
#10;x=-223850000;
#10;x=-223840000;
#10;x=-223830000;
#10;x=-223820000;
#10;x=-223810000;
#10;x=-223800000;
#10;x=-223790000;
#10;x=-223780000;
#10;x=-223770000;
#10;x=-223760000;
#10;x=-223750000;
#10;x=-223740000;
#10;x=-223730000;
#10;x=-223720000;
#10;x=-223710000;
#10;x=-223700000;
#10;x=-223690000;
#10;x=-223680000;
#10;x=-223670000;
#10;x=-223660000;
#10;x=-223650000;
#10;x=-223640000;
#10;x=-223630000;
#10;x=-223620000;
#10;x=-223610000;
#10;x=-223600000;
#10;x=-223590000;
#10;x=-223580000;
#10;x=-223570000;
#10;x=-223560000;
#10;x=-223550000;
#10;x=-223540000;
#10;x=-223530000;
#10;x=-223520000;
#10;x=-223510000;
#10;x=-223500000;
#10;x=-223490000;
#10;x=-223480000;
#10;x=-223470000;
#10;x=-223460000;
#10;x=-223450000;
#10;x=-223440000;
#10;x=-223430000;
#10;x=-223420000;
#10;x=-223410000;
#10;x=-223400000;
#10;x=-223390000;
#10;x=-223380000;
#10;x=-223370000;
#10;x=-223360000;
#10;x=-223350000;
#10;x=-223340000;
#10;x=-223330000;
#10;x=-223320000;
#10;x=-223310000;
#10;x=-223300000;
#10;x=-223290000;
#10;x=-223280000;
#10;x=-223270000;
#10;x=-223260000;
#10;x=-223250000;
#10;x=-223240000;
#10;x=-223230000;
#10;x=-223220000;
#10;x=-223210000;
#10;x=-223200000;
#10;x=-223190000;
#10;x=-223180000;
#10;x=-223170000;
#10;x=-223160000;
#10;x=-223150000;
#10;x=-223140000;
#10;x=-223130000;
#10;x=-223120000;
#10;x=-223110000;
#10;x=-223100000;
#10;x=-223090000;
#10;x=-223080000;
#10;x=-223070000;
#10;x=-223060000;
#10;x=-223050000;
#10;x=-223040000;
#10;x=-223030000;
#10;x=-223020000;
#10;x=-223010000;
#10;x=-223000000;
#10;x=-222990000;
#10;x=-222980000;
#10;x=-222970000;
#10;x=-222960000;
#10;x=-222950000;
#10;x=-222940000;
#10;x=-222930000;
#10;x=-222920000;
#10;x=-222910000;
#10;x=-222900000;
#10;x=-222890000;
#10;x=-222880000;
#10;x=-222870000;
#10;x=-222860000;
#10;x=-222850000;
#10;x=-222840000;
#10;x=-222830000;
#10;x=-222820000;
#10;x=-222810000;
#10;x=-222800000;
#10;x=-222790000;
#10;x=-222780000;
#10;x=-222770000;
#10;x=-222760000;
#10;x=-222750000;
#10;x=-222740000;
#10;x=-222730000;
#10;x=-222720000;
#10;x=-222710000;
#10;x=-222700000;
#10;x=-222690000;
#10;x=-222680000;
#10;x=-222670000;
#10;x=-222660000;
#10;x=-222650000;
#10;x=-222640000;
#10;x=-222630000;
#10;x=-222620000;
#10;x=-222610000;
#10;x=-222600000;
#10;x=-222590000;
#10;x=-222580000;
#10;x=-222570000;
#10;x=-222560000;
#10;x=-222550000;
#10;x=-222540000;
#10;x=-222530000;
#10;x=-222520000;
#10;x=-222510000;
#10;x=-222500000;
#10;x=-222490000;
#10;x=-222480000;
#10;x=-222470000;
#10;x=-222460000;
#10;x=-222450000;
#10;x=-222440000;
#10;x=-222430000;
#10;x=-222420000;
#10;x=-222410000;
#10;x=-222400000;
#10;x=-222390000;
#10;x=-222380000;
#10;x=-222370000;
#10;x=-222360000;
#10;x=-222350000;
#10;x=-222340000;
#10;x=-222330000;
#10;x=-222320000;
#10;x=-222310000;
#10;x=-222300000;
#10;x=-222290000;
#10;x=-222280000;
#10;x=-222270000;
#10;x=-222260000;
#10;x=-222250000;
#10;x=-222240000;
#10;x=-222230000;
#10;x=-222220000;
#10;x=-222210000;
#10;x=-222200000;
#10;x=-222190000;
#10;x=-222180000;
#10;x=-222170000;
#10;x=-222160000;
#10;x=-222150000;
#10;x=-222140000;
#10;x=-222130000;
#10;x=-222120000;
#10;x=-222110000;
#10;x=-222100000;
#10;x=-222090000;
#10;x=-222080000;
#10;x=-222070000;
#10;x=-222060000;
#10;x=-222050000;
#10;x=-222040000;
#10;x=-222030000;
#10;x=-222020000;
#10;x=-222010000;
#10;x=-222000000;
#10;x=-221990000;
#10;x=-221980000;
#10;x=-221970000;
#10;x=-221960000;
#10;x=-221950000;
#10;x=-221940000;
#10;x=-221930000;
#10;x=-221920000;
#10;x=-221910000;
#10;x=-221900000;
#10;x=-221890000;
#10;x=-221880000;
#10;x=-221870000;
#10;x=-221860000;
#10;x=-221850000;
#10;x=-221840000;
#10;x=-221830000;
#10;x=-221820000;
#10;x=-221810000;
#10;x=-221800000;
#10;x=-221790000;
#10;x=-221780000;
#10;x=-221770000;
#10;x=-221760000;
#10;x=-221750000;
#10;x=-221740000;
#10;x=-221730000;
#10;x=-221720000;
#10;x=-221710000;
#10;x=-221700000;
#10;x=-221690000;
#10;x=-221680000;
#10;x=-221670000;
#10;x=-221660000;
#10;x=-221650000;
#10;x=-221640000;
#10;x=-221630000;
#10;x=-221620000;
#10;x=-221610000;
#10;x=-221600000;
#10;x=-221590000;
#10;x=-221580000;
#10;x=-221570000;
#10;x=-221560000;
#10;x=-221550000;
#10;x=-221540000;
#10;x=-221530000;
#10;x=-221520000;
#10;x=-221510000;
#10;x=-221500000;
#10;x=-221490000;
#10;x=-221480000;
#10;x=-221470000;
#10;x=-221460000;
#10;x=-221450000;
#10;x=-221440000;
#10;x=-221430000;
#10;x=-221420000;
#10;x=-221410000;
#10;x=-221400000;
#10;x=-221390000;
#10;x=-221380000;
#10;x=-221370000;
#10;x=-221360000;
#10;x=-221350000;
#10;x=-221340000;
#10;x=-221330000;
#10;x=-221320000;
#10;x=-221310000;
#10;x=-221300000;
#10;x=-221290000;
#10;x=-221280000;
#10;x=-221270000;
#10;x=-221260000;
#10;x=-221250000;
#10;x=-221240000;
#10;x=-221230000;
#10;x=-221220000;
#10;x=-221210000;
#10;x=-221200000;
#10;x=-221190000;
#10;x=-221180000;
#10;x=-221170000;
#10;x=-221160000;
#10;x=-221150000;
#10;x=-221140000;
#10;x=-221130000;
#10;x=-221120000;
#10;x=-221110000;
#10;x=-221100000;
#10;x=-221090000;
#10;x=-221080000;
#10;x=-221070000;
#10;x=-221060000;
#10;x=-221050000;
#10;x=-221040000;
#10;x=-221030000;
#10;x=-221020000;
#10;x=-221010000;
#10;x=-221000000;
#10;x=-220990000;
#10;x=-220980000;
#10;x=-220970000;
#10;x=-220960000;
#10;x=-220950000;
#10;x=-220940000;
#10;x=-220930000;
#10;x=-220920000;
#10;x=-220910000;
#10;x=-220900000;
#10;x=-220890000;
#10;x=-220880000;
#10;x=-220870000;
#10;x=-220860000;
#10;x=-220850000;
#10;x=-220840000;
#10;x=-220830000;
#10;x=-220820000;
#10;x=-220810000;
#10;x=-220800000;
#10;x=-220790000;
#10;x=-220780000;
#10;x=-220770000;
#10;x=-220760000;
#10;x=-220750000;
#10;x=-220740000;
#10;x=-220730000;
#10;x=-220720000;
#10;x=-220710000;
#10;x=-220700000;
#10;x=-220690000;
#10;x=-220680000;
#10;x=-220670000;
#10;x=-220660000;
#10;x=-220650000;
#10;x=-220640000;
#10;x=-220630000;
#10;x=-220620000;
#10;x=-220610000;
#10;x=-220600000;
#10;x=-220590000;
#10;x=-220580000;
#10;x=-220570000;
#10;x=-220560000;
#10;x=-220550000;
#10;x=-220540000;
#10;x=-220530000;
#10;x=-220520000;
#10;x=-220510000;
#10;x=-220500000;
#10;x=-220490000;
#10;x=-220480000;
#10;x=-220470000;
#10;x=-220460000;
#10;x=-220450000;
#10;x=-220440000;
#10;x=-220430000;
#10;x=-220420000;
#10;x=-220410000;
#10;x=-220400000;
#10;x=-220390000;
#10;x=-220380000;
#10;x=-220370000;
#10;x=-220360000;
#10;x=-220350000;
#10;x=-220340000;
#10;x=-220330000;
#10;x=-220320000;
#10;x=-220310000;
#10;x=-220300000;
#10;x=-220290000;
#10;x=-220280000;
#10;x=-220270000;
#10;x=-220260000;
#10;x=-220250000;
#10;x=-220240000;
#10;x=-220230000;
#10;x=-220220000;
#10;x=-220210000;
#10;x=-220200000;
#10;x=-220190000;
#10;x=-220180000;
#10;x=-220170000;
#10;x=-220160000;
#10;x=-220150000;
#10;x=-220140000;
#10;x=-220130000;
#10;x=-220120000;
#10;x=-220110000;
#10;x=-220100000;
#10;x=-220090000;
#10;x=-220080000;
#10;x=-220070000;
#10;x=-220060000;
#10;x=-220050000;
#10;x=-220040000;
#10;x=-220030000;
#10;x=-220020000;
#10;x=-220010000;
#10;x=-220000000;
#10;x=-219990000;
#10;x=-219980000;
#10;x=-219970000;
#10;x=-219960000;
#10;x=-219950000;
#10;x=-219940000;
#10;x=-219930000;
#10;x=-219920000;
#10;x=-219910000;
#10;x=-219900000;
#10;x=-219890000;
#10;x=-219880000;
#10;x=-219870000;
#10;x=-219860000;
#10;x=-219850000;
#10;x=-219840000;
#10;x=-219830000;
#10;x=-219820000;
#10;x=-219810000;
#10;x=-219800000;
#10;x=-219790000;
#10;x=-219780000;
#10;x=-219770000;
#10;x=-219760000;
#10;x=-219750000;
#10;x=-219740000;
#10;x=-219730000;
#10;x=-219720000;
#10;x=-219710000;
#10;x=-219700000;
#10;x=-219690000;
#10;x=-219680000;
#10;x=-219670000;
#10;x=-219660000;
#10;x=-219650000;
#10;x=-219640000;
#10;x=-219630000;
#10;x=-219620000;
#10;x=-219610000;
#10;x=-219600000;
#10;x=-219590000;
#10;x=-219580000;
#10;x=-219570000;
#10;x=-219560000;
#10;x=-219550000;
#10;x=-219540000;
#10;x=-219530000;
#10;x=-219520000;
#10;x=-219510000;
#10;x=-219500000;
#10;x=-219490000;
#10;x=-219480000;
#10;x=-219470000;
#10;x=-219460000;
#10;x=-219450000;
#10;x=-219440000;
#10;x=-219430000;
#10;x=-219420000;
#10;x=-219410000;
#10;x=-219400000;
#10;x=-219390000;
#10;x=-219380000;
#10;x=-219370000;
#10;x=-219360000;
#10;x=-219350000;
#10;x=-219340000;
#10;x=-219330000;
#10;x=-219320000;
#10;x=-219310000;
#10;x=-219300000;
#10;x=-219290000;
#10;x=-219280000;
#10;x=-219270000;
#10;x=-219260000;
#10;x=-219250000;
#10;x=-219240000;
#10;x=-219230000;
#10;x=-219220000;
#10;x=-219210000;
#10;x=-219200000;
#10;x=-219190000;
#10;x=-219180000;
#10;x=-219170000;
#10;x=-219160000;
#10;x=-219150000;
#10;x=-219140000;
#10;x=-219130000;
#10;x=-219120000;
#10;x=-219110000;
#10;x=-219100000;
#10;x=-219090000;
#10;x=-219080000;
#10;x=-219070000;
#10;x=-219060000;
#10;x=-219050000;
#10;x=-219040000;
#10;x=-219030000;
#10;x=-219020000;
#10;x=-219010000;
#10;x=-219000000;
#10;x=-218990000;
#10;x=-218980000;
#10;x=-218970000;
#10;x=-218960000;
#10;x=-218950000;
#10;x=-218940000;
#10;x=-218930000;
#10;x=-218920000;
#10;x=-218910000;
#10;x=-218900000;
#10;x=-218890000;
#10;x=-218880000;
#10;x=-218870000;
#10;x=-218860000;
#10;x=-218850000;
#10;x=-218840000;
#10;x=-218830000;
#10;x=-218820000;
#10;x=-218810000;
#10;x=-218800000;
#10;x=-218790000;
#10;x=-218780000;
#10;x=-218770000;
#10;x=-218760000;
#10;x=-218750000;
#10;x=-218740000;
#10;x=-218730000;
#10;x=-218720000;
#10;x=-218710000;
#10;x=-218700000;
#10;x=-218690000;
#10;x=-218680000;
#10;x=-218670000;
#10;x=-218660000;
#10;x=-218650000;
#10;x=-218640000;
#10;x=-218630000;
#10;x=-218620000;
#10;x=-218610000;
#10;x=-218600000;
#10;x=-218590000;
#10;x=-218580000;
#10;x=-218570000;
#10;x=-218560000;
#10;x=-218550000;
#10;x=-218540000;
#10;x=-218530000;
#10;x=-218520000;
#10;x=-218510000;
#10;x=-218500000;
#10;x=-218490000;
#10;x=-218480000;
#10;x=-218470000;
#10;x=-218460000;
#10;x=-218450000;
#10;x=-218440000;
#10;x=-218430000;
#10;x=-218420000;
#10;x=-218410000;
#10;x=-218400000;
#10;x=-218390000;
#10;x=-218380000;
#10;x=-218370000;
#10;x=-218360000;
#10;x=-218350000;
#10;x=-218340000;
#10;x=-218330000;
#10;x=-218320000;
#10;x=-218310000;
#10;x=-218300000;
#10;x=-218290000;
#10;x=-218280000;
#10;x=-218270000;
#10;x=-218260000;
#10;x=-218250000;
#10;x=-218240000;
#10;x=-218230000;
#10;x=-218220000;
#10;x=-218210000;
#10;x=-218200000;
#10;x=-218190000;
#10;x=-218180000;
#10;x=-218170000;
#10;x=-218160000;
#10;x=-218150000;
#10;x=-218140000;
#10;x=-218130000;
#10;x=-218120000;
#10;x=-218110000;
#10;x=-218100000;
#10;x=-218090000;
#10;x=-218080000;
#10;x=-218070000;
#10;x=-218060000;
#10;x=-218050000;
#10;x=-218040000;
#10;x=-218030000;
#10;x=-218020000;
#10;x=-218010000;
#10;x=-218000000;
#10;x=-217990000;
#10;x=-217980000;
#10;x=-217970000;
#10;x=-217960000;
#10;x=-217950000;
#10;x=-217940000;
#10;x=-217930000;
#10;x=-217920000;
#10;x=-217910000;
#10;x=-217900000;
#10;x=-217890000;
#10;x=-217880000;
#10;x=-217870000;
#10;x=-217860000;
#10;x=-217850000;
#10;x=-217840000;
#10;x=-217830000;
#10;x=-217820000;
#10;x=-217810000;
#10;x=-217800000;
#10;x=-217790000;
#10;x=-217780000;
#10;x=-217770000;
#10;x=-217760000;
#10;x=-217750000;
#10;x=-217740000;
#10;x=-217730000;
#10;x=-217720000;
#10;x=-217710000;
#10;x=-217700000;
#10;x=-217690000;
#10;x=-217680000;
#10;x=-217670000;
#10;x=-217660000;
#10;x=-217650000;
#10;x=-217640000;
#10;x=-217630000;
#10;x=-217620000;
#10;x=-217610000;
#10;x=-217600000;
#10;x=-217590000;
#10;x=-217580000;
#10;x=-217570000;
#10;x=-217560000;
#10;x=-217550000;
#10;x=-217540000;
#10;x=-217530000;
#10;x=-217520000;
#10;x=-217510000;
#10;x=-217500000;
#10;x=-217490000;
#10;x=-217480000;
#10;x=-217470000;
#10;x=-217460000;
#10;x=-217450000;
#10;x=-217440000;
#10;x=-217430000;
#10;x=-217420000;
#10;x=-217410000;
#10;x=-217400000;
#10;x=-217390000;
#10;x=-217380000;
#10;x=-217370000;
#10;x=-217360000;
#10;x=-217350000;
#10;x=-217340000;
#10;x=-217330000;
#10;x=-217320000;
#10;x=-217310000;
#10;x=-217300000;
#10;x=-217290000;
#10;x=-217280000;
#10;x=-217270000;
#10;x=-217260000;
#10;x=-217250000;
#10;x=-217240000;
#10;x=-217230000;
#10;x=-217220000;
#10;x=-217210000;
#10;x=-217200000;
#10;x=-217190000;
#10;x=-217180000;
#10;x=-217170000;
#10;x=-217160000;
#10;x=-217150000;
#10;x=-217140000;
#10;x=-217130000;
#10;x=-217120000;
#10;x=-217110000;
#10;x=-217100000;
#10;x=-217090000;
#10;x=-217080000;
#10;x=-217070000;
#10;x=-217060000;
#10;x=-217050000;
#10;x=-217040000;
#10;x=-217030000;
#10;x=-217020000;
#10;x=-217010000;
#10;x=-217000000;
#10;x=-216990000;
#10;x=-216980000;
#10;x=-216970000;
#10;x=-216960000;
#10;x=-216950000;
#10;x=-216940000;
#10;x=-216930000;
#10;x=-216920000;
#10;x=-216910000;
#10;x=-216900000;
#10;x=-216890000;
#10;x=-216880000;
#10;x=-216870000;
#10;x=-216860000;
#10;x=-216850000;
#10;x=-216840000;
#10;x=-216830000;
#10;x=-216820000;
#10;x=-216810000;
#10;x=-216800000;
#10;x=-216790000;
#10;x=-216780000;
#10;x=-216770000;
#10;x=-216760000;
#10;x=-216750000;
#10;x=-216740000;
#10;x=-216730000;
#10;x=-216720000;
#10;x=-216710000;
#10;x=-216700000;
#10;x=-216690000;
#10;x=-216680000;
#10;x=-216670000;
#10;x=-216660000;
#10;x=-216650000;
#10;x=-216640000;
#10;x=-216630000;
#10;x=-216620000;
#10;x=-216610000;
#10;x=-216600000;
#10;x=-216590000;
#10;x=-216580000;
#10;x=-216570000;
#10;x=-216560000;
#10;x=-216550000;
#10;x=-216540000;
#10;x=-216530000;
#10;x=-216520000;
#10;x=-216510000;
#10;x=-216500000;
#10;x=-216490000;
#10;x=-216480000;
#10;x=-216470000;
#10;x=-216460000;
#10;x=-216450000;
#10;x=-216440000;
#10;x=-216430000;
#10;x=-216420000;
#10;x=-216410000;
#10;x=-216400000;
#10;x=-216390000;
#10;x=-216380000;
#10;x=-216370000;
#10;x=-216360000;
#10;x=-216350000;
#10;x=-216340000;
#10;x=-216330000;
#10;x=-216320000;
#10;x=-216310000;
#10;x=-216300000;
#10;x=-216290000;
#10;x=-216280000;
#10;x=-216270000;
#10;x=-216260000;
#10;x=-216250000;
#10;x=-216240000;
#10;x=-216230000;
#10;x=-216220000;
#10;x=-216210000;
#10;x=-216200000;
#10;x=-216190000;
#10;x=-216180000;
#10;x=-216170000;
#10;x=-216160000;
#10;x=-216150000;
#10;x=-216140000;
#10;x=-216130000;
#10;x=-216120000;
#10;x=-216110000;
#10;x=-216100000;
#10;x=-216090000;
#10;x=-216080000;
#10;x=-216070000;
#10;x=-216060000;
#10;x=-216050000;
#10;x=-216040000;
#10;x=-216030000;
#10;x=-216020000;
#10;x=-216010000;
#10;x=-216000000;
#10;x=-215990000;
#10;x=-215980000;
#10;x=-215970000;
#10;x=-215960000;
#10;x=-215950000;
#10;x=-215940000;
#10;x=-215930000;
#10;x=-215920000;
#10;x=-215910000;
#10;x=-215900000;
#10;x=-215890000;
#10;x=-215880000;
#10;x=-215870000;
#10;x=-215860000;
#10;x=-215850000;
#10;x=-215840000;
#10;x=-215830000;
#10;x=-215820000;
#10;x=-215810000;
#10;x=-215800000;
#10;x=-215790000;
#10;x=-215780000;
#10;x=-215770000;
#10;x=-215760000;
#10;x=-215750000;
#10;x=-215740000;
#10;x=-215730000;
#10;x=-215720000;
#10;x=-215710000;
#10;x=-215700000;
#10;x=-215690000;
#10;x=-215680000;
#10;x=-215670000;
#10;x=-215660000;
#10;x=-215650000;
#10;x=-215640000;
#10;x=-215630000;
#10;x=-215620000;
#10;x=-215610000;
#10;x=-215600000;
#10;x=-215590000;
#10;x=-215580000;
#10;x=-215570000;
#10;x=-215560000;
#10;x=-215550000;
#10;x=-215540000;
#10;x=-215530000;
#10;x=-215520000;
#10;x=-215510000;
#10;x=-215500000;
#10;x=-215490000;
#10;x=-215480000;
#10;x=-215470000;
#10;x=-215460000;
#10;x=-215450000;
#10;x=-215440000;
#10;x=-215430000;
#10;x=-215420000;
#10;x=-215410000;
#10;x=-215400000;
#10;x=-215390000;
#10;x=-215380000;
#10;x=-215370000;
#10;x=-215360000;
#10;x=-215350000;
#10;x=-215340000;
#10;x=-215330000;
#10;x=-215320000;
#10;x=-215310000;
#10;x=-215300000;
#10;x=-215290000;
#10;x=-215280000;
#10;x=-215270000;
#10;x=-215260000;
#10;x=-215250000;
#10;x=-215240000;
#10;x=-215230000;
#10;x=-215220000;
#10;x=-215210000;
#10;x=-215200000;
#10;x=-215190000;
#10;x=-215180000;
#10;x=-215170000;
#10;x=-215160000;
#10;x=-215150000;
#10;x=-215140000;
#10;x=-215130000;
#10;x=-215120000;
#10;x=-215110000;
#10;x=-215100000;
#10;x=-215090000;
#10;x=-215080000;
#10;x=-215070000;
#10;x=-215060000;
#10;x=-215050000;
#10;x=-215040000;
#10;x=-215030000;
#10;x=-215020000;
#10;x=-215010000;
#10;x=-215000000;
#10;x=-214990000;
#10;x=-214980000;
#10;x=-214970000;
#10;x=-214960000;
#10;x=-214950000;
#10;x=-214940000;
#10;x=-214930000;
#10;x=-214920000;
#10;x=-214910000;
#10;x=-214900000;
#10;x=-214890000;
#10;x=-214880000;
#10;x=-214870000;
#10;x=-214860000;
#10;x=-214850000;
#10;x=-214840000;
#10;x=-214830000;
#10;x=-214820000;
#10;x=-214810000;
#10;x=-214800000;
#10;x=-214790000;
#10;x=-214780000;
#10;x=-214770000;
#10;x=-214760000;
#10;x=-214750000;
#10;x=-214740000;
#10;x=-214730000;
#10;x=-214720000;
#10;x=-214710000;
#10;x=-214700000;
#10;x=-214690000;
#10;x=-214680000;
#10;x=-214670000;
#10;x=-214660000;
#10;x=-214650000;
#10;x=-214640000;
#10;x=-214630000;
#10;x=-214620000;
#10;x=-214610000;
#10;x=-214600000;
#10;x=-214590000;
#10;x=-214580000;
#10;x=-214570000;
#10;x=-214560000;
#10;x=-214550000;
#10;x=-214540000;
#10;x=-214530000;
#10;x=-214520000;
#10;x=-214510000;
#10;x=-214500000;
#10;x=-214490000;
#10;x=-214480000;
#10;x=-214470000;
#10;x=-214460000;
#10;x=-214450000;
#10;x=-214440000;
#10;x=-214430000;
#10;x=-214420000;
#10;x=-214410000;
#10;x=-214400000;
#10;x=-214390000;
#10;x=-214380000;
#10;x=-214370000;
#10;x=-214360000;
#10;x=-214350000;
#10;x=-214340000;
#10;x=-214330000;
#10;x=-214320000;
#10;x=-214310000;
#10;x=-214300000;
#10;x=-214290000;
#10;x=-214280000;
#10;x=-214270000;
#10;x=-214260000;
#10;x=-214250000;
#10;x=-214240000;
#10;x=-214230000;
#10;x=-214220000;
#10;x=-214210000;
#10;x=-214200000;
#10;x=-214190000;
#10;x=-214180000;
#10;x=-214170000;
#10;x=-214160000;
#10;x=-214150000;
#10;x=-214140000;
#10;x=-214130000;
#10;x=-214120000;
#10;x=-214110000;
#10;x=-214100000;
#10;x=-214090000;
#10;x=-214080000;
#10;x=-214070000;
#10;x=-214060000;
#10;x=-214050000;
#10;x=-214040000;
#10;x=-214030000;
#10;x=-214020000;
#10;x=-214010000;
#10;x=-214000000;
#10;x=-213990000;
#10;x=-213980000;
#10;x=-213970000;
#10;x=-213960000;
#10;x=-213950000;
#10;x=-213940000;
#10;x=-213930000;
#10;x=-213920000;
#10;x=-213910000;
#10;x=-213900000;
#10;x=-213890000;
#10;x=-213880000;
#10;x=-213870000;
#10;x=-213860000;
#10;x=-213850000;
#10;x=-213840000;
#10;x=-213830000;
#10;x=-213820000;
#10;x=-213810000;
#10;x=-213800000;
#10;x=-213790000;
#10;x=-213780000;
#10;x=-213770000;
#10;x=-213760000;
#10;x=-213750000;
#10;x=-213740000;
#10;x=-213730000;
#10;x=-213720000;
#10;x=-213710000;
#10;x=-213700000;
#10;x=-213690000;
#10;x=-213680000;
#10;x=-213670000;
#10;x=-213660000;
#10;x=-213650000;
#10;x=-213640000;
#10;x=-213630000;
#10;x=-213620000;
#10;x=-213610000;
#10;x=-213600000;
#10;x=-213590000;
#10;x=-213580000;
#10;x=-213570000;
#10;x=-213560000;
#10;x=-213550000;
#10;x=-213540000;
#10;x=-213530000;
#10;x=-213520000;
#10;x=-213510000;
#10;x=-213500000;
#10;x=-213490000;
#10;x=-213480000;
#10;x=-213470000;
#10;x=-213460000;
#10;x=-213450000;
#10;x=-213440000;
#10;x=-213430000;
#10;x=-213420000;
#10;x=-213410000;
#10;x=-213400000;
#10;x=-213390000;
#10;x=-213380000;
#10;x=-213370000;
#10;x=-213360000;
#10;x=-213350000;
#10;x=-213340000;
#10;x=-213330000;
#10;x=-213320000;
#10;x=-213310000;
#10;x=-213300000;
#10;x=-213290000;
#10;x=-213280000;
#10;x=-213270000;
#10;x=-213260000;
#10;x=-213250000;
#10;x=-213240000;
#10;x=-213230000;
#10;x=-213220000;
#10;x=-213210000;
#10;x=-213200000;
#10;x=-213190000;
#10;x=-213180000;
#10;x=-213170000;
#10;x=-213160000;
#10;x=-213150000;
#10;x=-213140000;
#10;x=-213130000;
#10;x=-213120000;
#10;x=-213110000;
#10;x=-213100000;
#10;x=-213090000;
#10;x=-213080000;
#10;x=-213070000;
#10;x=-213060000;
#10;x=-213050000;
#10;x=-213040000;
#10;x=-213030000;
#10;x=-213020000;
#10;x=-213010000;
#10;x=-213000000;
#10;x=-212990000;
#10;x=-212980000;
#10;x=-212970000;
#10;x=-212960000;
#10;x=-212950000;
#10;x=-212940000;
#10;x=-212930000;
#10;x=-212920000;
#10;x=-212910000;
#10;x=-212900000;
#10;x=-212890000;
#10;x=-212880000;
#10;x=-212870000;
#10;x=-212860000;
#10;x=-212850000;
#10;x=-212840000;
#10;x=-212830000;
#10;x=-212820000;
#10;x=-212810000;
#10;x=-212800000;
#10;x=-212790000;
#10;x=-212780000;
#10;x=-212770000;
#10;x=-212760000;
#10;x=-212750000;
#10;x=-212740000;
#10;x=-212730000;
#10;x=-212720000;
#10;x=-212710000;
#10;x=-212700000;
#10;x=-212690000;
#10;x=-212680000;
#10;x=-212670000;
#10;x=-212660000;
#10;x=-212650000;
#10;x=-212640000;
#10;x=-212630000;
#10;x=-212620000;
#10;x=-212610000;
#10;x=-212600000;
#10;x=-212590000;
#10;x=-212580000;
#10;x=-212570000;
#10;x=-212560000;
#10;x=-212550000;
#10;x=-212540000;
#10;x=-212530000;
#10;x=-212520000;
#10;x=-212510000;
#10;x=-212500000;
#10;x=-212490000;
#10;x=-212480000;
#10;x=-212470000;
#10;x=-212460000;
#10;x=-212450000;
#10;x=-212440000;
#10;x=-212430000;
#10;x=-212420000;
#10;x=-212410000;
#10;x=-212400000;
#10;x=-212390000;
#10;x=-212380000;
#10;x=-212370000;
#10;x=-212360000;
#10;x=-212350000;
#10;x=-212340000;
#10;x=-212330000;
#10;x=-212320000;
#10;x=-212310000;
#10;x=-212300000;
#10;x=-212290000;
#10;x=-212280000;
#10;x=-212270000;
#10;x=-212260000;
#10;x=-212250000;
#10;x=-212240000;
#10;x=-212230000;
#10;x=-212220000;
#10;x=-212210000;
#10;x=-212200000;
#10;x=-212190000;
#10;x=-212180000;
#10;x=-212170000;
#10;x=-212160000;
#10;x=-212150000;
#10;x=-212140000;
#10;x=-212130000;
#10;x=-212120000;
#10;x=-212110000;
#10;x=-212100000;
#10;x=-212090000;
#10;x=-212080000;
#10;x=-212070000;
#10;x=-212060000;
#10;x=-212050000;
#10;x=-212040000;
#10;x=-212030000;
#10;x=-212020000;
#10;x=-212010000;
#10;x=-212000000;
#10;x=-211990000;
#10;x=-211980000;
#10;x=-211970000;
#10;x=-211960000;
#10;x=-211950000;
#10;x=-211940000;
#10;x=-211930000;
#10;x=-211920000;
#10;x=-211910000;
#10;x=-211900000;
#10;x=-211890000;
#10;x=-211880000;
#10;x=-211870000;
#10;x=-211860000;
#10;x=-211850000;
#10;x=-211840000;
#10;x=-211830000;
#10;x=-211820000;
#10;x=-211810000;
#10;x=-211800000;
#10;x=-211790000;
#10;x=-211780000;
#10;x=-211770000;
#10;x=-211760000;
#10;x=-211750000;
#10;x=-211740000;
#10;x=-211730000;
#10;x=-211720000;
#10;x=-211710000;
#10;x=-211700000;
#10;x=-211690000;
#10;x=-211680000;
#10;x=-211670000;
#10;x=-211660000;
#10;x=-211650000;
#10;x=-211640000;
#10;x=-211630000;
#10;x=-211620000;
#10;x=-211610000;
#10;x=-211600000;
#10;x=-211590000;
#10;x=-211580000;
#10;x=-211570000;
#10;x=-211560000;
#10;x=-211550000;
#10;x=-211540000;
#10;x=-211530000;
#10;x=-211520000;
#10;x=-211510000;
#10;x=-211500000;
#10;x=-211490000;
#10;x=-211480000;
#10;x=-211470000;
#10;x=-211460000;
#10;x=-211450000;
#10;x=-211440000;
#10;x=-211430000;
#10;x=-211420000;
#10;x=-211410000;
#10;x=-211400000;
#10;x=-211390000;
#10;x=-211380000;
#10;x=-211370000;
#10;x=-211360000;
#10;x=-211350000;
#10;x=-211340000;
#10;x=-211330000;
#10;x=-211320000;
#10;x=-211310000;
#10;x=-211300000;
#10;x=-211290000;
#10;x=-211280000;
#10;x=-211270000;
#10;x=-211260000;
#10;x=-211250000;
#10;x=-211240000;
#10;x=-211230000;
#10;x=-211220000;
#10;x=-211210000;
#10;x=-211200000;
#10;x=-211190000;
#10;x=-211180000;
#10;x=-211170000;
#10;x=-211160000;
#10;x=-211150000;
#10;x=-211140000;
#10;x=-211130000;
#10;x=-211120000;
#10;x=-211110000;
#10;x=-211100000;
#10;x=-211090000;
#10;x=-211080000;
#10;x=-211070000;
#10;x=-211060000;
#10;x=-211050000;
#10;x=-211040000;
#10;x=-211030000;
#10;x=-211020000;
#10;x=-211010000;
#10;x=-211000000;
#10;x=-210990000;
#10;x=-210980000;
#10;x=-210970000;
#10;x=-210960000;
#10;x=-210950000;
#10;x=-210940000;
#10;x=-210930000;
#10;x=-210920000;
#10;x=-210910000;
#10;x=-210900000;
#10;x=-210890000;
#10;x=-210880000;
#10;x=-210870000;
#10;x=-210860000;
#10;x=-210850000;
#10;x=-210840000;
#10;x=-210830000;
#10;x=-210820000;
#10;x=-210810000;
#10;x=-210800000;
#10;x=-210790000;
#10;x=-210780000;
#10;x=-210770000;
#10;x=-210760000;
#10;x=-210750000;
#10;x=-210740000;
#10;x=-210730000;
#10;x=-210720000;
#10;x=-210710000;
#10;x=-210700000;
#10;x=-210690000;
#10;x=-210680000;
#10;x=-210670000;
#10;x=-210660000;
#10;x=-210650000;
#10;x=-210640000;
#10;x=-210630000;
#10;x=-210620000;
#10;x=-210610000;
#10;x=-210600000;
#10;x=-210590000;
#10;x=-210580000;
#10;x=-210570000;
#10;x=-210560000;
#10;x=-210550000;
#10;x=-210540000;
#10;x=-210530000;
#10;x=-210520000;
#10;x=-210510000;
#10;x=-210500000;
#10;x=-210490000;
#10;x=-210480000;
#10;x=-210470000;
#10;x=-210460000;
#10;x=-210450000;
#10;x=-210440000;
#10;x=-210430000;
#10;x=-210420000;
#10;x=-210410000;
#10;x=-210400000;
#10;x=-210390000;
#10;x=-210380000;
#10;x=-210370000;
#10;x=-210360000;
#10;x=-210350000;
#10;x=-210340000;
#10;x=-210330000;
#10;x=-210320000;
#10;x=-210310000;
#10;x=-210300000;
#10;x=-210290000;
#10;x=-210280000;
#10;x=-210270000;
#10;x=-210260000;
#10;x=-210250000;
#10;x=-210240000;
#10;x=-210230000;
#10;x=-210220000;
#10;x=-210210000;
#10;x=-210200000;
#10;x=-210190000;
#10;x=-210180000;
#10;x=-210170000;
#10;x=-210160000;
#10;x=-210150000;
#10;x=-210140000;
#10;x=-210130000;
#10;x=-210120000;
#10;x=-210110000;
#10;x=-210100000;
#10;x=-210090000;
#10;x=-210080000;
#10;x=-210070000;
#10;x=-210060000;
#10;x=-210050000;
#10;x=-210040000;
#10;x=-210030000;
#10;x=-210020000;
#10;x=-210010000;
#10;x=-210000000;
#10;x=-209990000;
#10;x=-209980000;
#10;x=-209970000;
#10;x=-209960000;
#10;x=-209950000;
#10;x=-209940000;
#10;x=-209930000;
#10;x=-209920000;
#10;x=-209910000;
#10;x=-209900000;
#10;x=-209890000;
#10;x=-209880000;
#10;x=-209870000;
#10;x=-209860000;
#10;x=-209850000;
#10;x=-209840000;
#10;x=-209830000;
#10;x=-209820000;
#10;x=-209810000;
#10;x=-209800000;
#10;x=-209790000;
#10;x=-209780000;
#10;x=-209770000;
#10;x=-209760000;
#10;x=-209750000;
#10;x=-209740000;
#10;x=-209730000;
#10;x=-209720000;
#10;x=-209710000;
#10;x=-209700000;
#10;x=-209690000;
#10;x=-209680000;
#10;x=-209670000;
#10;x=-209660000;
#10;x=-209650000;
#10;x=-209640000;
#10;x=-209630000;
#10;x=-209620000;
#10;x=-209610000;
#10;x=-209600000;
#10;x=-209590000;
#10;x=-209580000;
#10;x=-209570000;
#10;x=-209560000;
#10;x=-209550000;
#10;x=-209540000;
#10;x=-209530000;
#10;x=-209520000;
#10;x=-209510000;
#10;x=-209500000;
#10;x=-209490000;
#10;x=-209480000;
#10;x=-209470000;
#10;x=-209460000;
#10;x=-209450000;
#10;x=-209440000;
#10;x=-209430000;
#10;x=-209420000;
#10;x=-209410000;
#10;x=-209400000;
#10;x=-209390000;
#10;x=-209380000;
#10;x=-209370000;
#10;x=-209360000;
#10;x=-209350000;
#10;x=-209340000;
#10;x=-209330000;
#10;x=-209320000;
#10;x=-209310000;
#10;x=-209300000;
#10;x=-209290000;
#10;x=-209280000;
#10;x=-209270000;
#10;x=-209260000;
#10;x=-209250000;
#10;x=-209240000;
#10;x=-209230000;
#10;x=-209220000;
#10;x=-209210000;
#10;x=-209200000;
#10;x=-209190000;
#10;x=-209180000;
#10;x=-209170000;
#10;x=-209160000;
#10;x=-209150000;
#10;x=-209140000;
#10;x=-209130000;
#10;x=-209120000;
#10;x=-209110000;
#10;x=-209100000;
#10;x=-209090000;
#10;x=-209080000;
#10;x=-209070000;
#10;x=-209060000;
#10;x=-209050000;
#10;x=-209040000;
#10;x=-209030000;
#10;x=-209020000;
#10;x=-209010000;
#10;x=-209000000;
#10;x=-208990000;
#10;x=-208980000;
#10;x=-208970000;
#10;x=-208960000;
#10;x=-208950000;
#10;x=-208940000;
#10;x=-208930000;
#10;x=-208920000;
#10;x=-208910000;
#10;x=-208900000;
#10;x=-208890000;
#10;x=-208880000;
#10;x=-208870000;
#10;x=-208860000;
#10;x=-208850000;
#10;x=-208840000;
#10;x=-208830000;
#10;x=-208820000;
#10;x=-208810000;
#10;x=-208800000;
#10;x=-208790000;
#10;x=-208780000;
#10;x=-208770000;
#10;x=-208760000;
#10;x=-208750000;
#10;x=-208740000;
#10;x=-208730000;
#10;x=-208720000;
#10;x=-208710000;
#10;x=-208700000;
#10;x=-208690000;
#10;x=-208680000;
#10;x=-208670000;
#10;x=-208660000;
#10;x=-208650000;
#10;x=-208640000;
#10;x=-208630000;
#10;x=-208620000;
#10;x=-208610000;
#10;x=-208600000;
#10;x=-208590000;
#10;x=-208580000;
#10;x=-208570000;
#10;x=-208560000;
#10;x=-208550000;
#10;x=-208540000;
#10;x=-208530000;
#10;x=-208520000;
#10;x=-208510000;
#10;x=-208500000;
#10;x=-208490000;
#10;x=-208480000;
#10;x=-208470000;
#10;x=-208460000;
#10;x=-208450000;
#10;x=-208440000;
#10;x=-208430000;
#10;x=-208420000;
#10;x=-208410000;
#10;x=-208400000;
#10;x=-208390000;
#10;x=-208380000;
#10;x=-208370000;
#10;x=-208360000;
#10;x=-208350000;
#10;x=-208340000;
#10;x=-208330000;
#10;x=-208320000;
#10;x=-208310000;
#10;x=-208300000;
#10;x=-208290000;
#10;x=-208280000;
#10;x=-208270000;
#10;x=-208260000;
#10;x=-208250000;
#10;x=-208240000;
#10;x=-208230000;
#10;x=-208220000;
#10;x=-208210000;
#10;x=-208200000;
#10;x=-208190000;
#10;x=-208180000;
#10;x=-208170000;
#10;x=-208160000;
#10;x=-208150000;
#10;x=-208140000;
#10;x=-208130000;
#10;x=-208120000;
#10;x=-208110000;
#10;x=-208100000;
#10;x=-208090000;
#10;x=-208080000;
#10;x=-208070000;
#10;x=-208060000;
#10;x=-208050000;
#10;x=-208040000;
#10;x=-208030000;
#10;x=-208020000;
#10;x=-208010000;
#10;x=-208000000;
#10;x=-207990000;
#10;x=-207980000;
#10;x=-207970000;
#10;x=-207960000;
#10;x=-207950000;
#10;x=-207940000;
#10;x=-207930000;
#10;x=-207920000;
#10;x=-207910000;
#10;x=-207900000;
#10;x=-207890000;
#10;x=-207880000;
#10;x=-207870000;
#10;x=-207860000;
#10;x=-207850000;
#10;x=-207840000;
#10;x=-207830000;
#10;x=-207820000;
#10;x=-207810000;
#10;x=-207800000;
#10;x=-207790000;
#10;x=-207780000;
#10;x=-207770000;
#10;x=-207760000;
#10;x=-207750000;
#10;x=-207740000;
#10;x=-207730000;
#10;x=-207720000;
#10;x=-207710000;
#10;x=-207700000;
#10;x=-207690000;
#10;x=-207680000;
#10;x=-207670000;
#10;x=-207660000;
#10;x=-207650000;
#10;x=-207640000;
#10;x=-207630000;
#10;x=-207620000;
#10;x=-207610000;
#10;x=-207600000;
#10;x=-207590000;
#10;x=-207580000;
#10;x=-207570000;
#10;x=-207560000;
#10;x=-207550000;
#10;x=-207540000;
#10;x=-207530000;
#10;x=-207520000;
#10;x=-207510000;
#10;x=-207500000;
#10;x=-207490000;
#10;x=-207480000;
#10;x=-207470000;
#10;x=-207460000;
#10;x=-207450000;
#10;x=-207440000;
#10;x=-207430000;
#10;x=-207420000;
#10;x=-207410000;
#10;x=-207400000;
#10;x=-207390000;
#10;x=-207380000;
#10;x=-207370000;
#10;x=-207360000;
#10;x=-207350000;
#10;x=-207340000;
#10;x=-207330000;
#10;x=-207320000;
#10;x=-207310000;
#10;x=-207300000;
#10;x=-207290000;
#10;x=-207280000;
#10;x=-207270000;
#10;x=-207260000;
#10;x=-207250000;
#10;x=-207240000;
#10;x=-207230000;
#10;x=-207220000;
#10;x=-207210000;
#10;x=-207200000;
#10;x=-207190000;
#10;x=-207180000;
#10;x=-207170000;
#10;x=-207160000;
#10;x=-207150000;
#10;x=-207140000;
#10;x=-207130000;
#10;x=-207120000;
#10;x=-207110000;
#10;x=-207100000;
#10;x=-207090000;
#10;x=-207080000;
#10;x=-207070000;
#10;x=-207060000;
#10;x=-207050000;
#10;x=-207040000;
#10;x=-207030000;
#10;x=-207020000;
#10;x=-207010000;
#10;x=-207000000;
#10;x=-206990000;
#10;x=-206980000;
#10;x=-206970000;
#10;x=-206960000;
#10;x=-206950000;
#10;x=-206940000;
#10;x=-206930000;
#10;x=-206920000;
#10;x=-206910000;
#10;x=-206900000;
#10;x=-206890000;
#10;x=-206880000;
#10;x=-206870000;
#10;x=-206860000;
#10;x=-206850000;
#10;x=-206840000;
#10;x=-206830000;
#10;x=-206820000;
#10;x=-206810000;
#10;x=-206800000;
#10;x=-206790000;
#10;x=-206780000;
#10;x=-206770000;
#10;x=-206760000;
#10;x=-206750000;
#10;x=-206740000;
#10;x=-206730000;
#10;x=-206720000;
#10;x=-206710000;
#10;x=-206700000;
#10;x=-206690000;
#10;x=-206680000;
#10;x=-206670000;
#10;x=-206660000;
#10;x=-206650000;
#10;x=-206640000;
#10;x=-206630000;
#10;x=-206620000;
#10;x=-206610000;
#10;x=-206600000;
#10;x=-206590000;
#10;x=-206580000;
#10;x=-206570000;
#10;x=-206560000;
#10;x=-206550000;
#10;x=-206540000;
#10;x=-206530000;
#10;x=-206520000;
#10;x=-206510000;
#10;x=-206500000;
#10;x=-206490000;
#10;x=-206480000;
#10;x=-206470000;
#10;x=-206460000;
#10;x=-206450000;
#10;x=-206440000;
#10;x=-206430000;
#10;x=-206420000;
#10;x=-206410000;
#10;x=-206400000;
#10;x=-206390000;
#10;x=-206380000;
#10;x=-206370000;
#10;x=-206360000;
#10;x=-206350000;
#10;x=-206340000;
#10;x=-206330000;
#10;x=-206320000;
#10;x=-206310000;
#10;x=-206300000;
#10;x=-206290000;
#10;x=-206280000;
#10;x=-206270000;
#10;x=-206260000;
#10;x=-206250000;
#10;x=-206240000;
#10;x=-206230000;
#10;x=-206220000;
#10;x=-206210000;
#10;x=-206200000;
#10;x=-206190000;
#10;x=-206180000;
#10;x=-206170000;
#10;x=-206160000;
#10;x=-206150000;
#10;x=-206140000;
#10;x=-206130000;
#10;x=-206120000;
#10;x=-206110000;
#10;x=-206100000;
#10;x=-206090000;
#10;x=-206080000;
#10;x=-206070000;
#10;x=-206060000;
#10;x=-206050000;
#10;x=-206040000;
#10;x=-206030000;
#10;x=-206020000;
#10;x=-206010000;
#10;x=-206000000;
#10;x=-205990000;
#10;x=-205980000;
#10;x=-205970000;
#10;x=-205960000;
#10;x=-205950000;
#10;x=-205940000;
#10;x=-205930000;
#10;x=-205920000;
#10;x=-205910000;
#10;x=-205900000;
#10;x=-205890000;
#10;x=-205880000;
#10;x=-205870000;
#10;x=-205860000;
#10;x=-205850000;
#10;x=-205840000;
#10;x=-205830000;
#10;x=-205820000;
#10;x=-205810000;
#10;x=-205800000;
#10;x=-205790000;
#10;x=-205780000;
#10;x=-205770000;
#10;x=-205760000;
#10;x=-205750000;
#10;x=-205740000;
#10;x=-205730000;
#10;x=-205720000;
#10;x=-205710000;
#10;x=-205700000;
#10;x=-205690000;
#10;x=-205680000;
#10;x=-205670000;
#10;x=-205660000;
#10;x=-205650000;
#10;x=-205640000;
#10;x=-205630000;
#10;x=-205620000;
#10;x=-205610000;
#10;x=-205600000;
#10;x=-205590000;
#10;x=-205580000;
#10;x=-205570000;
#10;x=-205560000;
#10;x=-205550000;
#10;x=-205540000;
#10;x=-205530000;
#10;x=-205520000;
#10;x=-205510000;
#10;x=-205500000;
#10;x=-205490000;
#10;x=-205480000;
#10;x=-205470000;
#10;x=-205460000;
#10;x=-205450000;
#10;x=-205440000;
#10;x=-205430000;
#10;x=-205420000;
#10;x=-205410000;
#10;x=-205400000;
#10;x=-205390000;
#10;x=-205380000;
#10;x=-205370000;
#10;x=-205360000;
#10;x=-205350000;
#10;x=-205340000;
#10;x=-205330000;
#10;x=-205320000;
#10;x=-205310000;
#10;x=-205300000;
#10;x=-205290000;
#10;x=-205280000;
#10;x=-205270000;
#10;x=-205260000;
#10;x=-205250000;
#10;x=-205240000;
#10;x=-205230000;
#10;x=-205220000;
#10;x=-205210000;
#10;x=-205200000;
#10;x=-205190000;
#10;x=-205180000;
#10;x=-205170000;
#10;x=-205160000;
#10;x=-205150000;
#10;x=-205140000;
#10;x=-205130000;
#10;x=-205120000;
#10;x=-205110000;
#10;x=-205100000;
#10;x=-205090000;
#10;x=-205080000;
#10;x=-205070000;
#10;x=-205060000;
#10;x=-205050000;
#10;x=-205040000;
#10;x=-205030000;
#10;x=-205020000;
#10;x=-205010000;
#10;x=-205000000;
#10;x=-204990000;
#10;x=-204980000;
#10;x=-204970000;
#10;x=-204960000;
#10;x=-204950000;
#10;x=-204940000;
#10;x=-204930000;
#10;x=-204920000;
#10;x=-204910000;
#10;x=-204900000;
#10;x=-204890000;
#10;x=-204880000;
#10;x=-204870000;
#10;x=-204860000;
#10;x=-204850000;
#10;x=-204840000;
#10;x=-204830000;
#10;x=-204820000;
#10;x=-204810000;
#10;x=-204800000;
#10;x=-204790000;
#10;x=-204780000;
#10;x=-204770000;
#10;x=-204760000;
#10;x=-204750000;
#10;x=-204740000;
#10;x=-204730000;
#10;x=-204720000;
#10;x=-204710000;
#10;x=-204700000;
#10;x=-204690000;
#10;x=-204680000;
#10;x=-204670000;
#10;x=-204660000;
#10;x=-204650000;
#10;x=-204640000;
#10;x=-204630000;
#10;x=-204620000;
#10;x=-204610000;
#10;x=-204600000;
#10;x=-204590000;
#10;x=-204580000;
#10;x=-204570000;
#10;x=-204560000;
#10;x=-204550000;
#10;x=-204540000;
#10;x=-204530000;
#10;x=-204520000;
#10;x=-204510000;
#10;x=-204500000;
#10;x=-204490000;
#10;x=-204480000;
#10;x=-204470000;
#10;x=-204460000;
#10;x=-204450000;
#10;x=-204440000;
#10;x=-204430000;
#10;x=-204420000;
#10;x=-204410000;
#10;x=-204400000;
#10;x=-204390000;
#10;x=-204380000;
#10;x=-204370000;
#10;x=-204360000;
#10;x=-204350000;
#10;x=-204340000;
#10;x=-204330000;
#10;x=-204320000;
#10;x=-204310000;
#10;x=-204300000;
#10;x=-204290000;
#10;x=-204280000;
#10;x=-204270000;
#10;x=-204260000;
#10;x=-204250000;
#10;x=-204240000;
#10;x=-204230000;
#10;x=-204220000;
#10;x=-204210000;
#10;x=-204200000;
#10;x=-204190000;
#10;x=-204180000;
#10;x=-204170000;
#10;x=-204160000;
#10;x=-204150000;
#10;x=-204140000;
#10;x=-204130000;
#10;x=-204120000;
#10;x=-204110000;
#10;x=-204100000;
#10;x=-204090000;
#10;x=-204080000;
#10;x=-204070000;
#10;x=-204060000;
#10;x=-204050000;
#10;x=-204040000;
#10;x=-204030000;
#10;x=-204020000;
#10;x=-204010000;
#10;x=-204000000;
#10;x=-203990000;
#10;x=-203980000;
#10;x=-203970000;
#10;x=-203960000;
#10;x=-203950000;
#10;x=-203940000;
#10;x=-203930000;
#10;x=-203920000;
#10;x=-203910000;
#10;x=-203900000;
#10;x=-203890000;
#10;x=-203880000;
#10;x=-203870000;
#10;x=-203860000;
#10;x=-203850000;
#10;x=-203840000;
#10;x=-203830000;
#10;x=-203820000;
#10;x=-203810000;
#10;x=-203800000;
#10;x=-203790000;
#10;x=-203780000;
#10;x=-203770000;
#10;x=-203760000;
#10;x=-203750000;
#10;x=-203740000;
#10;x=-203730000;
#10;x=-203720000;
#10;x=-203710000;
#10;x=-203700000;
#10;x=-203690000;
#10;x=-203680000;
#10;x=-203670000;
#10;x=-203660000;
#10;x=-203650000;
#10;x=-203640000;
#10;x=-203630000;
#10;x=-203620000;
#10;x=-203610000;
#10;x=-203600000;
#10;x=-203590000;
#10;x=-203580000;
#10;x=-203570000;
#10;x=-203560000;
#10;x=-203550000;
#10;x=-203540000;
#10;x=-203530000;
#10;x=-203520000;
#10;x=-203510000;
#10;x=-203500000;
#10;x=-203490000;
#10;x=-203480000;
#10;x=-203470000;
#10;x=-203460000;
#10;x=-203450000;
#10;x=-203440000;
#10;x=-203430000;
#10;x=-203420000;
#10;x=-203410000;
#10;x=-203400000;
#10;x=-203390000;
#10;x=-203380000;
#10;x=-203370000;
#10;x=-203360000;
#10;x=-203350000;
#10;x=-203340000;
#10;x=-203330000;
#10;x=-203320000;
#10;x=-203310000;
#10;x=-203300000;
#10;x=-203290000;
#10;x=-203280000;
#10;x=-203270000;
#10;x=-203260000;
#10;x=-203250000;
#10;x=-203240000;
#10;x=-203230000;
#10;x=-203220000;
#10;x=-203210000;
#10;x=-203200000;
#10;x=-203190000;
#10;x=-203180000;
#10;x=-203170000;
#10;x=-203160000;
#10;x=-203150000;
#10;x=-203140000;
#10;x=-203130000;
#10;x=-203120000;
#10;x=-203110000;
#10;x=-203100000;
#10;x=-203090000;
#10;x=-203080000;
#10;x=-203070000;
#10;x=-203060000;
#10;x=-203050000;
#10;x=-203040000;
#10;x=-203030000;
#10;x=-203020000;
#10;x=-203010000;
#10;x=-203000000;
#10;x=-202990000;
#10;x=-202980000;
#10;x=-202970000;
#10;x=-202960000;
#10;x=-202950000;
#10;x=-202940000;
#10;x=-202930000;
#10;x=-202920000;
#10;x=-202910000;
#10;x=-202900000;
#10;x=-202890000;
#10;x=-202880000;
#10;x=-202870000;
#10;x=-202860000;
#10;x=-202850000;
#10;x=-202840000;
#10;x=-202830000;
#10;x=-202820000;
#10;x=-202810000;
#10;x=-202800000;
#10;x=-202790000;
#10;x=-202780000;
#10;x=-202770000;
#10;x=-202760000;
#10;x=-202750000;
#10;x=-202740000;
#10;x=-202730000;
#10;x=-202720000;
#10;x=-202710000;
#10;x=-202700000;
#10;x=-202690000;
#10;x=-202680000;
#10;x=-202670000;
#10;x=-202660000;
#10;x=-202650000;
#10;x=-202640000;
#10;x=-202630000;
#10;x=-202620000;
#10;x=-202610000;
#10;x=-202600000;
#10;x=-202590000;
#10;x=-202580000;
#10;x=-202570000;
#10;x=-202560000;
#10;x=-202550000;
#10;x=-202540000;
#10;x=-202530000;
#10;x=-202520000;
#10;x=-202510000;
#10;x=-202500000;
#10;x=-202490000;
#10;x=-202480000;
#10;x=-202470000;
#10;x=-202460000;
#10;x=-202450000;
#10;x=-202440000;
#10;x=-202430000;
#10;x=-202420000;
#10;x=-202410000;
#10;x=-202400000;
#10;x=-202390000;
#10;x=-202380000;
#10;x=-202370000;
#10;x=-202360000;
#10;x=-202350000;
#10;x=-202340000;
#10;x=-202330000;
#10;x=-202320000;
#10;x=-202310000;
#10;x=-202300000;
#10;x=-202290000;
#10;x=-202280000;
#10;x=-202270000;
#10;x=-202260000;
#10;x=-202250000;
#10;x=-202240000;
#10;x=-202230000;
#10;x=-202220000;
#10;x=-202210000;
#10;x=-202200000;
#10;x=-202190000;
#10;x=-202180000;
#10;x=-202170000;
#10;x=-202160000;
#10;x=-202150000;
#10;x=-202140000;
#10;x=-202130000;
#10;x=-202120000;
#10;x=-202110000;
#10;x=-202100000;
#10;x=-202090000;
#10;x=-202080000;
#10;x=-202070000;
#10;x=-202060000;
#10;x=-202050000;
#10;x=-202040000;
#10;x=-202030000;
#10;x=-202020000;
#10;x=-202010000;
#10;x=-202000000;
#10;x=-201990000;
#10;x=-201980000;
#10;x=-201970000;
#10;x=-201960000;
#10;x=-201950000;
#10;x=-201940000;
#10;x=-201930000;
#10;x=-201920000;
#10;x=-201910000;
#10;x=-201900000;
#10;x=-201890000;
#10;x=-201880000;
#10;x=-201870000;
#10;x=-201860000;
#10;x=-201850000;
#10;x=-201840000;
#10;x=-201830000;
#10;x=-201820000;
#10;x=-201810000;
#10;x=-201800000;
#10;x=-201790000;
#10;x=-201780000;
#10;x=-201770000;
#10;x=-201760000;
#10;x=-201750000;
#10;x=-201740000;
#10;x=-201730000;
#10;x=-201720000;
#10;x=-201710000;
#10;x=-201700000;
#10;x=-201690000;
#10;x=-201680000;
#10;x=-201670000;
#10;x=-201660000;
#10;x=-201650000;
#10;x=-201640000;
#10;x=-201630000;
#10;x=-201620000;
#10;x=-201610000;
#10;x=-201600000;
#10;x=-201590000;
#10;x=-201580000;
#10;x=-201570000;
#10;x=-201560000;
#10;x=-201550000;
#10;x=-201540000;
#10;x=-201530000;
#10;x=-201520000;
#10;x=-201510000;
#10;x=-201500000;
#10;x=-201490000;
#10;x=-201480000;
#10;x=-201470000;
#10;x=-201460000;
#10;x=-201450000;
#10;x=-201440000;
#10;x=-201430000;
#10;x=-201420000;
#10;x=-201410000;
#10;x=-201400000;
#10;x=-201390000;
#10;x=-201380000;
#10;x=-201370000;
#10;x=-201360000;
#10;x=-201350000;
#10;x=-201340000;
#10;x=-201330000;
#10;x=-201320000;
#10;x=-201310000;
#10;x=-201300000;
#10;x=-201290000;
#10;x=-201280000;
#10;x=-201270000;
#10;x=-201260000;
#10;x=-201250000;
#10;x=-201240000;
#10;x=-201230000;
#10;x=-201220000;
#10;x=-201210000;
#10;x=-201200000;
#10;x=-201190000;
#10;x=-201180000;
#10;x=-201170000;
#10;x=-201160000;
#10;x=-201150000;
#10;x=-201140000;
#10;x=-201130000;
#10;x=-201120000;
#10;x=-201110000;
#10;x=-201100000;
#10;x=-201090000;
#10;x=-201080000;
#10;x=-201070000;
#10;x=-201060000;
#10;x=-201050000;
#10;x=-201040000;
#10;x=-201030000;
#10;x=-201020000;
#10;x=-201010000;
#10;x=-201000000;
#10;x=-200990000;
#10;x=-200980000;
#10;x=-200970000;
#10;x=-200960000;
#10;x=-200950000;
#10;x=-200940000;
#10;x=-200930000;
#10;x=-200920000;
#10;x=-200910000;
#10;x=-200900000;
#10;x=-200890000;
#10;x=-200880000;
#10;x=-200870000;
#10;x=-200860000;
#10;x=-200850000;
#10;x=-200840000;
#10;x=-200830000;
#10;x=-200820000;
#10;x=-200810000;
#10;x=-200800000;
#10;x=-200790000;
#10;x=-200780000;
#10;x=-200770000;
#10;x=-200760000;
#10;x=-200750000;
#10;x=-200740000;
#10;x=-200730000;
#10;x=-200720000;
#10;x=-200710000;
#10;x=-200700000;
#10;x=-200690000;
#10;x=-200680000;
#10;x=-200670000;
#10;x=-200660000;
#10;x=-200650000;
#10;x=-200640000;
#10;x=-200630000;
#10;x=-200620000;
#10;x=-200610000;
#10;x=-200600000;
#10;x=-200590000;
#10;x=-200580000;
#10;x=-200570000;
#10;x=-200560000;
#10;x=-200550000;
#10;x=-200540000;
#10;x=-200530000;
#10;x=-200520000;
#10;x=-200510000;
#10;x=-200500000;
#10;x=-200490000;
#10;x=-200480000;
#10;x=-200470000;
#10;x=-200460000;
#10;x=-200450000;
#10;x=-200440000;
#10;x=-200430000;
#10;x=-200420000;
#10;x=-200410000;
#10;x=-200400000;
#10;x=-200390000;
#10;x=-200380000;
#10;x=-200370000;
#10;x=-200360000;
#10;x=-200350000;
#10;x=-200340000;
#10;x=-200330000;
#10;x=-200320000;
#10;x=-200310000;
#10;x=-200300000;
#10;x=-200290000;
#10;x=-200280000;
#10;x=-200270000;
#10;x=-200260000;
#10;x=-200250000;
#10;x=-200240000;
#10;x=-200230000;
#10;x=-200220000;
#10;x=-200210000;
#10;x=-200200000;
#10;x=-200190000;
#10;x=-200180000;
#10;x=-200170000;
#10;x=-200160000;
#10;x=-200150000;
#10;x=-200140000;
#10;x=-200130000;
#10;x=-200120000;
#10;x=-200110000;
#10;x=-200100000;
#10;x=-200090000;
#10;x=-200080000;
#10;x=-200070000;
#10;x=-200060000;
#10;x=-200050000;
#10;x=-200040000;
#10;x=-200030000;
#10;x=-200020000;
#10;x=-200010000;
#10;x=-200000000;
#10;x=-199990000;
#10;x=-199980000;
#10;x=-199970000;
#10;x=-199960000;
#10;x=-199950000;
#10;x=-199940000;
#10;x=-199930000;
#10;x=-199920000;
#10;x=-199910000;
#10;x=-199900000;
#10;x=-199890000;
#10;x=-199880000;
#10;x=-199870000;
#10;x=-199860000;
#10;x=-199850000;
#10;x=-199840000;
#10;x=-199830000;
#10;x=-199820000;
#10;x=-199810000;
#10;x=-199800000;
#10;x=-199790000;
#10;x=-199780000;
#10;x=-199770000;
#10;x=-199760000;
#10;x=-199750000;
#10;x=-199740000;
#10;x=-199730000;
#10;x=-199720000;
#10;x=-199710000;
#10;x=-199700000;
#10;x=-199690000;
#10;x=-199680000;
#10;x=-199670000;
#10;x=-199660000;
#10;x=-199650000;
#10;x=-199640000;
#10;x=-199630000;
#10;x=-199620000;
#10;x=-199610000;
#10;x=-199600000;
#10;x=-199590000;
#10;x=-199580000;
#10;x=-199570000;
#10;x=-199560000;
#10;x=-199550000;
#10;x=-199540000;
#10;x=-199530000;
#10;x=-199520000;
#10;x=-199510000;
#10;x=-199500000;
#10;x=-199490000;
#10;x=-199480000;
#10;x=-199470000;
#10;x=-199460000;
#10;x=-199450000;
#10;x=-199440000;
#10;x=-199430000;
#10;x=-199420000;
#10;x=-199410000;
#10;x=-199400000;
#10;x=-199390000;
#10;x=-199380000;
#10;x=-199370000;
#10;x=-199360000;
#10;x=-199350000;
#10;x=-199340000;
#10;x=-199330000;
#10;x=-199320000;
#10;x=-199310000;
#10;x=-199300000;
#10;x=-199290000;
#10;x=-199280000;
#10;x=-199270000;
#10;x=-199260000;
#10;x=-199250000;
#10;x=-199240000;
#10;x=-199230000;
#10;x=-199220000;
#10;x=-199210000;
#10;x=-199200000;
#10;x=-199190000;
#10;x=-199180000;
#10;x=-199170000;
#10;x=-199160000;
#10;x=-199150000;
#10;x=-199140000;
#10;x=-199130000;
#10;x=-199120000;
#10;x=-199110000;
#10;x=-199100000;
#10;x=-199090000;
#10;x=-199080000;
#10;x=-199070000;
#10;x=-199060000;
#10;x=-199050000;
#10;x=-199040000;
#10;x=-199030000;
#10;x=-199020000;
#10;x=-199010000;
#10;x=-199000000;
#10;x=-198990000;
#10;x=-198980000;
#10;x=-198970000;
#10;x=-198960000;
#10;x=-198950000;
#10;x=-198940000;
#10;x=-198930000;
#10;x=-198920000;
#10;x=-198910000;
#10;x=-198900000;
#10;x=-198890000;
#10;x=-198880000;
#10;x=-198870000;
#10;x=-198860000;
#10;x=-198850000;
#10;x=-198840000;
#10;x=-198830000;
#10;x=-198820000;
#10;x=-198810000;
#10;x=-198800000;
#10;x=-198790000;
#10;x=-198780000;
#10;x=-198770000;
#10;x=-198760000;
#10;x=-198750000;
#10;x=-198740000;
#10;x=-198730000;
#10;x=-198720000;
#10;x=-198710000;
#10;x=-198700000;
#10;x=-198690000;
#10;x=-198680000;
#10;x=-198670000;
#10;x=-198660000;
#10;x=-198650000;
#10;x=-198640000;
#10;x=-198630000;
#10;x=-198620000;
#10;x=-198610000;
#10;x=-198600000;
#10;x=-198590000;
#10;x=-198580000;
#10;x=-198570000;
#10;x=-198560000;
#10;x=-198550000;
#10;x=-198540000;
#10;x=-198530000;
#10;x=-198520000;
#10;x=-198510000;
#10;x=-198500000;
#10;x=-198490000;
#10;x=-198480000;
#10;x=-198470000;
#10;x=-198460000;
#10;x=-198450000;
#10;x=-198440000;
#10;x=-198430000;
#10;x=-198420000;
#10;x=-198410000;
#10;x=-198400000;
#10;x=-198390000;
#10;x=-198380000;
#10;x=-198370000;
#10;x=-198360000;
#10;x=-198350000;
#10;x=-198340000;
#10;x=-198330000;
#10;x=-198320000;
#10;x=-198310000;
#10;x=-198300000;
#10;x=-198290000;
#10;x=-198280000;
#10;x=-198270000;
#10;x=-198260000;
#10;x=-198250000;
#10;x=-198240000;
#10;x=-198230000;
#10;x=-198220000;
#10;x=-198210000;
#10;x=-198200000;
#10;x=-198190000;
#10;x=-198180000;
#10;x=-198170000;
#10;x=-198160000;
#10;x=-198150000;
#10;x=-198140000;
#10;x=-198130000;
#10;x=-198120000;
#10;x=-198110000;
#10;x=-198100000;
#10;x=-198090000;
#10;x=-198080000;
#10;x=-198070000;
#10;x=-198060000;
#10;x=-198050000;
#10;x=-198040000;
#10;x=-198030000;
#10;x=-198020000;
#10;x=-198010000;
#10;x=-198000000;
#10;x=-197990000;
#10;x=-197980000;
#10;x=-197970000;
#10;x=-197960000;
#10;x=-197950000;
#10;x=-197940000;
#10;x=-197930000;
#10;x=-197920000;
#10;x=-197910000;
#10;x=-197900000;
#10;x=-197890000;
#10;x=-197880000;
#10;x=-197870000;
#10;x=-197860000;
#10;x=-197850000;
#10;x=-197840000;
#10;x=-197830000;
#10;x=-197820000;
#10;x=-197810000;
#10;x=-197800000;
#10;x=-197790000;
#10;x=-197780000;
#10;x=-197770000;
#10;x=-197760000;
#10;x=-197750000;
#10;x=-197740000;
#10;x=-197730000;
#10;x=-197720000;
#10;x=-197710000;
#10;x=-197700000;
#10;x=-197690000;
#10;x=-197680000;
#10;x=-197670000;
#10;x=-197660000;
#10;x=-197650000;
#10;x=-197640000;
#10;x=-197630000;
#10;x=-197620000;
#10;x=-197610000;
#10;x=-197600000;
#10;x=-197590000;
#10;x=-197580000;
#10;x=-197570000;
#10;x=-197560000;
#10;x=-197550000;
#10;x=-197540000;
#10;x=-197530000;
#10;x=-197520000;
#10;x=-197510000;
#10;x=-197500000;
#10;x=-197490000;
#10;x=-197480000;
#10;x=-197470000;
#10;x=-197460000;
#10;x=-197450000;
#10;x=-197440000;
#10;x=-197430000;
#10;x=-197420000;
#10;x=-197410000;
#10;x=-197400000;
#10;x=-197390000;
#10;x=-197380000;
#10;x=-197370000;
#10;x=-197360000;
#10;x=-197350000;
#10;x=-197340000;
#10;x=-197330000;
#10;x=-197320000;
#10;x=-197310000;
#10;x=-197300000;
#10;x=-197290000;
#10;x=-197280000;
#10;x=-197270000;
#10;x=-197260000;
#10;x=-197250000;
#10;x=-197240000;
#10;x=-197230000;
#10;x=-197220000;
#10;x=-197210000;
#10;x=-197200000;
#10;x=-197190000;
#10;x=-197180000;
#10;x=-197170000;
#10;x=-197160000;
#10;x=-197150000;
#10;x=-197140000;
#10;x=-197130000;
#10;x=-197120000;
#10;x=-197110000;
#10;x=-197100000;
#10;x=-197090000;
#10;x=-197080000;
#10;x=-197070000;
#10;x=-197060000;
#10;x=-197050000;
#10;x=-197040000;
#10;x=-197030000;
#10;x=-197020000;
#10;x=-197010000;
#10;x=-197000000;
#10;x=-196990000;
#10;x=-196980000;
#10;x=-196970000;
#10;x=-196960000;
#10;x=-196950000;
#10;x=-196940000;
#10;x=-196930000;
#10;x=-196920000;
#10;x=-196910000;
#10;x=-196900000;
#10;x=-196890000;
#10;x=-196880000;
#10;x=-196870000;
#10;x=-196860000;
#10;x=-196850000;
#10;x=-196840000;
#10;x=-196830000;
#10;x=-196820000;
#10;x=-196810000;
#10;x=-196800000;
#10;x=-196790000;
#10;x=-196780000;
#10;x=-196770000;
#10;x=-196760000;
#10;x=-196750000;
#10;x=-196740000;
#10;x=-196730000;
#10;x=-196720000;
#10;x=-196710000;
#10;x=-196700000;
#10;x=-196690000;
#10;x=-196680000;
#10;x=-196670000;
#10;x=-196660000;
#10;x=-196650000;
#10;x=-196640000;
#10;x=-196630000;
#10;x=-196620000;
#10;x=-196610000;
#10;x=-196600000;
#10;x=-196590000;
#10;x=-196580000;
#10;x=-196570000;
#10;x=-196560000;
#10;x=-196550000;
#10;x=-196540000;
#10;x=-196530000;
#10;x=-196520000;
#10;x=-196510000;
#10;x=-196500000;
#10;x=-196490000;
#10;x=-196480000;
#10;x=-196470000;
#10;x=-196460000;
#10;x=-196450000;
#10;x=-196440000;
#10;x=-196430000;
#10;x=-196420000;
#10;x=-196410000;
#10;x=-196400000;
#10;x=-196390000;
#10;x=-196380000;
#10;x=-196370000;
#10;x=-196360000;
#10;x=-196350000;
#10;x=-196340000;
#10;x=-196330000;
#10;x=-196320000;
#10;x=-196310000;
#10;x=-196300000;
#10;x=-196290000;
#10;x=-196280000;
#10;x=-196270000;
#10;x=-196260000;
#10;x=-196250000;
#10;x=-196240000;
#10;x=-196230000;
#10;x=-196220000;
#10;x=-196210000;
#10;x=-196200000;
#10;x=-196190000;
#10;x=-196180000;
#10;x=-196170000;
#10;x=-196160000;
#10;x=-196150000;
#10;x=-196140000;
#10;x=-196130000;
#10;x=-196120000;
#10;x=-196110000;
#10;x=-196100000;
#10;x=-196090000;
#10;x=-196080000;
#10;x=-196070000;
#10;x=-196060000;
#10;x=-196050000;
#10;x=-196040000;
#10;x=-196030000;
#10;x=-196020000;
#10;x=-196010000;
#10;x=-196000000;
#10;x=-195990000;
#10;x=-195980000;
#10;x=-195970000;
#10;x=-195960000;
#10;x=-195950000;
#10;x=-195940000;
#10;x=-195930000;
#10;x=-195920000;
#10;x=-195910000;
#10;x=-195900000;
#10;x=-195890000;
#10;x=-195880000;
#10;x=-195870000;
#10;x=-195860000;
#10;x=-195850000;
#10;x=-195840000;
#10;x=-195830000;
#10;x=-195820000;
#10;x=-195810000;
#10;x=-195800000;
#10;x=-195790000;
#10;x=-195780000;
#10;x=-195770000;
#10;x=-195760000;
#10;x=-195750000;
#10;x=-195740000;
#10;x=-195730000;
#10;x=-195720000;
#10;x=-195710000;
#10;x=-195700000;
#10;x=-195690000;
#10;x=-195680000;
#10;x=-195670000;
#10;x=-195660000;
#10;x=-195650000;
#10;x=-195640000;
#10;x=-195630000;
#10;x=-195620000;
#10;x=-195610000;
#10;x=-195600000;
#10;x=-195590000;
#10;x=-195580000;
#10;x=-195570000;
#10;x=-195560000;
#10;x=-195550000;
#10;x=-195540000;
#10;x=-195530000;
#10;x=-195520000;
#10;x=-195510000;
#10;x=-195500000;
#10;x=-195490000;
#10;x=-195480000;
#10;x=-195470000;
#10;x=-195460000;
#10;x=-195450000;
#10;x=-195440000;
#10;x=-195430000;
#10;x=-195420000;
#10;x=-195410000;
#10;x=-195400000;
#10;x=-195390000;
#10;x=-195380000;
#10;x=-195370000;
#10;x=-195360000;
#10;x=-195350000;
#10;x=-195340000;
#10;x=-195330000;
#10;x=-195320000;
#10;x=-195310000;
#10;x=-195300000;
#10;x=-195290000;
#10;x=-195280000;
#10;x=-195270000;
#10;x=-195260000;
#10;x=-195250000;
#10;x=-195240000;
#10;x=-195230000;
#10;x=-195220000;
#10;x=-195210000;
#10;x=-195200000;
#10;x=-195190000;
#10;x=-195180000;
#10;x=-195170000;
#10;x=-195160000;
#10;x=-195150000;
#10;x=-195140000;
#10;x=-195130000;
#10;x=-195120000;
#10;x=-195110000;
#10;x=-195100000;
#10;x=-195090000;
#10;x=-195080000;
#10;x=-195070000;
#10;x=-195060000;
#10;x=-195050000;
#10;x=-195040000;
#10;x=-195030000;
#10;x=-195020000;
#10;x=-195010000;
#10;x=-195000000;
#10;x=-194990000;
#10;x=-194980000;
#10;x=-194970000;
#10;x=-194960000;
#10;x=-194950000;
#10;x=-194940000;
#10;x=-194930000;
#10;x=-194920000;
#10;x=-194910000;
#10;x=-194900000;
#10;x=-194890000;
#10;x=-194880000;
#10;x=-194870000;
#10;x=-194860000;
#10;x=-194850000;
#10;x=-194840000;
#10;x=-194830000;
#10;x=-194820000;
#10;x=-194810000;
#10;x=-194800000;
#10;x=-194790000;
#10;x=-194780000;
#10;x=-194770000;
#10;x=-194760000;
#10;x=-194750000;
#10;x=-194740000;
#10;x=-194730000;
#10;x=-194720000;
#10;x=-194710000;
#10;x=-194700000;
#10;x=-194690000;
#10;x=-194680000;
#10;x=-194670000;
#10;x=-194660000;
#10;x=-194650000;
#10;x=-194640000;
#10;x=-194630000;
#10;x=-194620000;
#10;x=-194610000;
#10;x=-194600000;
#10;x=-194590000;
#10;x=-194580000;
#10;x=-194570000;
#10;x=-194560000;
#10;x=-194550000;
#10;x=-194540000;
#10;x=-194530000;
#10;x=-194520000;
#10;x=-194510000;
#10;x=-194500000;
#10;x=-194490000;
#10;x=-194480000;
#10;x=-194470000;
#10;x=-194460000;
#10;x=-194450000;
#10;x=-194440000;
#10;x=-194430000;
#10;x=-194420000;
#10;x=-194410000;
#10;x=-194400000;
#10;x=-194390000;
#10;x=-194380000;
#10;x=-194370000;
#10;x=-194360000;
#10;x=-194350000;
#10;x=-194340000;
#10;x=-194330000;
#10;x=-194320000;
#10;x=-194310000;
#10;x=-194300000;
#10;x=-194290000;
#10;x=-194280000;
#10;x=-194270000;
#10;x=-194260000;
#10;x=-194250000;
#10;x=-194240000;
#10;x=-194230000;
#10;x=-194220000;
#10;x=-194210000;
#10;x=-194200000;
#10;x=-194190000;
#10;x=-194180000;
#10;x=-194170000;
#10;x=-194160000;
#10;x=-194150000;
#10;x=-194140000;
#10;x=-194130000;
#10;x=-194120000;
#10;x=-194110000;
#10;x=-194100000;
#10;x=-194090000;
#10;x=-194080000;
#10;x=-194070000;
#10;x=-194060000;
#10;x=-194050000;
#10;x=-194040000;
#10;x=-194030000;
#10;x=-194020000;
#10;x=-194010000;
#10;x=-194000000;
#10;x=-193990000;
#10;x=-193980000;
#10;x=-193970000;
#10;x=-193960000;
#10;x=-193950000;
#10;x=-193940000;
#10;x=-193930000;
#10;x=-193920000;
#10;x=-193910000;
#10;x=-193900000;
#10;x=-193890000;
#10;x=-193880000;
#10;x=-193870000;
#10;x=-193860000;
#10;x=-193850000;
#10;x=-193840000;
#10;x=-193830000;
#10;x=-193820000;
#10;x=-193810000;
#10;x=-193800000;
#10;x=-193790000;
#10;x=-193780000;
#10;x=-193770000;
#10;x=-193760000;
#10;x=-193750000;
#10;x=-193740000;
#10;x=-193730000;
#10;x=-193720000;
#10;x=-193710000;
#10;x=-193700000;
#10;x=-193690000;
#10;x=-193680000;
#10;x=-193670000;
#10;x=-193660000;
#10;x=-193650000;
#10;x=-193640000;
#10;x=-193630000;
#10;x=-193620000;
#10;x=-193610000;
#10;x=-193600000;
#10;x=-193590000;
#10;x=-193580000;
#10;x=-193570000;
#10;x=-193560000;
#10;x=-193550000;
#10;x=-193540000;
#10;x=-193530000;
#10;x=-193520000;
#10;x=-193510000;
#10;x=-193500000;
#10;x=-193490000;
#10;x=-193480000;
#10;x=-193470000;
#10;x=-193460000;
#10;x=-193450000;
#10;x=-193440000;
#10;x=-193430000;
#10;x=-193420000;
#10;x=-193410000;
#10;x=-193400000;
#10;x=-193390000;
#10;x=-193380000;
#10;x=-193370000;
#10;x=-193360000;
#10;x=-193350000;
#10;x=-193340000;
#10;x=-193330000;
#10;x=-193320000;
#10;x=-193310000;
#10;x=-193300000;
#10;x=-193290000;
#10;x=-193280000;
#10;x=-193270000;
#10;x=-193260000;
#10;x=-193250000;
#10;x=-193240000;
#10;x=-193230000;
#10;x=-193220000;
#10;x=-193210000;
#10;x=-193200000;
#10;x=-193190000;
#10;x=-193180000;
#10;x=-193170000;
#10;x=-193160000;
#10;x=-193150000;
#10;x=-193140000;
#10;x=-193130000;
#10;x=-193120000;
#10;x=-193110000;
#10;x=-193100000;
#10;x=-193090000;
#10;x=-193080000;
#10;x=-193070000;
#10;x=-193060000;
#10;x=-193050000;
#10;x=-193040000;
#10;x=-193030000;
#10;x=-193020000;
#10;x=-193010000;
#10;x=-193000000;
#10;x=-192990000;
#10;x=-192980000;
#10;x=-192970000;
#10;x=-192960000;
#10;x=-192950000;
#10;x=-192940000;
#10;x=-192930000;
#10;x=-192920000;
#10;x=-192910000;
#10;x=-192900000;
#10;x=-192890000;
#10;x=-192880000;
#10;x=-192870000;
#10;x=-192860000;
#10;x=-192850000;
#10;x=-192840000;
#10;x=-192830000;
#10;x=-192820000;
#10;x=-192810000;
#10;x=-192800000;
#10;x=-192790000;
#10;x=-192780000;
#10;x=-192770000;
#10;x=-192760000;
#10;x=-192750000;
#10;x=-192740000;
#10;x=-192730000;
#10;x=-192720000;
#10;x=-192710000;
#10;x=-192700000;
#10;x=-192690000;
#10;x=-192680000;
#10;x=-192670000;
#10;x=-192660000;
#10;x=-192650000;
#10;x=-192640000;
#10;x=-192630000;
#10;x=-192620000;
#10;x=-192610000;
#10;x=-192600000;
#10;x=-192590000;
#10;x=-192580000;
#10;x=-192570000;
#10;x=-192560000;
#10;x=-192550000;
#10;x=-192540000;
#10;x=-192530000;
#10;x=-192520000;
#10;x=-192510000;
#10;x=-192500000;
#10;x=-192490000;
#10;x=-192480000;
#10;x=-192470000;
#10;x=-192460000;
#10;x=-192450000;
#10;x=-192440000;
#10;x=-192430000;
#10;x=-192420000;
#10;x=-192410000;
#10;x=-192400000;
#10;x=-192390000;
#10;x=-192380000;
#10;x=-192370000;
#10;x=-192360000;
#10;x=-192350000;
#10;x=-192340000;
#10;x=-192330000;
#10;x=-192320000;
#10;x=-192310000;
#10;x=-192300000;
#10;x=-192290000;
#10;x=-192280000;
#10;x=-192270000;
#10;x=-192260000;
#10;x=-192250000;
#10;x=-192240000;
#10;x=-192230000;
#10;x=-192220000;
#10;x=-192210000;
#10;x=-192200000;
#10;x=-192190000;
#10;x=-192180000;
#10;x=-192170000;
#10;x=-192160000;
#10;x=-192150000;
#10;x=-192140000;
#10;x=-192130000;
#10;x=-192120000;
#10;x=-192110000;
#10;x=-192100000;
#10;x=-192090000;
#10;x=-192080000;
#10;x=-192070000;
#10;x=-192060000;
#10;x=-192050000;
#10;x=-192040000;
#10;x=-192030000;
#10;x=-192020000;
#10;x=-192010000;
#10;x=-192000000;
#10;x=-191990000;
#10;x=-191980000;
#10;x=-191970000;
#10;x=-191960000;
#10;x=-191950000;
#10;x=-191940000;
#10;x=-191930000;
#10;x=-191920000;
#10;x=-191910000;
#10;x=-191900000;
#10;x=-191890000;
#10;x=-191880000;
#10;x=-191870000;
#10;x=-191860000;
#10;x=-191850000;
#10;x=-191840000;
#10;x=-191830000;
#10;x=-191820000;
#10;x=-191810000;
#10;x=-191800000;
#10;x=-191790000;
#10;x=-191780000;
#10;x=-191770000;
#10;x=-191760000;
#10;x=-191750000;
#10;x=-191740000;
#10;x=-191730000;
#10;x=-191720000;
#10;x=-191710000;
#10;x=-191700000;
#10;x=-191690000;
#10;x=-191680000;
#10;x=-191670000;
#10;x=-191660000;
#10;x=-191650000;
#10;x=-191640000;
#10;x=-191630000;
#10;x=-191620000;
#10;x=-191610000;
#10;x=-191600000;
#10;x=-191590000;
#10;x=-191580000;
#10;x=-191570000;
#10;x=-191560000;
#10;x=-191550000;
#10;x=-191540000;
#10;x=-191530000;
#10;x=-191520000;
#10;x=-191510000;
#10;x=-191500000;
#10;x=-191490000;
#10;x=-191480000;
#10;x=-191470000;
#10;x=-191460000;
#10;x=-191450000;
#10;x=-191440000;
#10;x=-191430000;
#10;x=-191420000;
#10;x=-191410000;
#10;x=-191400000;
#10;x=-191390000;
#10;x=-191380000;
#10;x=-191370000;
#10;x=-191360000;
#10;x=-191350000;
#10;x=-191340000;
#10;x=-191330000;
#10;x=-191320000;
#10;x=-191310000;
#10;x=-191300000;
#10;x=-191290000;
#10;x=-191280000;
#10;x=-191270000;
#10;x=-191260000;
#10;x=-191250000;
#10;x=-191240000;
#10;x=-191230000;
#10;x=-191220000;
#10;x=-191210000;
#10;x=-191200000;
#10;x=-191190000;
#10;x=-191180000;
#10;x=-191170000;
#10;x=-191160000;
#10;x=-191150000;
#10;x=-191140000;
#10;x=-191130000;
#10;x=-191120000;
#10;x=-191110000;
#10;x=-191100000;
#10;x=-191090000;
#10;x=-191080000;
#10;x=-191070000;
#10;x=-191060000;
#10;x=-191050000;
#10;x=-191040000;
#10;x=-191030000;
#10;x=-191020000;
#10;x=-191010000;
#10;x=-191000000;
#10;x=-190990000;
#10;x=-190980000;
#10;x=-190970000;
#10;x=-190960000;
#10;x=-190950000;
#10;x=-190940000;
#10;x=-190930000;
#10;x=-190920000;
#10;x=-190910000;
#10;x=-190900000;
#10;x=-190890000;
#10;x=-190880000;
#10;x=-190870000;
#10;x=-190860000;
#10;x=-190850000;
#10;x=-190840000;
#10;x=-190830000;
#10;x=-190820000;
#10;x=-190810000;
#10;x=-190800000;
#10;x=-190790000;
#10;x=-190780000;
#10;x=-190770000;
#10;x=-190760000;
#10;x=-190750000;
#10;x=-190740000;
#10;x=-190730000;
#10;x=-190720000;
#10;x=-190710000;
#10;x=-190700000;
#10;x=-190690000;
#10;x=-190680000;
#10;x=-190670000;
#10;x=-190660000;
#10;x=-190650000;
#10;x=-190640000;
#10;x=-190630000;
#10;x=-190620000;
#10;x=-190610000;
#10;x=-190600000;
#10;x=-190590000;
#10;x=-190580000;
#10;x=-190570000;
#10;x=-190560000;
#10;x=-190550000;
#10;x=-190540000;
#10;x=-190530000;
#10;x=-190520000;
#10;x=-190510000;
#10;x=-190500000;
#10;x=-190490000;
#10;x=-190480000;
#10;x=-190470000;
#10;x=-190460000;
#10;x=-190450000;
#10;x=-190440000;
#10;x=-190430000;
#10;x=-190420000;
#10;x=-190410000;
#10;x=-190400000;
#10;x=-190390000;
#10;x=-190380000;
#10;x=-190370000;
#10;x=-190360000;
#10;x=-190350000;
#10;x=-190340000;
#10;x=-190330000;
#10;x=-190320000;
#10;x=-190310000;
#10;x=-190300000;
#10;x=-190290000;
#10;x=-190280000;
#10;x=-190270000;
#10;x=-190260000;
#10;x=-190250000;
#10;x=-190240000;
#10;x=-190230000;
#10;x=-190220000;
#10;x=-190210000;
#10;x=-190200000;
#10;x=-190190000;
#10;x=-190180000;
#10;x=-190170000;
#10;x=-190160000;
#10;x=-190150000;
#10;x=-190140000;
#10;x=-190130000;
#10;x=-190120000;
#10;x=-190110000;
#10;x=-190100000;
#10;x=-190090000;
#10;x=-190080000;
#10;x=-190070000;
#10;x=-190060000;
#10;x=-190050000;
#10;x=-190040000;
#10;x=-190030000;
#10;x=-190020000;
#10;x=-190010000;
#10;x=-190000000;
#10;x=-189990000;
#10;x=-189980000;
#10;x=-189970000;
#10;x=-189960000;
#10;x=-189950000;
#10;x=-189940000;
#10;x=-189930000;
#10;x=-189920000;
#10;x=-189910000;
#10;x=-189900000;
#10;x=-189890000;
#10;x=-189880000;
#10;x=-189870000;
#10;x=-189860000;
#10;x=-189850000;
#10;x=-189840000;
#10;x=-189830000;
#10;x=-189820000;
#10;x=-189810000;
#10;x=-189800000;
#10;x=-189790000;
#10;x=-189780000;
#10;x=-189770000;
#10;x=-189760000;
#10;x=-189750000;
#10;x=-189740000;
#10;x=-189730000;
#10;x=-189720000;
#10;x=-189710000;
#10;x=-189700000;
#10;x=-189690000;
#10;x=-189680000;
#10;x=-189670000;
#10;x=-189660000;
#10;x=-189650000;
#10;x=-189640000;
#10;x=-189630000;
#10;x=-189620000;
#10;x=-189610000;
#10;x=-189600000;
#10;x=-189590000;
#10;x=-189580000;
#10;x=-189570000;
#10;x=-189560000;
#10;x=-189550000;
#10;x=-189540000;
#10;x=-189530000;
#10;x=-189520000;
#10;x=-189510000;
#10;x=-189500000;
#10;x=-189490000;
#10;x=-189480000;
#10;x=-189470000;
#10;x=-189460000;
#10;x=-189450000;
#10;x=-189440000;
#10;x=-189430000;
#10;x=-189420000;
#10;x=-189410000;
#10;x=-189400000;
#10;x=-189390000;
#10;x=-189380000;
#10;x=-189370000;
#10;x=-189360000;
#10;x=-189350000;
#10;x=-189340000;
#10;x=-189330000;
#10;x=-189320000;
#10;x=-189310000;
#10;x=-189300000;
#10;x=-189290000;
#10;x=-189280000;
#10;x=-189270000;
#10;x=-189260000;
#10;x=-189250000;
#10;x=-189240000;
#10;x=-189230000;
#10;x=-189220000;
#10;x=-189210000;
#10;x=-189200000;
#10;x=-189190000;
#10;x=-189180000;
#10;x=-189170000;
#10;x=-189160000;
#10;x=-189150000;
#10;x=-189140000;
#10;x=-189130000;
#10;x=-189120000;
#10;x=-189110000;
#10;x=-189100000;
#10;x=-189090000;
#10;x=-189080000;
#10;x=-189070000;
#10;x=-189060000;
#10;x=-189050000;
#10;x=-189040000;
#10;x=-189030000;
#10;x=-189020000;
#10;x=-189010000;
#10;x=-189000000;
#10;x=-188990000;
#10;x=-188980000;
#10;x=-188970000;
#10;x=-188960000;
#10;x=-188950000;
#10;x=-188940000;
#10;x=-188930000;
#10;x=-188920000;
#10;x=-188910000;
#10;x=-188900000;
#10;x=-188890000;
#10;x=-188880000;
#10;x=-188870000;
#10;x=-188860000;
#10;x=-188850000;
#10;x=-188840000;
#10;x=-188830000;
#10;x=-188820000;
#10;x=-188810000;
#10;x=-188800000;
#10;x=-188790000;
#10;x=-188780000;
#10;x=-188770000;
#10;x=-188760000;
#10;x=-188750000;
#10;x=-188740000;
#10;x=-188730000;
#10;x=-188720000;
#10;x=-188710000;
#10;x=-188700000;
#10;x=-188690000;
#10;x=-188680000;
#10;x=-188670000;
#10;x=-188660000;
#10;x=-188650000;
#10;x=-188640000;
#10;x=-188630000;
#10;x=-188620000;
#10;x=-188610000;
#10;x=-188600000;
#10;x=-188590000;
#10;x=-188580000;
#10;x=-188570000;
#10;x=-188560000;
#10;x=-188550000;
#10;x=-188540000;
#10;x=-188530000;
#10;x=-188520000;
#10;x=-188510000;
#10;x=-188500000;
#10;x=-188490000;
#10;x=-188480000;
#10;x=-188470000;
#10;x=-188460000;
#10;x=-188450000;
#10;x=-188440000;
#10;x=-188430000;
#10;x=-188420000;
#10;x=-188410000;
#10;x=-188400000;
#10;x=-188390000;
#10;x=-188380000;
#10;x=-188370000;
#10;x=-188360000;
#10;x=-188350000;
#10;x=-188340000;
#10;x=-188330000;
#10;x=-188320000;
#10;x=-188310000;
#10;x=-188300000;
#10;x=-188290000;
#10;x=-188280000;
#10;x=-188270000;
#10;x=-188260000;
#10;x=-188250000;
#10;x=-188240000;
#10;x=-188230000;
#10;x=-188220000;
#10;x=-188210000;
#10;x=-188200000;
#10;x=-188190000;
#10;x=-188180000;
#10;x=-188170000;
#10;x=-188160000;
#10;x=-188150000;
#10;x=-188140000;
#10;x=-188130000;
#10;x=-188120000;
#10;x=-188110000;
#10;x=-188100000;
#10;x=-188090000;
#10;x=-188080000;
#10;x=-188070000;
#10;x=-188060000;
#10;x=-188050000;
#10;x=-188040000;
#10;x=-188030000;
#10;x=-188020000;
#10;x=-188010000;
#10;x=-188000000;
#10;x=-187990000;
#10;x=-187980000;
#10;x=-187970000;
#10;x=-187960000;
#10;x=-187950000;
#10;x=-187940000;
#10;x=-187930000;
#10;x=-187920000;
#10;x=-187910000;
#10;x=-187900000;
#10;x=-187890000;
#10;x=-187880000;
#10;x=-187870000;
#10;x=-187860000;
#10;x=-187850000;
#10;x=-187840000;
#10;x=-187830000;
#10;x=-187820000;
#10;x=-187810000;
#10;x=-187800000;
#10;x=-187790000;
#10;x=-187780000;
#10;x=-187770000;
#10;x=-187760000;
#10;x=-187750000;
#10;x=-187740000;
#10;x=-187730000;
#10;x=-187720000;
#10;x=-187710000;
#10;x=-187700000;
#10;x=-187690000;
#10;x=-187680000;
#10;x=-187670000;
#10;x=-187660000;
#10;x=-187650000;
#10;x=-187640000;
#10;x=-187630000;
#10;x=-187620000;
#10;x=-187610000;
#10;x=-187600000;
#10;x=-187590000;
#10;x=-187580000;
#10;x=-187570000;
#10;x=-187560000;
#10;x=-187550000;
#10;x=-187540000;
#10;x=-187530000;
#10;x=-187520000;
#10;x=-187510000;
#10;x=-187500000;
#10;x=-187490000;
#10;x=-187480000;
#10;x=-187470000;
#10;x=-187460000;
#10;x=-187450000;
#10;x=-187440000;
#10;x=-187430000;
#10;x=-187420000;
#10;x=-187410000;
#10;x=-187400000;
#10;x=-187390000;
#10;x=-187380000;
#10;x=-187370000;
#10;x=-187360000;
#10;x=-187350000;
#10;x=-187340000;
#10;x=-187330000;
#10;x=-187320000;
#10;x=-187310000;
#10;x=-187300000;
#10;x=-187290000;
#10;x=-187280000;
#10;x=-187270000;
#10;x=-187260000;
#10;x=-187250000;
#10;x=-187240000;
#10;x=-187230000;
#10;x=-187220000;
#10;x=-187210000;
#10;x=-187200000;
#10;x=-187190000;
#10;x=-187180000;
#10;x=-187170000;
#10;x=-187160000;
#10;x=-187150000;
#10;x=-187140000;
#10;x=-187130000;
#10;x=-187120000;
#10;x=-187110000;
#10;x=-187100000;
#10;x=-187090000;
#10;x=-187080000;
#10;x=-187070000;
#10;x=-187060000;
#10;x=-187050000;
#10;x=-187040000;
#10;x=-187030000;
#10;x=-187020000;
#10;x=-187010000;
#10;x=-187000000;
#10;x=-186990000;
#10;x=-186980000;
#10;x=-186970000;
#10;x=-186960000;
#10;x=-186950000;
#10;x=-186940000;
#10;x=-186930000;
#10;x=-186920000;
#10;x=-186910000;
#10;x=-186900000;
#10;x=-186890000;
#10;x=-186880000;
#10;x=-186870000;
#10;x=-186860000;
#10;x=-186850000;
#10;x=-186840000;
#10;x=-186830000;
#10;x=-186820000;
#10;x=-186810000;
#10;x=-186800000;
#10;x=-186790000;
#10;x=-186780000;
#10;x=-186770000;
#10;x=-186760000;
#10;x=-186750000;
#10;x=-186740000;
#10;x=-186730000;
#10;x=-186720000;
#10;x=-186710000;
#10;x=-186700000;
#10;x=-186690000;
#10;x=-186680000;
#10;x=-186670000;
#10;x=-186660000;
#10;x=-186650000;
#10;x=-186640000;
#10;x=-186630000;
#10;x=-186620000;
#10;x=-186610000;
#10;x=-186600000;
#10;x=-186590000;
#10;x=-186580000;
#10;x=-186570000;
#10;x=-186560000;
#10;x=-186550000;
#10;x=-186540000;
#10;x=-186530000;
#10;x=-186520000;
#10;x=-186510000;
#10;x=-186500000;
#10;x=-186490000;
#10;x=-186480000;
#10;x=-186470000;
#10;x=-186460000;
#10;x=-186450000;
#10;x=-186440000;
#10;x=-186430000;
#10;x=-186420000;
#10;x=-186410000;
#10;x=-186400000;
#10;x=-186390000;
#10;x=-186380000;
#10;x=-186370000;
#10;x=-186360000;
#10;x=-186350000;
#10;x=-186340000;
#10;x=-186330000;
#10;x=-186320000;
#10;x=-186310000;
#10;x=-186300000;
#10;x=-186290000;
#10;x=-186280000;
#10;x=-186270000;
#10;x=-186260000;
#10;x=-186250000;
#10;x=-186240000;
#10;x=-186230000;
#10;x=-186220000;
#10;x=-186210000;
#10;x=-186200000;
#10;x=-186190000;
#10;x=-186180000;
#10;x=-186170000;
#10;x=-186160000;
#10;x=-186150000;
#10;x=-186140000;
#10;x=-186130000;
#10;x=-186120000;
#10;x=-186110000;
#10;x=-186100000;
#10;x=-186090000;
#10;x=-186080000;
#10;x=-186070000;
#10;x=-186060000;
#10;x=-186050000;
#10;x=-186040000;
#10;x=-186030000;
#10;x=-186020000;
#10;x=-186010000;
#10;x=-186000000;
#10;x=-185990000;
#10;x=-185980000;
#10;x=-185970000;
#10;x=-185960000;
#10;x=-185950000;
#10;x=-185940000;
#10;x=-185930000;
#10;x=-185920000;
#10;x=-185910000;
#10;x=-185900000;
#10;x=-185890000;
#10;x=-185880000;
#10;x=-185870000;
#10;x=-185860000;
#10;x=-185850000;
#10;x=-185840000;
#10;x=-185830000;
#10;x=-185820000;
#10;x=-185810000;
#10;x=-185800000;
#10;x=-185790000;
#10;x=-185780000;
#10;x=-185770000;
#10;x=-185760000;
#10;x=-185750000;
#10;x=-185740000;
#10;x=-185730000;
#10;x=-185720000;
#10;x=-185710000;
#10;x=-185700000;
#10;x=-185690000;
#10;x=-185680000;
#10;x=-185670000;
#10;x=-185660000;
#10;x=-185650000;
#10;x=-185640000;
#10;x=-185630000;
#10;x=-185620000;
#10;x=-185610000;
#10;x=-185600000;
#10;x=-185590000;
#10;x=-185580000;
#10;x=-185570000;
#10;x=-185560000;
#10;x=-185550000;
#10;x=-185540000;
#10;x=-185530000;
#10;x=-185520000;
#10;x=-185510000;
#10;x=-185500000;
#10;x=-185490000;
#10;x=-185480000;
#10;x=-185470000;
#10;x=-185460000;
#10;x=-185450000;
#10;x=-185440000;
#10;x=-185430000;
#10;x=-185420000;
#10;x=-185410000;
#10;x=-185400000;
#10;x=-185390000;
#10;x=-185380000;
#10;x=-185370000;
#10;x=-185360000;
#10;x=-185350000;
#10;x=-185340000;
#10;x=-185330000;
#10;x=-185320000;
#10;x=-185310000;
#10;x=-185300000;
#10;x=-185290000;
#10;x=-185280000;
#10;x=-185270000;
#10;x=-185260000;
#10;x=-185250000;
#10;x=-185240000;
#10;x=-185230000;
#10;x=-185220000;
#10;x=-185210000;
#10;x=-185200000;
#10;x=-185190000;
#10;x=-185180000;
#10;x=-185170000;
#10;x=-185160000;
#10;x=-185150000;
#10;x=-185140000;
#10;x=-185130000;
#10;x=-185120000;
#10;x=-185110000;
#10;x=-185100000;
#10;x=-185090000;
#10;x=-185080000;
#10;x=-185070000;
#10;x=-185060000;
#10;x=-185050000;
#10;x=-185040000;
#10;x=-185030000;
#10;x=-185020000;
#10;x=-185010000;
#10;x=-185000000;
#10;x=-184990000;
#10;x=-184980000;
#10;x=-184970000;
#10;x=-184960000;
#10;x=-184950000;
#10;x=-184940000;
#10;x=-184930000;
#10;x=-184920000;
#10;x=-184910000;
#10;x=-184900000;
#10;x=-184890000;
#10;x=-184880000;
#10;x=-184870000;
#10;x=-184860000;
#10;x=-184850000;
#10;x=-184840000;
#10;x=-184830000;
#10;x=-184820000;
#10;x=-184810000;
#10;x=-184800000;
#10;x=-184790000;
#10;x=-184780000;
#10;x=-184770000;
#10;x=-184760000;
#10;x=-184750000;
#10;x=-184740000;
#10;x=-184730000;
#10;x=-184720000;
#10;x=-184710000;
#10;x=-184700000;
#10;x=-184690000;
#10;x=-184680000;
#10;x=-184670000;
#10;x=-184660000;
#10;x=-184650000;
#10;x=-184640000;
#10;x=-184630000;
#10;x=-184620000;
#10;x=-184610000;
#10;x=-184600000;
#10;x=-184590000;
#10;x=-184580000;
#10;x=-184570000;
#10;x=-184560000;
#10;x=-184550000;
#10;x=-184540000;
#10;x=-184530000;
#10;x=-184520000;
#10;x=-184510000;
#10;x=-184500000;
#10;x=-184490000;
#10;x=-184480000;
#10;x=-184470000;
#10;x=-184460000;
#10;x=-184450000;
#10;x=-184440000;
#10;x=-184430000;
#10;x=-184420000;
#10;x=-184410000;
#10;x=-184400000;
#10;x=-184390000;
#10;x=-184380000;
#10;x=-184370000;
#10;x=-184360000;
#10;x=-184350000;
#10;x=-184340000;
#10;x=-184330000;
#10;x=-184320000;
#10;x=-184310000;
#10;x=-184300000;
#10;x=-184290000;
#10;x=-184280000;
#10;x=-184270000;
#10;x=-184260000;
#10;x=-184250000;
#10;x=-184240000;
#10;x=-184230000;
#10;x=-184220000;
#10;x=-184210000;
#10;x=-184200000;
#10;x=-184190000;
#10;x=-184180000;
#10;x=-184170000;
#10;x=-184160000;
#10;x=-184150000;
#10;x=-184140000;
#10;x=-184130000;
#10;x=-184120000;
#10;x=-184110000;
#10;x=-184100000;
#10;x=-184090000;
#10;x=-184080000;
#10;x=-184070000;
#10;x=-184060000;
#10;x=-184050000;
#10;x=-184040000;
#10;x=-184030000;
#10;x=-184020000;
#10;x=-184010000;
#10;x=-184000000;
#10;x=-183990000;
#10;x=-183980000;
#10;x=-183970000;
#10;x=-183960000;
#10;x=-183950000;
#10;x=-183940000;
#10;x=-183930000;
#10;x=-183920000;
#10;x=-183910000;
#10;x=-183900000;
#10;x=-183890000;
#10;x=-183880000;
#10;x=-183870000;
#10;x=-183860000;
#10;x=-183850000;
#10;x=-183840000;
#10;x=-183830000;
#10;x=-183820000;
#10;x=-183810000;
#10;x=-183800000;
#10;x=-183790000;
#10;x=-183780000;
#10;x=-183770000;
#10;x=-183760000;
#10;x=-183750000;
#10;x=-183740000;
#10;x=-183730000;
#10;x=-183720000;
#10;x=-183710000;
#10;x=-183700000;
#10;x=-183690000;
#10;x=-183680000;
#10;x=-183670000;
#10;x=-183660000;
#10;x=-183650000;
#10;x=-183640000;
#10;x=-183630000;
#10;x=-183620000;
#10;x=-183610000;
#10;x=-183600000;
#10;x=-183590000;
#10;x=-183580000;
#10;x=-183570000;
#10;x=-183560000;
#10;x=-183550000;
#10;x=-183540000;
#10;x=-183530000;
#10;x=-183520000;
#10;x=-183510000;
#10;x=-183500000;
#10;x=-183490000;
#10;x=-183480000;
#10;x=-183470000;
#10;x=-183460000;
#10;x=-183450000;
#10;x=-183440000;
#10;x=-183430000;
#10;x=-183420000;
#10;x=-183410000;
#10;x=-183400000;
#10;x=-183390000;
#10;x=-183380000;
#10;x=-183370000;
#10;x=-183360000;
#10;x=-183350000;
#10;x=-183340000;
#10;x=-183330000;
#10;x=-183320000;
#10;x=-183310000;
#10;x=-183300000;
#10;x=-183290000;
#10;x=-183280000;
#10;x=-183270000;
#10;x=-183260000;
#10;x=-183250000;
#10;x=-183240000;
#10;x=-183230000;
#10;x=-183220000;
#10;x=-183210000;
#10;x=-183200000;
#10;x=-183190000;
#10;x=-183180000;
#10;x=-183170000;
#10;x=-183160000;
#10;x=-183150000;
#10;x=-183140000;
#10;x=-183130000;
#10;x=-183120000;
#10;x=-183110000;
#10;x=-183100000;
#10;x=-183090000;
#10;x=-183080000;
#10;x=-183070000;
#10;x=-183060000;
#10;x=-183050000;
#10;x=-183040000;
#10;x=-183030000;
#10;x=-183020000;
#10;x=-183010000;
#10;x=-183000000;
#10;x=-182990000;
#10;x=-182980000;
#10;x=-182970000;
#10;x=-182960000;
#10;x=-182950000;
#10;x=-182940000;
#10;x=-182930000;
#10;x=-182920000;
#10;x=-182910000;
#10;x=-182900000;
#10;x=-182890000;
#10;x=-182880000;
#10;x=-182870000;
#10;x=-182860000;
#10;x=-182850000;
#10;x=-182840000;
#10;x=-182830000;
#10;x=-182820000;
#10;x=-182810000;
#10;x=-182800000;
#10;x=-182790000;
#10;x=-182780000;
#10;x=-182770000;
#10;x=-182760000;
#10;x=-182750000;
#10;x=-182740000;
#10;x=-182730000;
#10;x=-182720000;
#10;x=-182710000;
#10;x=-182700000;
#10;x=-182690000;
#10;x=-182680000;
#10;x=-182670000;
#10;x=-182660000;
#10;x=-182650000;
#10;x=-182640000;
#10;x=-182630000;
#10;x=-182620000;
#10;x=-182610000;
#10;x=-182600000;
#10;x=-182590000;
#10;x=-182580000;
#10;x=-182570000;
#10;x=-182560000;
#10;x=-182550000;
#10;x=-182540000;
#10;x=-182530000;
#10;x=-182520000;
#10;x=-182510000;
#10;x=-182500000;
#10;x=-182490000;
#10;x=-182480000;
#10;x=-182470000;
#10;x=-182460000;
#10;x=-182450000;
#10;x=-182440000;
#10;x=-182430000;
#10;x=-182420000;
#10;x=-182410000;
#10;x=-182400000;
#10;x=-182390000;
#10;x=-182380000;
#10;x=-182370000;
#10;x=-182360000;
#10;x=-182350000;
#10;x=-182340000;
#10;x=-182330000;
#10;x=-182320000;
#10;x=-182310000;
#10;x=-182300000;
#10;x=-182290000;
#10;x=-182280000;
#10;x=-182270000;
#10;x=-182260000;
#10;x=-182250000;
#10;x=-182240000;
#10;x=-182230000;
#10;x=-182220000;
#10;x=-182210000;
#10;x=-182200000;
#10;x=-182190000;
#10;x=-182180000;
#10;x=-182170000;
#10;x=-182160000;
#10;x=-182150000;
#10;x=-182140000;
#10;x=-182130000;
#10;x=-182120000;
#10;x=-182110000;
#10;x=-182100000;
#10;x=-182090000;
#10;x=-182080000;
#10;x=-182070000;
#10;x=-182060000;
#10;x=-182050000;
#10;x=-182040000;
#10;x=-182030000;
#10;x=-182020000;
#10;x=-182010000;
#10;x=-182000000;
#10;x=-181990000;
#10;x=-181980000;
#10;x=-181970000;
#10;x=-181960000;
#10;x=-181950000;
#10;x=-181940000;
#10;x=-181930000;
#10;x=-181920000;
#10;x=-181910000;
#10;x=-181900000;
#10;x=-181890000;
#10;x=-181880000;
#10;x=-181870000;
#10;x=-181860000;
#10;x=-181850000;
#10;x=-181840000;
#10;x=-181830000;
#10;x=-181820000;
#10;x=-181810000;
#10;x=-181800000;
#10;x=-181790000;
#10;x=-181780000;
#10;x=-181770000;
#10;x=-181760000;
#10;x=-181750000;
#10;x=-181740000;
#10;x=-181730000;
#10;x=-181720000;
#10;x=-181710000;
#10;x=-181700000;
#10;x=-181690000;
#10;x=-181680000;
#10;x=-181670000;
#10;x=-181660000;
#10;x=-181650000;
#10;x=-181640000;
#10;x=-181630000;
#10;x=-181620000;
#10;x=-181610000;
#10;x=-181600000;
#10;x=-181590000;
#10;x=-181580000;
#10;x=-181570000;
#10;x=-181560000;
#10;x=-181550000;
#10;x=-181540000;
#10;x=-181530000;
#10;x=-181520000;
#10;x=-181510000;
#10;x=-181500000;
#10;x=-181490000;
#10;x=-181480000;
#10;x=-181470000;
#10;x=-181460000;
#10;x=-181450000;
#10;x=-181440000;
#10;x=-181430000;
#10;x=-181420000;
#10;x=-181410000;
#10;x=-181400000;
#10;x=-181390000;
#10;x=-181380000;
#10;x=-181370000;
#10;x=-181360000;
#10;x=-181350000;
#10;x=-181340000;
#10;x=-181330000;
#10;x=-181320000;
#10;x=-181310000;
#10;x=-181300000;
#10;x=-181290000;
#10;x=-181280000;
#10;x=-181270000;
#10;x=-181260000;
#10;x=-181250000;
#10;x=-181240000;
#10;x=-181230000;
#10;x=-181220000;
#10;x=-181210000;
#10;x=-181200000;
#10;x=-181190000;
#10;x=-181180000;
#10;x=-181170000;
#10;x=-181160000;
#10;x=-181150000;
#10;x=-181140000;
#10;x=-181130000;
#10;x=-181120000;
#10;x=-181110000;
#10;x=-181100000;
#10;x=-181090000;
#10;x=-181080000;
#10;x=-181070000;
#10;x=-181060000;
#10;x=-181050000;
#10;x=-181040000;
#10;x=-181030000;
#10;x=-181020000;
#10;x=-181010000;
#10;x=-181000000;
#10;x=-180990000;
#10;x=-180980000;
#10;x=-180970000;
#10;x=-180960000;
#10;x=-180950000;
#10;x=-180940000;
#10;x=-180930000;
#10;x=-180920000;
#10;x=-180910000;
#10;x=-180900000;
#10;x=-180890000;
#10;x=-180880000;
#10;x=-180870000;
#10;x=-180860000;
#10;x=-180850000;
#10;x=-180840000;
#10;x=-180830000;
#10;x=-180820000;
#10;x=-180810000;
#10;x=-180800000;
#10;x=-180790000;
#10;x=-180780000;
#10;x=-180770000;
#10;x=-180760000;
#10;x=-180750000;
#10;x=-180740000;
#10;x=-180730000;
#10;x=-180720000;
#10;x=-180710000;
#10;x=-180700000;
#10;x=-180690000;
#10;x=-180680000;
#10;x=-180670000;
#10;x=-180660000;
#10;x=-180650000;
#10;x=-180640000;
#10;x=-180630000;
#10;x=-180620000;
#10;x=-180610000;
#10;x=-180600000;
#10;x=-180590000;
#10;x=-180580000;
#10;x=-180570000;
#10;x=-180560000;
#10;x=-180550000;
#10;x=-180540000;
#10;x=-180530000;
#10;x=-180520000;
#10;x=-180510000;
#10;x=-180500000;
#10;x=-180490000;
#10;x=-180480000;
#10;x=-180470000;
#10;x=-180460000;
#10;x=-180450000;
#10;x=-180440000;
#10;x=-180430000;
#10;x=-180420000;
#10;x=-180410000;
#10;x=-180400000;
#10;x=-180390000;
#10;x=-180380000;
#10;x=-180370000;
#10;x=-180360000;
#10;x=-180350000;
#10;x=-180340000;
#10;x=-180330000;
#10;x=-180320000;
#10;x=-180310000;
#10;x=-180300000;
#10;x=-180290000;
#10;x=-180280000;
#10;x=-180270000;
#10;x=-180260000;
#10;x=-180250000;
#10;x=-180240000;
#10;x=-180230000;
#10;x=-180220000;
#10;x=-180210000;
#10;x=-180200000;
#10;x=-180190000;
#10;x=-180180000;
#10;x=-180170000;
#10;x=-180160000;
#10;x=-180150000;
#10;x=-180140000;
#10;x=-180130000;
#10;x=-180120000;
#10;x=-180110000;
#10;x=-180100000;
#10;x=-180090000;
#10;x=-180080000;
#10;x=-180070000;
#10;x=-180060000;
#10;x=-180050000;
#10;x=-180040000;
#10;x=-180030000;
#10;x=-180020000;
#10;x=-180010000;
#10;x=-180000000;
#10;x=-179990000;
#10;x=-179980000;
#10;x=-179970000;
#10;x=-179960000;
#10;x=-179950000;
#10;x=-179940000;
#10;x=-179930000;
#10;x=-179920000;
#10;x=-179910000;
#10;x=-179900000;
#10;x=-179890000;
#10;x=-179880000;
#10;x=-179870000;
#10;x=-179860000;
#10;x=-179850000;
#10;x=-179840000;
#10;x=-179830000;
#10;x=-179820000;
#10;x=-179810000;
#10;x=-179800000;
#10;x=-179790000;
#10;x=-179780000;
#10;x=-179770000;
#10;x=-179760000;
#10;x=-179750000;
#10;x=-179740000;
#10;x=-179730000;
#10;x=-179720000;
#10;x=-179710000;
#10;x=-179700000;
#10;x=-179690000;
#10;x=-179680000;
#10;x=-179670000;
#10;x=-179660000;
#10;x=-179650000;
#10;x=-179640000;
#10;x=-179630000;
#10;x=-179620000;
#10;x=-179610000;
#10;x=-179600000;
#10;x=-179590000;
#10;x=-179580000;
#10;x=-179570000;
#10;x=-179560000;
#10;x=-179550000;
#10;x=-179540000;
#10;x=-179530000;
#10;x=-179520000;
#10;x=-179510000;
#10;x=-179500000;
#10;x=-179490000;
#10;x=-179480000;
#10;x=-179470000;
#10;x=-179460000;
#10;x=-179450000;
#10;x=-179440000;
#10;x=-179430000;
#10;x=-179420000;
#10;x=-179410000;
#10;x=-179400000;
#10;x=-179390000;
#10;x=-179380000;
#10;x=-179370000;
#10;x=-179360000;
#10;x=-179350000;
#10;x=-179340000;
#10;x=-179330000;
#10;x=-179320000;
#10;x=-179310000;
#10;x=-179300000;
#10;x=-179290000;
#10;x=-179280000;
#10;x=-179270000;
#10;x=-179260000;
#10;x=-179250000;
#10;x=-179240000;
#10;x=-179230000;
#10;x=-179220000;
#10;x=-179210000;
#10;x=-179200000;
#10;x=-179190000;
#10;x=-179180000;
#10;x=-179170000;
#10;x=-179160000;
#10;x=-179150000;
#10;x=-179140000;
#10;x=-179130000;
#10;x=-179120000;
#10;x=-179110000;
#10;x=-179100000;
#10;x=-179090000;
#10;x=-179080000;
#10;x=-179070000;
#10;x=-179060000;
#10;x=-179050000;
#10;x=-179040000;
#10;x=-179030000;
#10;x=-179020000;
#10;x=-179010000;
#10;x=-179000000;
#10;x=-178990000;
#10;x=-178980000;
#10;x=-178970000;
#10;x=-178960000;
#10;x=-178950000;
#10;x=-178940000;
#10;x=-178930000;
#10;x=-178920000;
#10;x=-178910000;
#10;x=-178900000;
#10;x=-178890000;
#10;x=-178880000;
#10;x=-178870000;
#10;x=-178860000;
#10;x=-178850000;
#10;x=-178840000;
#10;x=-178830000;
#10;x=-178820000;
#10;x=-178810000;
#10;x=-178800000;
#10;x=-178790000;
#10;x=-178780000;
#10;x=-178770000;
#10;x=-178760000;
#10;x=-178750000;
#10;x=-178740000;
#10;x=-178730000;
#10;x=-178720000;
#10;x=-178710000;
#10;x=-178700000;
#10;x=-178690000;
#10;x=-178680000;
#10;x=-178670000;
#10;x=-178660000;
#10;x=-178650000;
#10;x=-178640000;
#10;x=-178630000;
#10;x=-178620000;
#10;x=-178610000;
#10;x=-178600000;
#10;x=-178590000;
#10;x=-178580000;
#10;x=-178570000;
#10;x=-178560000;
#10;x=-178550000;
#10;x=-178540000;
#10;x=-178530000;
#10;x=-178520000;
#10;x=-178510000;
#10;x=-178500000;
#10;x=-178490000;
#10;x=-178480000;
#10;x=-178470000;
#10;x=-178460000;
#10;x=-178450000;
#10;x=-178440000;
#10;x=-178430000;
#10;x=-178420000;
#10;x=-178410000;
#10;x=-178400000;
#10;x=-178390000;
#10;x=-178380000;
#10;x=-178370000;
#10;x=-178360000;
#10;x=-178350000;
#10;x=-178340000;
#10;x=-178330000;
#10;x=-178320000;
#10;x=-178310000;
#10;x=-178300000;
#10;x=-178290000;
#10;x=-178280000;
#10;x=-178270000;
#10;x=-178260000;
#10;x=-178250000;
#10;x=-178240000;
#10;x=-178230000;
#10;x=-178220000;
#10;x=-178210000;
#10;x=-178200000;
#10;x=-178190000;
#10;x=-178180000;
#10;x=-178170000;
#10;x=-178160000;
#10;x=-178150000;
#10;x=-178140000;
#10;x=-178130000;
#10;x=-178120000;
#10;x=-178110000;
#10;x=-178100000;
#10;x=-178090000;
#10;x=-178080000;
#10;x=-178070000;
#10;x=-178060000;
#10;x=-178050000;
#10;x=-178040000;
#10;x=-178030000;
#10;x=-178020000;
#10;x=-178010000;
#10;x=-178000000;
#10;x=-177990000;
#10;x=-177980000;
#10;x=-177970000;
#10;x=-177960000;
#10;x=-177950000;
#10;x=-177940000;
#10;x=-177930000;
#10;x=-177920000;
#10;x=-177910000;
#10;x=-177900000;
#10;x=-177890000;
#10;x=-177880000;
#10;x=-177870000;
#10;x=-177860000;
#10;x=-177850000;
#10;x=-177840000;
#10;x=-177830000;
#10;x=-177820000;
#10;x=-177810000;
#10;x=-177800000;
#10;x=-177790000;
#10;x=-177780000;
#10;x=-177770000;
#10;x=-177760000;
#10;x=-177750000;
#10;x=-177740000;
#10;x=-177730000;
#10;x=-177720000;
#10;x=-177710000;
#10;x=-177700000;
#10;x=-177690000;
#10;x=-177680000;
#10;x=-177670000;
#10;x=-177660000;
#10;x=-177650000;
#10;x=-177640000;
#10;x=-177630000;
#10;x=-177620000;
#10;x=-177610000;
#10;x=-177600000;
#10;x=-177590000;
#10;x=-177580000;
#10;x=-177570000;
#10;x=-177560000;
#10;x=-177550000;
#10;x=-177540000;
#10;x=-177530000;
#10;x=-177520000;
#10;x=-177510000;
#10;x=-177500000;
#10;x=-177490000;
#10;x=-177480000;
#10;x=-177470000;
#10;x=-177460000;
#10;x=-177450000;
#10;x=-177440000;
#10;x=-177430000;
#10;x=-177420000;
#10;x=-177410000;
#10;x=-177400000;
#10;x=-177390000;
#10;x=-177380000;
#10;x=-177370000;
#10;x=-177360000;
#10;x=-177350000;
#10;x=-177340000;
#10;x=-177330000;
#10;x=-177320000;
#10;x=-177310000;
#10;x=-177300000;
#10;x=-177290000;
#10;x=-177280000;
#10;x=-177270000;
#10;x=-177260000;
#10;x=-177250000;
#10;x=-177240000;
#10;x=-177230000;
#10;x=-177220000;
#10;x=-177210000;
#10;x=-177200000;
#10;x=-177190000;
#10;x=-177180000;
#10;x=-177170000;
#10;x=-177160000;
#10;x=-177150000;
#10;x=-177140000;
#10;x=-177130000;
#10;x=-177120000;
#10;x=-177110000;
#10;x=-177100000;
#10;x=-177090000;
#10;x=-177080000;
#10;x=-177070000;
#10;x=-177060000;
#10;x=-177050000;
#10;x=-177040000;
#10;x=-177030000;
#10;x=-177020000;
#10;x=-177010000;
#10;x=-177000000;
#10;x=-176990000;
#10;x=-176980000;
#10;x=-176970000;
#10;x=-176960000;
#10;x=-176950000;
#10;x=-176940000;
#10;x=-176930000;
#10;x=-176920000;
#10;x=-176910000;
#10;x=-176900000;
#10;x=-176890000;
#10;x=-176880000;
#10;x=-176870000;
#10;x=-176860000;
#10;x=-176850000;
#10;x=-176840000;
#10;x=-176830000;
#10;x=-176820000;
#10;x=-176810000;
#10;x=-176800000;
#10;x=-176790000;
#10;x=-176780000;
#10;x=-176770000;
#10;x=-176760000;
#10;x=-176750000;
#10;x=-176740000;
#10;x=-176730000;
#10;x=-176720000;
#10;x=-176710000;
#10;x=-176700000;
#10;x=-176690000;
#10;x=-176680000;
#10;x=-176670000;
#10;x=-176660000;
#10;x=-176650000;
#10;x=-176640000;
#10;x=-176630000;
#10;x=-176620000;
#10;x=-176610000;
#10;x=-176600000;
#10;x=-176590000;
#10;x=-176580000;
#10;x=-176570000;
#10;x=-176560000;
#10;x=-176550000;
#10;x=-176540000;
#10;x=-176530000;
#10;x=-176520000;
#10;x=-176510000;
#10;x=-176500000;
#10;x=-176490000;
#10;x=-176480000;
#10;x=-176470000;
#10;x=-176460000;
#10;x=-176450000;
#10;x=-176440000;
#10;x=-176430000;
#10;x=-176420000;
#10;x=-176410000;
#10;x=-176400000;
#10;x=-176390000;
#10;x=-176380000;
#10;x=-176370000;
#10;x=-176360000;
#10;x=-176350000;
#10;x=-176340000;
#10;x=-176330000;
#10;x=-176320000;
#10;x=-176310000;
#10;x=-176300000;
#10;x=-176290000;
#10;x=-176280000;
#10;x=-176270000;
#10;x=-176260000;
#10;x=-176250000;
#10;x=-176240000;
#10;x=-176230000;
#10;x=-176220000;
#10;x=-176210000;
#10;x=-176200000;
#10;x=-176190000;
#10;x=-176180000;
#10;x=-176170000;
#10;x=-176160000;
#10;x=-176150000;
#10;x=-176140000;
#10;x=-176130000;
#10;x=-176120000;
#10;x=-176110000;
#10;x=-176100000;
#10;x=-176090000;
#10;x=-176080000;
#10;x=-176070000;
#10;x=-176060000;
#10;x=-176050000;
#10;x=-176040000;
#10;x=-176030000;
#10;x=-176020000;
#10;x=-176010000;
#10;x=-176000000;
#10;x=-175990000;
#10;x=-175980000;
#10;x=-175970000;
#10;x=-175960000;
#10;x=-175950000;
#10;x=-175940000;
#10;x=-175930000;
#10;x=-175920000;
#10;x=-175910000;
#10;x=-175900000;
#10;x=-175890000;
#10;x=-175880000;
#10;x=-175870000;
#10;x=-175860000;
#10;x=-175850000;
#10;x=-175840000;
#10;x=-175830000;
#10;x=-175820000;
#10;x=-175810000;
#10;x=-175800000;
#10;x=-175790000;
#10;x=-175780000;
#10;x=-175770000;
#10;x=-175760000;
#10;x=-175750000;
#10;x=-175740000;
#10;x=-175730000;
#10;x=-175720000;
#10;x=-175710000;
#10;x=-175700000;
#10;x=-175690000;
#10;x=-175680000;
#10;x=-175670000;
#10;x=-175660000;
#10;x=-175650000;
#10;x=-175640000;
#10;x=-175630000;
#10;x=-175620000;
#10;x=-175610000;
#10;x=-175600000;
#10;x=-175590000;
#10;x=-175580000;
#10;x=-175570000;
#10;x=-175560000;
#10;x=-175550000;
#10;x=-175540000;
#10;x=-175530000;
#10;x=-175520000;
#10;x=-175510000;
#10;x=-175500000;
#10;x=-175490000;
#10;x=-175480000;
#10;x=-175470000;
#10;x=-175460000;
#10;x=-175450000;
#10;x=-175440000;
#10;x=-175430000;
#10;x=-175420000;
#10;x=-175410000;
#10;x=-175400000;
#10;x=-175390000;
#10;x=-175380000;
#10;x=-175370000;
#10;x=-175360000;
#10;x=-175350000;
#10;x=-175340000;
#10;x=-175330000;
#10;x=-175320000;
#10;x=-175310000;
#10;x=-175300000;
#10;x=-175290000;
#10;x=-175280000;
#10;x=-175270000;
#10;x=-175260000;
#10;x=-175250000;
#10;x=-175240000;
#10;x=-175230000;
#10;x=-175220000;
#10;x=-175210000;
#10;x=-175200000;
#10;x=-175190000;
#10;x=-175180000;
#10;x=-175170000;
#10;x=-175160000;
#10;x=-175150000;
#10;x=-175140000;
#10;x=-175130000;
#10;x=-175120000;
#10;x=-175110000;
#10;x=-175100000;
#10;x=-175090000;
#10;x=-175080000;
#10;x=-175070000;
#10;x=-175060000;
#10;x=-175050000;
#10;x=-175040000;
#10;x=-175030000;
#10;x=-175020000;
#10;x=-175010000;
#10;x=-175000000;
#10;x=-174990000;
#10;x=-174980000;
#10;x=-174970000;
#10;x=-174960000;
#10;x=-174950000;
#10;x=-174940000;
#10;x=-174930000;
#10;x=-174920000;
#10;x=-174910000;
#10;x=-174900000;
#10;x=-174890000;
#10;x=-174880000;
#10;x=-174870000;
#10;x=-174860000;
#10;x=-174850000;
#10;x=-174840000;
#10;x=-174830000;
#10;x=-174820000;
#10;x=-174810000;
#10;x=-174800000;
#10;x=-174790000;
#10;x=-174780000;
#10;x=-174770000;
#10;x=-174760000;
#10;x=-174750000;
#10;x=-174740000;
#10;x=-174730000;
#10;x=-174720000;
#10;x=-174710000;
#10;x=-174700000;
#10;x=-174690000;
#10;x=-174680000;
#10;x=-174670000;
#10;x=-174660000;
#10;x=-174650000;
#10;x=-174640000;
#10;x=-174630000;
#10;x=-174620000;
#10;x=-174610000;
#10;x=-174600000;
#10;x=-174590000;
#10;x=-174580000;
#10;x=-174570000;
#10;x=-174560000;
#10;x=-174550000;
#10;x=-174540000;
#10;x=-174530000;
#10;x=-174520000;
#10;x=-174510000;
#10;x=-174500000;
#10;x=-174490000;
#10;x=-174480000;
#10;x=-174470000;
#10;x=-174460000;
#10;x=-174450000;
#10;x=-174440000;
#10;x=-174430000;
#10;x=-174420000;
#10;x=-174410000;
#10;x=-174400000;
#10;x=-174390000;
#10;x=-174380000;
#10;x=-174370000;
#10;x=-174360000;
#10;x=-174350000;
#10;x=-174340000;
#10;x=-174330000;
#10;x=-174320000;
#10;x=-174310000;
#10;x=-174300000;
#10;x=-174290000;
#10;x=-174280000;
#10;x=-174270000;
#10;x=-174260000;
#10;x=-174250000;
#10;x=-174240000;
#10;x=-174230000;
#10;x=-174220000;
#10;x=-174210000;
#10;x=-174200000;
#10;x=-174190000;
#10;x=-174180000;
#10;x=-174170000;
#10;x=-174160000;
#10;x=-174150000;
#10;x=-174140000;
#10;x=-174130000;
#10;x=-174120000;
#10;x=-174110000;
#10;x=-174100000;
#10;x=-174090000;
#10;x=-174080000;
#10;x=-174070000;
#10;x=-174060000;
#10;x=-174050000;
#10;x=-174040000;
#10;x=-174030000;
#10;x=-174020000;
#10;x=-174010000;
#10;x=-174000000;
#10;x=-173990000;
#10;x=-173980000;
#10;x=-173970000;
#10;x=-173960000;
#10;x=-173950000;
#10;x=-173940000;
#10;x=-173930000;
#10;x=-173920000;
#10;x=-173910000;
#10;x=-173900000;
#10;x=-173890000;
#10;x=-173880000;
#10;x=-173870000;
#10;x=-173860000;
#10;x=-173850000;
#10;x=-173840000;
#10;x=-173830000;
#10;x=-173820000;
#10;x=-173810000;
#10;x=-173800000;
#10;x=-173790000;
#10;x=-173780000;
#10;x=-173770000;
#10;x=-173760000;
#10;x=-173750000;
#10;x=-173740000;
#10;x=-173730000;
#10;x=-173720000;
#10;x=-173710000;
#10;x=-173700000;
#10;x=-173690000;
#10;x=-173680000;
#10;x=-173670000;
#10;x=-173660000;
#10;x=-173650000;
#10;x=-173640000;
#10;x=-173630000;
#10;x=-173620000;
#10;x=-173610000;
#10;x=-173600000;
#10;x=-173590000;
#10;x=-173580000;
#10;x=-173570000;
#10;x=-173560000;
#10;x=-173550000;
#10;x=-173540000;
#10;x=-173530000;
#10;x=-173520000;
#10;x=-173510000;
#10;x=-173500000;
#10;x=-173490000;
#10;x=-173480000;
#10;x=-173470000;
#10;x=-173460000;
#10;x=-173450000;
#10;x=-173440000;
#10;x=-173430000;
#10;x=-173420000;
#10;x=-173410000;
#10;x=-173400000;
#10;x=-173390000;
#10;x=-173380000;
#10;x=-173370000;
#10;x=-173360000;
#10;x=-173350000;
#10;x=-173340000;
#10;x=-173330000;
#10;x=-173320000;
#10;x=-173310000;
#10;x=-173300000;
#10;x=-173290000;
#10;x=-173280000;
#10;x=-173270000;
#10;x=-173260000;
#10;x=-173250000;
#10;x=-173240000;
#10;x=-173230000;
#10;x=-173220000;
#10;x=-173210000;
#10;x=-173200000;
#10;x=-173190000;
#10;x=-173180000;
#10;x=-173170000;
#10;x=-173160000;
#10;x=-173150000;
#10;x=-173140000;
#10;x=-173130000;
#10;x=-173120000;
#10;x=-173110000;
#10;x=-173100000;
#10;x=-173090000;
#10;x=-173080000;
#10;x=-173070000;
#10;x=-173060000;
#10;x=-173050000;
#10;x=-173040000;
#10;x=-173030000;
#10;x=-173020000;
#10;x=-173010000;
#10;x=-173000000;
#10;x=-172990000;
#10;x=-172980000;
#10;x=-172970000;
#10;x=-172960000;
#10;x=-172950000;
#10;x=-172940000;
#10;x=-172930000;
#10;x=-172920000;
#10;x=-172910000;
#10;x=-172900000;
#10;x=-172890000;
#10;x=-172880000;
#10;x=-172870000;
#10;x=-172860000;
#10;x=-172850000;
#10;x=-172840000;
#10;x=-172830000;
#10;x=-172820000;
#10;x=-172810000;
#10;x=-172800000;
#10;x=-172790000;
#10;x=-172780000;
#10;x=-172770000;
#10;x=-172760000;
#10;x=-172750000;
#10;x=-172740000;
#10;x=-172730000;
#10;x=-172720000;
#10;x=-172710000;
#10;x=-172700000;
#10;x=-172690000;
#10;x=-172680000;
#10;x=-172670000;
#10;x=-172660000;
#10;x=-172650000;
#10;x=-172640000;
#10;x=-172630000;
#10;x=-172620000;
#10;x=-172610000;
#10;x=-172600000;
#10;x=-172590000;
#10;x=-172580000;
#10;x=-172570000;
#10;x=-172560000;
#10;x=-172550000;
#10;x=-172540000;
#10;x=-172530000;
#10;x=-172520000;
#10;x=-172510000;
#10;x=-172500000;
#10;x=-172490000;
#10;x=-172480000;
#10;x=-172470000;
#10;x=-172460000;
#10;x=-172450000;
#10;x=-172440000;
#10;x=-172430000;
#10;x=-172420000;
#10;x=-172410000;
#10;x=-172400000;
#10;x=-172390000;
#10;x=-172380000;
#10;x=-172370000;
#10;x=-172360000;
#10;x=-172350000;
#10;x=-172340000;
#10;x=-172330000;
#10;x=-172320000;
#10;x=-172310000;
#10;x=-172300000;
#10;x=-172290000;
#10;x=-172280000;
#10;x=-172270000;
#10;x=-172260000;
#10;x=-172250000;
#10;x=-172240000;
#10;x=-172230000;
#10;x=-172220000;
#10;x=-172210000;
#10;x=-172200000;
#10;x=-172190000;
#10;x=-172180000;
#10;x=-172170000;
#10;x=-172160000;
#10;x=-172150000;
#10;x=-172140000;
#10;x=-172130000;
#10;x=-172120000;
#10;x=-172110000;
#10;x=-172100000;
#10;x=-172090000;
#10;x=-172080000;
#10;x=-172070000;
#10;x=-172060000;
#10;x=-172050000;
#10;x=-172040000;
#10;x=-172030000;
#10;x=-172020000;
#10;x=-172010000;
#10;x=-172000000;
#10;x=-171990000;
#10;x=-171980000;
#10;x=-171970000;
#10;x=-171960000;
#10;x=-171950000;
#10;x=-171940000;
#10;x=-171930000;
#10;x=-171920000;
#10;x=-171910000;
#10;x=-171900000;
#10;x=-171890000;
#10;x=-171880000;
#10;x=-171870000;
#10;x=-171860000;
#10;x=-171850000;
#10;x=-171840000;
#10;x=-171830000;
#10;x=-171820000;
#10;x=-171810000;
#10;x=-171800000;
#10;x=-171790000;
#10;x=-171780000;
#10;x=-171770000;
#10;x=-171760000;
#10;x=-171750000;
#10;x=-171740000;
#10;x=-171730000;
#10;x=-171720000;
#10;x=-171710000;
#10;x=-171700000;
#10;x=-171690000;
#10;x=-171680000;
#10;x=-171670000;
#10;x=-171660000;
#10;x=-171650000;
#10;x=-171640000;
#10;x=-171630000;
#10;x=-171620000;
#10;x=-171610000;
#10;x=-171600000;
#10;x=-171590000;
#10;x=-171580000;
#10;x=-171570000;
#10;x=-171560000;
#10;x=-171550000;
#10;x=-171540000;
#10;x=-171530000;
#10;x=-171520000;
#10;x=-171510000;
#10;x=-171500000;
#10;x=-171490000;
#10;x=-171480000;
#10;x=-171470000;
#10;x=-171460000;
#10;x=-171450000;
#10;x=-171440000;
#10;x=-171430000;
#10;x=-171420000;
#10;x=-171410000;
#10;x=-171400000;
#10;x=-171390000;
#10;x=-171380000;
#10;x=-171370000;
#10;x=-171360000;
#10;x=-171350000;
#10;x=-171340000;
#10;x=-171330000;
#10;x=-171320000;
#10;x=-171310000;
#10;x=-171300000;
#10;x=-171290000;
#10;x=-171280000;
#10;x=-171270000;
#10;x=-171260000;
#10;x=-171250000;
#10;x=-171240000;
#10;x=-171230000;
#10;x=-171220000;
#10;x=-171210000;
#10;x=-171200000;
#10;x=-171190000;
#10;x=-171180000;
#10;x=-171170000;
#10;x=-171160000;
#10;x=-171150000;
#10;x=-171140000;
#10;x=-171130000;
#10;x=-171120000;
#10;x=-171110000;
#10;x=-171100000;
#10;x=-171090000;
#10;x=-171080000;
#10;x=-171070000;
#10;x=-171060000;
#10;x=-171050000;
#10;x=-171040000;
#10;x=-171030000;
#10;x=-171020000;
#10;x=-171010000;
#10;x=-171000000;
#10;x=-170990000;
#10;x=-170980000;
#10;x=-170970000;
#10;x=-170960000;
#10;x=-170950000;
#10;x=-170940000;
#10;x=-170930000;
#10;x=-170920000;
#10;x=-170910000;
#10;x=-170900000;
#10;x=-170890000;
#10;x=-170880000;
#10;x=-170870000;
#10;x=-170860000;
#10;x=-170850000;
#10;x=-170840000;
#10;x=-170830000;
#10;x=-170820000;
#10;x=-170810000;
#10;x=-170800000;
#10;x=-170790000;
#10;x=-170780000;
#10;x=-170770000;
#10;x=-170760000;
#10;x=-170750000;
#10;x=-170740000;
#10;x=-170730000;
#10;x=-170720000;
#10;x=-170710000;
#10;x=-170700000;
#10;x=-170690000;
#10;x=-170680000;
#10;x=-170670000;
#10;x=-170660000;
#10;x=-170650000;
#10;x=-170640000;
#10;x=-170630000;
#10;x=-170620000;
#10;x=-170610000;
#10;x=-170600000;
#10;x=-170590000;
#10;x=-170580000;
#10;x=-170570000;
#10;x=-170560000;
#10;x=-170550000;
#10;x=-170540000;
#10;x=-170530000;
#10;x=-170520000;
#10;x=-170510000;
#10;x=-170500000;
#10;x=-170490000;
#10;x=-170480000;
#10;x=-170470000;
#10;x=-170460000;
#10;x=-170450000;
#10;x=-170440000;
#10;x=-170430000;
#10;x=-170420000;
#10;x=-170410000;
#10;x=-170400000;
#10;x=-170390000;
#10;x=-170380000;
#10;x=-170370000;
#10;x=-170360000;
#10;x=-170350000;
#10;x=-170340000;
#10;x=-170330000;
#10;x=-170320000;
#10;x=-170310000;
#10;x=-170300000;
#10;x=-170290000;
#10;x=-170280000;
#10;x=-170270000;
#10;x=-170260000;
#10;x=-170250000;
#10;x=-170240000;
#10;x=-170230000;
#10;x=-170220000;
#10;x=-170210000;
#10;x=-170200000;
#10;x=-170190000;
#10;x=-170180000;
#10;x=-170170000;
#10;x=-170160000;
#10;x=-170150000;
#10;x=-170140000;
#10;x=-170130000;
#10;x=-170120000;
#10;x=-170110000;
#10;x=-170100000;
#10;x=-170090000;
#10;x=-170080000;
#10;x=-170070000;
#10;x=-170060000;
#10;x=-170050000;
#10;x=-170040000;
#10;x=-170030000;
#10;x=-170020000;
#10;x=-170010000;
#10;x=-170000000;
#10;x=-169990000;
#10;x=-169980000;
#10;x=-169970000;
#10;x=-169960000;
#10;x=-169950000;
#10;x=-169940000;
#10;x=-169930000;
#10;x=-169920000;
#10;x=-169910000;
#10;x=-169900000;
#10;x=-169890000;
#10;x=-169880000;
#10;x=-169870000;
#10;x=-169860000;
#10;x=-169850000;
#10;x=-169840000;
#10;x=-169830000;
#10;x=-169820000;
#10;x=-169810000;
#10;x=-169800000;
#10;x=-169790000;
#10;x=-169780000;
#10;x=-169770000;
#10;x=-169760000;
#10;x=-169750000;
#10;x=-169740000;
#10;x=-169730000;
#10;x=-169720000;
#10;x=-169710000;
#10;x=-169700000;
#10;x=-169690000;
#10;x=-169680000;
#10;x=-169670000;
#10;x=-169660000;
#10;x=-169650000;
#10;x=-169640000;
#10;x=-169630000;
#10;x=-169620000;
#10;x=-169610000;
#10;x=-169600000;
#10;x=-169590000;
#10;x=-169580000;
#10;x=-169570000;
#10;x=-169560000;
#10;x=-169550000;
#10;x=-169540000;
#10;x=-169530000;
#10;x=-169520000;
#10;x=-169510000;
#10;x=-169500000;
#10;x=-169490000;
#10;x=-169480000;
#10;x=-169470000;
#10;x=-169460000;
#10;x=-169450000;
#10;x=-169440000;
#10;x=-169430000;
#10;x=-169420000;
#10;x=-169410000;
#10;x=-169400000;
#10;x=-169390000;
#10;x=-169380000;
#10;x=-169370000;
#10;x=-169360000;
#10;x=-169350000;
#10;x=-169340000;
#10;x=-169330000;
#10;x=-169320000;
#10;x=-169310000;
#10;x=-169300000;
#10;x=-169290000;
#10;x=-169280000;
#10;x=-169270000;
#10;x=-169260000;
#10;x=-169250000;
#10;x=-169240000;
#10;x=-169230000;
#10;x=-169220000;
#10;x=-169210000;
#10;x=-169200000;
#10;x=-169190000;
#10;x=-169180000;
#10;x=-169170000;
#10;x=-169160000;
#10;x=-169150000;
#10;x=-169140000;
#10;x=-169130000;
#10;x=-169120000;
#10;x=-169110000;
#10;x=-169100000;
#10;x=-169090000;
#10;x=-169080000;
#10;x=-169070000;
#10;x=-169060000;
#10;x=-169050000;
#10;x=-169040000;
#10;x=-169030000;
#10;x=-169020000;
#10;x=-169010000;
#10;x=-169000000;
#10;x=-168990000;
#10;x=-168980000;
#10;x=-168970000;
#10;x=-168960000;
#10;x=-168950000;
#10;x=-168940000;
#10;x=-168930000;
#10;x=-168920000;
#10;x=-168910000;
#10;x=-168900000;
#10;x=-168890000;
#10;x=-168880000;
#10;x=-168870000;
#10;x=-168860000;
#10;x=-168850000;
#10;x=-168840000;
#10;x=-168830000;
#10;x=-168820000;
#10;x=-168810000;
#10;x=-168800000;
#10;x=-168790000;
#10;x=-168780000;
#10;x=-168770000;
#10;x=-168760000;
#10;x=-168750000;
#10;x=-168740000;
#10;x=-168730000;
#10;x=-168720000;
#10;x=-168710000;
#10;x=-168700000;
#10;x=-168690000;
#10;x=-168680000;
#10;x=-168670000;
#10;x=-168660000;
#10;x=-168650000;
#10;x=-168640000;
#10;x=-168630000;
#10;x=-168620000;
#10;x=-168610000;
#10;x=-168600000;
#10;x=-168590000;
#10;x=-168580000;
#10;x=-168570000;
#10;x=-168560000;
#10;x=-168550000;
#10;x=-168540000;
#10;x=-168530000;
#10;x=-168520000;
#10;x=-168510000;
#10;x=-168500000;
#10;x=-168490000;
#10;x=-168480000;
#10;x=-168470000;
#10;x=-168460000;
#10;x=-168450000;
#10;x=-168440000;
#10;x=-168430000;
#10;x=-168420000;
#10;x=-168410000;
#10;x=-168400000;
#10;x=-168390000;
#10;x=-168380000;
#10;x=-168370000;
#10;x=-168360000;
#10;x=-168350000;
#10;x=-168340000;
#10;x=-168330000;
#10;x=-168320000;
#10;x=-168310000;
#10;x=-168300000;
#10;x=-168290000;
#10;x=-168280000;
#10;x=-168270000;
#10;x=-168260000;
#10;x=-168250000;
#10;x=-168240000;
#10;x=-168230000;
#10;x=-168220000;
#10;x=-168210000;
#10;x=-168200000;
#10;x=-168190000;
#10;x=-168180000;
#10;x=-168170000;
#10;x=-168160000;
#10;x=-168150000;
#10;x=-168140000;
#10;x=-168130000;
#10;x=-168120000;
#10;x=-168110000;
#10;x=-168100000;
#10;x=-168090000;
#10;x=-168080000;
#10;x=-168070000;
#10;x=-168060000;
#10;x=-168050000;
#10;x=-168040000;
#10;x=-168030000;
#10;x=-168020000;
#10;x=-168010000;
#10;x=-168000000;
#10;x=-167990000;
#10;x=-167980000;
#10;x=-167970000;
#10;x=-167960000;
#10;x=-167950000;
#10;x=-167940000;
#10;x=-167930000;
#10;x=-167920000;
#10;x=-167910000;
#10;x=-167900000;
#10;x=-167890000;
#10;x=-167880000;
#10;x=-167870000;
#10;x=-167860000;
#10;x=-167850000;
#10;x=-167840000;
#10;x=-167830000;
#10;x=-167820000;
#10;x=-167810000;
#10;x=-167800000;
#10;x=-167790000;
#10;x=-167780000;
#10;x=-167770000;
#10;x=-167760000;
#10;x=-167750000;
#10;x=-167740000;
#10;x=-167730000;
#10;x=-167720000;
#10;x=-167710000;
#10;x=-167700000;
#10;x=-167690000;
#10;x=-167680000;
#10;x=-167670000;
#10;x=-167660000;
#10;x=-167650000;
#10;x=-167640000;
#10;x=-167630000;
#10;x=-167620000;
#10;x=-167610000;
#10;x=-167600000;
#10;x=-167590000;
#10;x=-167580000;
#10;x=-167570000;
#10;x=-167560000;
#10;x=-167550000;
#10;x=-167540000;
#10;x=-167530000;
#10;x=-167520000;
#10;x=-167510000;
#10;x=-167500000;
#10;x=-167490000;
#10;x=-167480000;
#10;x=-167470000;
#10;x=-167460000;
#10;x=-167450000;
#10;x=-167440000;
#10;x=-167430000;
#10;x=-167420000;
#10;x=-167410000;
#10;x=-167400000;
#10;x=-167390000;
#10;x=-167380000;
#10;x=-167370000;
#10;x=-167360000;
#10;x=-167350000;
#10;x=-167340000;
#10;x=-167330000;
#10;x=-167320000;
#10;x=-167310000;
#10;x=-167300000;
#10;x=-167290000;
#10;x=-167280000;
#10;x=-167270000;
#10;x=-167260000;
#10;x=-167250000;
#10;x=-167240000;
#10;x=-167230000;
#10;x=-167220000;
#10;x=-167210000;
#10;x=-167200000;
#10;x=-167190000;
#10;x=-167180000;
#10;x=-167170000;
#10;x=-167160000;
#10;x=-167150000;
#10;x=-167140000;
#10;x=-167130000;
#10;x=-167120000;
#10;x=-167110000;
#10;x=-167100000;
#10;x=-167090000;
#10;x=-167080000;
#10;x=-167070000;
#10;x=-167060000;
#10;x=-167050000;
#10;x=-167040000;
#10;x=-167030000;
#10;x=-167020000;
#10;x=-167010000;
#10;x=-167000000;
#10;x=-166990000;
#10;x=-166980000;
#10;x=-166970000;
#10;x=-166960000;
#10;x=-166950000;
#10;x=-166940000;
#10;x=-166930000;
#10;x=-166920000;
#10;x=-166910000;
#10;x=-166900000;
#10;x=-166890000;
#10;x=-166880000;
#10;x=-166870000;
#10;x=-166860000;
#10;x=-166850000;
#10;x=-166840000;
#10;x=-166830000;
#10;x=-166820000;
#10;x=-166810000;
#10;x=-166800000;
#10;x=-166790000;
#10;x=-166780000;
#10;x=-166770000;
#10;x=-166760000;
#10;x=-166750000;
#10;x=-166740000;
#10;x=-166730000;
#10;x=-166720000;
#10;x=-166710000;
#10;x=-166700000;
#10;x=-166690000;
#10;x=-166680000;
#10;x=-166670000;
#10;x=-166660000;
#10;x=-166650000;
#10;x=-166640000;
#10;x=-166630000;
#10;x=-166620000;
#10;x=-166610000;
#10;x=-166600000;
#10;x=-166590000;
#10;x=-166580000;
#10;x=-166570000;
#10;x=-166560000;
#10;x=-166550000;
#10;x=-166540000;
#10;x=-166530000;
#10;x=-166520000;
#10;x=-166510000;
#10;x=-166500000;
#10;x=-166490000;
#10;x=-166480000;
#10;x=-166470000;
#10;x=-166460000;
#10;x=-166450000;
#10;x=-166440000;
#10;x=-166430000;
#10;x=-166420000;
#10;x=-166410000;
#10;x=-166400000;
#10;x=-166390000;
#10;x=-166380000;
#10;x=-166370000;
#10;x=-166360000;
#10;x=-166350000;
#10;x=-166340000;
#10;x=-166330000;
#10;x=-166320000;
#10;x=-166310000;
#10;x=-166300000;
#10;x=-166290000;
#10;x=-166280000;
#10;x=-166270000;
#10;x=-166260000;
#10;x=-166250000;
#10;x=-166240000;
#10;x=-166230000;
#10;x=-166220000;
#10;x=-166210000;
#10;x=-166200000;
#10;x=-166190000;
#10;x=-166180000;
#10;x=-166170000;
#10;x=-166160000;
#10;x=-166150000;
#10;x=-166140000;
#10;x=-166130000;
#10;x=-166120000;
#10;x=-166110000;
#10;x=-166100000;
#10;x=-166090000;
#10;x=-166080000;
#10;x=-166070000;
#10;x=-166060000;
#10;x=-166050000;
#10;x=-166040000;
#10;x=-166030000;
#10;x=-166020000;
#10;x=-166010000;
#10;x=-166000000;
#10;x=-165990000;
#10;x=-165980000;
#10;x=-165970000;
#10;x=-165960000;
#10;x=-165950000;
#10;x=-165940000;
#10;x=-165930000;
#10;x=-165920000;
#10;x=-165910000;
#10;x=-165900000;
#10;x=-165890000;
#10;x=-165880000;
#10;x=-165870000;
#10;x=-165860000;
#10;x=-165850000;
#10;x=-165840000;
#10;x=-165830000;
#10;x=-165820000;
#10;x=-165810000;
#10;x=-165800000;
#10;x=-165790000;
#10;x=-165780000;
#10;x=-165770000;
#10;x=-165760000;
#10;x=-165750000;
#10;x=-165740000;
#10;x=-165730000;
#10;x=-165720000;
#10;x=-165710000;
#10;x=-165700000;
#10;x=-165690000;
#10;x=-165680000;
#10;x=-165670000;
#10;x=-165660000;
#10;x=-165650000;
#10;x=-165640000;
#10;x=-165630000;
#10;x=-165620000;
#10;x=-165610000;
#10;x=-165600000;
#10;x=-165590000;
#10;x=-165580000;
#10;x=-165570000;
#10;x=-165560000;
#10;x=-165550000;
#10;x=-165540000;
#10;x=-165530000;
#10;x=-165520000;
#10;x=-165510000;
#10;x=-165500000;
#10;x=-165490000;
#10;x=-165480000;
#10;x=-165470000;
#10;x=-165460000;
#10;x=-165450000;
#10;x=-165440000;
#10;x=-165430000;
#10;x=-165420000;
#10;x=-165410000;
#10;x=-165400000;
#10;x=-165390000;
#10;x=-165380000;
#10;x=-165370000;
#10;x=-165360000;
#10;x=-165350000;
#10;x=-165340000;
#10;x=-165330000;
#10;x=-165320000;
#10;x=-165310000;
#10;x=-165300000;
#10;x=-165290000;
#10;x=-165280000;
#10;x=-165270000;
#10;x=-165260000;
#10;x=-165250000;
#10;x=-165240000;
#10;x=-165230000;
#10;x=-165220000;
#10;x=-165210000;
#10;x=-165200000;
#10;x=-165190000;
#10;x=-165180000;
#10;x=-165170000;
#10;x=-165160000;
#10;x=-165150000;
#10;x=-165140000;
#10;x=-165130000;
#10;x=-165120000;
#10;x=-165110000;
#10;x=-165100000;
#10;x=-165090000;
#10;x=-165080000;
#10;x=-165070000;
#10;x=-165060000;
#10;x=-165050000;
#10;x=-165040000;
#10;x=-165030000;
#10;x=-165020000;
#10;x=-165010000;
#10;x=-165000000;
#10;x=-164990000;
#10;x=-164980000;
#10;x=-164970000;
#10;x=-164960000;
#10;x=-164950000;
#10;x=-164940000;
#10;x=-164930000;
#10;x=-164920000;
#10;x=-164910000;
#10;x=-164900000;
#10;x=-164890000;
#10;x=-164880000;
#10;x=-164870000;
#10;x=-164860000;
#10;x=-164850000;
#10;x=-164840000;
#10;x=-164830000;
#10;x=-164820000;
#10;x=-164810000;
#10;x=-164800000;
#10;x=-164790000;
#10;x=-164780000;
#10;x=-164770000;
#10;x=-164760000;
#10;x=-164750000;
#10;x=-164740000;
#10;x=-164730000;
#10;x=-164720000;
#10;x=-164710000;
#10;x=-164700000;
#10;x=-164690000;
#10;x=-164680000;
#10;x=-164670000;
#10;x=-164660000;
#10;x=-164650000;
#10;x=-164640000;
#10;x=-164630000;
#10;x=-164620000;
#10;x=-164610000;
#10;x=-164600000;
#10;x=-164590000;
#10;x=-164580000;
#10;x=-164570000;
#10;x=-164560000;
#10;x=-164550000;
#10;x=-164540000;
#10;x=-164530000;
#10;x=-164520000;
#10;x=-164510000;
#10;x=-164500000;
#10;x=-164490000;
#10;x=-164480000;
#10;x=-164470000;
#10;x=-164460000;
#10;x=-164450000;
#10;x=-164440000;
#10;x=-164430000;
#10;x=-164420000;
#10;x=-164410000;
#10;x=-164400000;
#10;x=-164390000;
#10;x=-164380000;
#10;x=-164370000;
#10;x=-164360000;
#10;x=-164350000;
#10;x=-164340000;
#10;x=-164330000;
#10;x=-164320000;
#10;x=-164310000;
#10;x=-164300000;
#10;x=-164290000;
#10;x=-164280000;
#10;x=-164270000;
#10;x=-164260000;
#10;x=-164250000;
#10;x=-164240000;
#10;x=-164230000;
#10;x=-164220000;
#10;x=-164210000;
#10;x=-164200000;
#10;x=-164190000;
#10;x=-164180000;
#10;x=-164170000;
#10;x=-164160000;
#10;x=-164150000;
#10;x=-164140000;
#10;x=-164130000;
#10;x=-164120000;
#10;x=-164110000;
#10;x=-164100000;
#10;x=-164090000;
#10;x=-164080000;
#10;x=-164070000;
#10;x=-164060000;
#10;x=-164050000;
#10;x=-164040000;
#10;x=-164030000;
#10;x=-164020000;
#10;x=-164010000;
#10;x=-164000000;
#10;x=-163990000;
#10;x=-163980000;
#10;x=-163970000;
#10;x=-163960000;
#10;x=-163950000;
#10;x=-163940000;
#10;x=-163930000;
#10;x=-163920000;
#10;x=-163910000;
#10;x=-163900000;
#10;x=-163890000;
#10;x=-163880000;
#10;x=-163870000;
#10;x=-163860000;
#10;x=-163850000;
#10;x=-163840000;
#10;x=-163830000;
#10;x=-163820000;
#10;x=-163810000;
#10;x=-163800000;
#10;x=-163790000;
#10;x=-163780000;
#10;x=-163770000;
#10;x=-163760000;
#10;x=-163750000;
#10;x=-163740000;
#10;x=-163730000;
#10;x=-163720000;
#10;x=-163710000;
#10;x=-163700000;
#10;x=-163690000;
#10;x=-163680000;
#10;x=-163670000;
#10;x=-163660000;
#10;x=-163650000;
#10;x=-163640000;
#10;x=-163630000;
#10;x=-163620000;
#10;x=-163610000;
#10;x=-163600000;
#10;x=-163590000;
#10;x=-163580000;
#10;x=-163570000;
#10;x=-163560000;
#10;x=-163550000;
#10;x=-163540000;
#10;x=-163530000;
#10;x=-163520000;
#10;x=-163510000;
#10;x=-163500000;
#10;x=-163490000;
#10;x=-163480000;
#10;x=-163470000;
#10;x=-163460000;
#10;x=-163450000;
#10;x=-163440000;
#10;x=-163430000;
#10;x=-163420000;
#10;x=-163410000;
#10;x=-163400000;
#10;x=-163390000;
#10;x=-163380000;
#10;x=-163370000;
#10;x=-163360000;
#10;x=-163350000;
#10;x=-163340000;
#10;x=-163330000;
#10;x=-163320000;
#10;x=-163310000;
#10;x=-163300000;
#10;x=-163290000;
#10;x=-163280000;
#10;x=-163270000;
#10;x=-163260000;
#10;x=-163250000;
#10;x=-163240000;
#10;x=-163230000;
#10;x=-163220000;
#10;x=-163210000;
#10;x=-163200000;
#10;x=-163190000;
#10;x=-163180000;
#10;x=-163170000;
#10;x=-163160000;
#10;x=-163150000;
#10;x=-163140000;
#10;x=-163130000;
#10;x=-163120000;
#10;x=-163110000;
#10;x=-163100000;
#10;x=-163090000;
#10;x=-163080000;
#10;x=-163070000;
#10;x=-163060000;
#10;x=-163050000;
#10;x=-163040000;
#10;x=-163030000;
#10;x=-163020000;
#10;x=-163010000;
#10;x=-163000000;
#10;x=-162990000;
#10;x=-162980000;
#10;x=-162970000;
#10;x=-162960000;
#10;x=-162950000;
#10;x=-162940000;
#10;x=-162930000;
#10;x=-162920000;
#10;x=-162910000;
#10;x=-162900000;
#10;x=-162890000;
#10;x=-162880000;
#10;x=-162870000;
#10;x=-162860000;
#10;x=-162850000;
#10;x=-162840000;
#10;x=-162830000;
#10;x=-162820000;
#10;x=-162810000;
#10;x=-162800000;
#10;x=-162790000;
#10;x=-162780000;
#10;x=-162770000;
#10;x=-162760000;
#10;x=-162750000;
#10;x=-162740000;
#10;x=-162730000;
#10;x=-162720000;
#10;x=-162710000;
#10;x=-162700000;
#10;x=-162690000;
#10;x=-162680000;
#10;x=-162670000;
#10;x=-162660000;
#10;x=-162650000;
#10;x=-162640000;
#10;x=-162630000;
#10;x=-162620000;
#10;x=-162610000;
#10;x=-162600000;
#10;x=-162590000;
#10;x=-162580000;
#10;x=-162570000;
#10;x=-162560000;
#10;x=-162550000;
#10;x=-162540000;
#10;x=-162530000;
#10;x=-162520000;
#10;x=-162510000;
#10;x=-162500000;
#10;x=-162490000;
#10;x=-162480000;
#10;x=-162470000;
#10;x=-162460000;
#10;x=-162450000;
#10;x=-162440000;
#10;x=-162430000;
#10;x=-162420000;
#10;x=-162410000;
#10;x=-162400000;
#10;x=-162390000;
#10;x=-162380000;
#10;x=-162370000;
#10;x=-162360000;
#10;x=-162350000;
#10;x=-162340000;
#10;x=-162330000;
#10;x=-162320000;
#10;x=-162310000;
#10;x=-162300000;
#10;x=-162290000;
#10;x=-162280000;
#10;x=-162270000;
#10;x=-162260000;
#10;x=-162250000;
#10;x=-162240000;
#10;x=-162230000;
#10;x=-162220000;
#10;x=-162210000;
#10;x=-162200000;
#10;x=-162190000;
#10;x=-162180000;
#10;x=-162170000;
#10;x=-162160000;
#10;x=-162150000;
#10;x=-162140000;
#10;x=-162130000;
#10;x=-162120000;
#10;x=-162110000;
#10;x=-162100000;
#10;x=-162090000;
#10;x=-162080000;
#10;x=-162070000;
#10;x=-162060000;
#10;x=-162050000;
#10;x=-162040000;
#10;x=-162030000;
#10;x=-162020000;
#10;x=-162010000;
#10;x=-162000000;
#10;x=-161990000;
#10;x=-161980000;
#10;x=-161970000;
#10;x=-161960000;
#10;x=-161950000;
#10;x=-161940000;
#10;x=-161930000;
#10;x=-161920000;
#10;x=-161910000;
#10;x=-161900000;
#10;x=-161890000;
#10;x=-161880000;
#10;x=-161870000;
#10;x=-161860000;
#10;x=-161850000;
#10;x=-161840000;
#10;x=-161830000;
#10;x=-161820000;
#10;x=-161810000;
#10;x=-161800000;
#10;x=-161790000;
#10;x=-161780000;
#10;x=-161770000;
#10;x=-161760000;
#10;x=-161750000;
#10;x=-161740000;
#10;x=-161730000;
#10;x=-161720000;
#10;x=-161710000;
#10;x=-161700000;
#10;x=-161690000;
#10;x=-161680000;
#10;x=-161670000;
#10;x=-161660000;
#10;x=-161650000;
#10;x=-161640000;
#10;x=-161630000;
#10;x=-161620000;
#10;x=-161610000;
#10;x=-161600000;
#10;x=-161590000;
#10;x=-161580000;
#10;x=-161570000;
#10;x=-161560000;
#10;x=-161550000;
#10;x=-161540000;
#10;x=-161530000;
#10;x=-161520000;
#10;x=-161510000;
#10;x=-161500000;
#10;x=-161490000;
#10;x=-161480000;
#10;x=-161470000;
#10;x=-161460000;
#10;x=-161450000;
#10;x=-161440000;
#10;x=-161430000;
#10;x=-161420000;
#10;x=-161410000;
#10;x=-161400000;
#10;x=-161390000;
#10;x=-161380000;
#10;x=-161370000;
#10;x=-161360000;
#10;x=-161350000;
#10;x=-161340000;
#10;x=-161330000;
#10;x=-161320000;
#10;x=-161310000;
#10;x=-161300000;
#10;x=-161290000;
#10;x=-161280000;
#10;x=-161270000;
#10;x=-161260000;
#10;x=-161250000;
#10;x=-161240000;
#10;x=-161230000;
#10;x=-161220000;
#10;x=-161210000;
#10;x=-161200000;
#10;x=-161190000;
#10;x=-161180000;
#10;x=-161170000;
#10;x=-161160000;
#10;x=-161150000;
#10;x=-161140000;
#10;x=-161130000;
#10;x=-161120000;
#10;x=-161110000;
#10;x=-161100000;
#10;x=-161090000;
#10;x=-161080000;
#10;x=-161070000;
#10;x=-161060000;
#10;x=-161050000;
#10;x=-161040000;
#10;x=-161030000;
#10;x=-161020000;
#10;x=-161010000;
#10;x=-161000000;
#10;x=-160990000;
#10;x=-160980000;
#10;x=-160970000;
#10;x=-160960000;
#10;x=-160950000;
#10;x=-160940000;
#10;x=-160930000;
#10;x=-160920000;
#10;x=-160910000;
#10;x=-160900000;
#10;x=-160890000;
#10;x=-160880000;
#10;x=-160870000;
#10;x=-160860000;
#10;x=-160850000;
#10;x=-160840000;
#10;x=-160830000;
#10;x=-160820000;
#10;x=-160810000;
#10;x=-160800000;
#10;x=-160790000;
#10;x=-160780000;
#10;x=-160770000;
#10;x=-160760000;
#10;x=-160750000;
#10;x=-160740000;
#10;x=-160730000;
#10;x=-160720000;
#10;x=-160710000;
#10;x=-160700000;
#10;x=-160690000;
#10;x=-160680000;
#10;x=-160670000;
#10;x=-160660000;
#10;x=-160650000;
#10;x=-160640000;
#10;x=-160630000;
#10;x=-160620000;
#10;x=-160610000;
#10;x=-160600000;
#10;x=-160590000;
#10;x=-160580000;
#10;x=-160570000;
#10;x=-160560000;
#10;x=-160550000;
#10;x=-160540000;
#10;x=-160530000;
#10;x=-160520000;
#10;x=-160510000;
#10;x=-160500000;
#10;x=-160490000;
#10;x=-160480000;
#10;x=-160470000;
#10;x=-160460000;
#10;x=-160450000;
#10;x=-160440000;
#10;x=-160430000;
#10;x=-160420000;
#10;x=-160410000;
#10;x=-160400000;
#10;x=-160390000;
#10;x=-160380000;
#10;x=-160370000;
#10;x=-160360000;
#10;x=-160350000;
#10;x=-160340000;
#10;x=-160330000;
#10;x=-160320000;
#10;x=-160310000;
#10;x=-160300000;
#10;x=-160290000;
#10;x=-160280000;
#10;x=-160270000;
#10;x=-160260000;
#10;x=-160250000;
#10;x=-160240000;
#10;x=-160230000;
#10;x=-160220000;
#10;x=-160210000;
#10;x=-160200000;
#10;x=-160190000;
#10;x=-160180000;
#10;x=-160170000;
#10;x=-160160000;
#10;x=-160150000;
#10;x=-160140000;
#10;x=-160130000;
#10;x=-160120000;
#10;x=-160110000;
#10;x=-160100000;
#10;x=-160090000;
#10;x=-160080000;
#10;x=-160070000;
#10;x=-160060000;
#10;x=-160050000;
#10;x=-160040000;
#10;x=-160030000;
#10;x=-160020000;
#10;x=-160010000;
#10;x=-160000000;
#10;x=-159990000;
#10;x=-159980000;
#10;x=-159970000;
#10;x=-159960000;
#10;x=-159950000;
#10;x=-159940000;
#10;x=-159930000;
#10;x=-159920000;
#10;x=-159910000;
#10;x=-159900000;
#10;x=-159890000;
#10;x=-159880000;
#10;x=-159870000;
#10;x=-159860000;
#10;x=-159850000;
#10;x=-159840000;
#10;x=-159830000;
#10;x=-159820000;
#10;x=-159810000;
#10;x=-159800000;
#10;x=-159790000;
#10;x=-159780000;
#10;x=-159770000;
#10;x=-159760000;
#10;x=-159750000;
#10;x=-159740000;
#10;x=-159730000;
#10;x=-159720000;
#10;x=-159710000;
#10;x=-159700000;
#10;x=-159690000;
#10;x=-159680000;
#10;x=-159670000;
#10;x=-159660000;
#10;x=-159650000;
#10;x=-159640000;
#10;x=-159630000;
#10;x=-159620000;
#10;x=-159610000;
#10;x=-159600000;
#10;x=-159590000;
#10;x=-159580000;
#10;x=-159570000;
#10;x=-159560000;
#10;x=-159550000;
#10;x=-159540000;
#10;x=-159530000;
#10;x=-159520000;
#10;x=-159510000;
#10;x=-159500000;
#10;x=-159490000;
#10;x=-159480000;
#10;x=-159470000;
#10;x=-159460000;
#10;x=-159450000;
#10;x=-159440000;
#10;x=-159430000;
#10;x=-159420000;
#10;x=-159410000;
#10;x=-159400000;
#10;x=-159390000;
#10;x=-159380000;
#10;x=-159370000;
#10;x=-159360000;
#10;x=-159350000;
#10;x=-159340000;
#10;x=-159330000;
#10;x=-159320000;
#10;x=-159310000;
#10;x=-159300000;
#10;x=-159290000;
#10;x=-159280000;
#10;x=-159270000;
#10;x=-159260000;
#10;x=-159250000;
#10;x=-159240000;
#10;x=-159230000;
#10;x=-159220000;
#10;x=-159210000;
#10;x=-159200000;
#10;x=-159190000;
#10;x=-159180000;
#10;x=-159170000;
#10;x=-159160000;
#10;x=-159150000;
#10;x=-159140000;
#10;x=-159130000;
#10;x=-159120000;
#10;x=-159110000;
#10;x=-159100000;
#10;x=-159090000;
#10;x=-159080000;
#10;x=-159070000;
#10;x=-159060000;
#10;x=-159050000;
#10;x=-159040000;
#10;x=-159030000;
#10;x=-159020000;
#10;x=-159010000;
#10;x=-159000000;
#10;x=-158990000;
#10;x=-158980000;
#10;x=-158970000;
#10;x=-158960000;
#10;x=-158950000;
#10;x=-158940000;
#10;x=-158930000;
#10;x=-158920000;
#10;x=-158910000;
#10;x=-158900000;
#10;x=-158890000;
#10;x=-158880000;
#10;x=-158870000;
#10;x=-158860000;
#10;x=-158850000;
#10;x=-158840000;
#10;x=-158830000;
#10;x=-158820000;
#10;x=-158810000;
#10;x=-158800000;
#10;x=-158790000;
#10;x=-158780000;
#10;x=-158770000;
#10;x=-158760000;
#10;x=-158750000;
#10;x=-158740000;
#10;x=-158730000;
#10;x=-158720000;
#10;x=-158710000;
#10;x=-158700000;
#10;x=-158690000;
#10;x=-158680000;
#10;x=-158670000;
#10;x=-158660000;
#10;x=-158650000;
#10;x=-158640000;
#10;x=-158630000;
#10;x=-158620000;
#10;x=-158610000;
#10;x=-158600000;
#10;x=-158590000;
#10;x=-158580000;
#10;x=-158570000;
#10;x=-158560000;
#10;x=-158550000;
#10;x=-158540000;
#10;x=-158530000;
#10;x=-158520000;
#10;x=-158510000;
#10;x=-158500000;
#10;x=-158490000;
#10;x=-158480000;
#10;x=-158470000;
#10;x=-158460000;
#10;x=-158450000;
#10;x=-158440000;
#10;x=-158430000;
#10;x=-158420000;
#10;x=-158410000;
#10;x=-158400000;
#10;x=-158390000;
#10;x=-158380000;
#10;x=-158370000;
#10;x=-158360000;
#10;x=-158350000;
#10;x=-158340000;
#10;x=-158330000;
#10;x=-158320000;
#10;x=-158310000;
#10;x=-158300000;
#10;x=-158290000;
#10;x=-158280000;
#10;x=-158270000;
#10;x=-158260000;
#10;x=-158250000;
#10;x=-158240000;
#10;x=-158230000;
#10;x=-158220000;
#10;x=-158210000;
#10;x=-158200000;
#10;x=-158190000;
#10;x=-158180000;
#10;x=-158170000;
#10;x=-158160000;
#10;x=-158150000;
#10;x=-158140000;
#10;x=-158130000;
#10;x=-158120000;
#10;x=-158110000;
#10;x=-158100000;
#10;x=-158090000;
#10;x=-158080000;
#10;x=-158070000;
#10;x=-158060000;
#10;x=-158050000;
#10;x=-158040000;
#10;x=-158030000;
#10;x=-158020000;
#10;x=-158010000;
#10;x=-158000000;
#10;x=-157990000;
#10;x=-157980000;
#10;x=-157970000;
#10;x=-157960000;
#10;x=-157950000;
#10;x=-157940000;
#10;x=-157930000;
#10;x=-157920000;
#10;x=-157910000;
#10;x=-157900000;
#10;x=-157890000;
#10;x=-157880000;
#10;x=-157870000;
#10;x=-157860000;
#10;x=-157850000;
#10;x=-157840000;
#10;x=-157830000;
#10;x=-157820000;
#10;x=-157810000;
#10;x=-157800000;
#10;x=-157790000;
#10;x=-157780000;
#10;x=-157770000;
#10;x=-157760000;
#10;x=-157750000;
#10;x=-157740000;
#10;x=-157730000;
#10;x=-157720000;
#10;x=-157710000;
#10;x=-157700000;
#10;x=-157690000;
#10;x=-157680000;
#10;x=-157670000;
#10;x=-157660000;
#10;x=-157650000;
#10;x=-157640000;
#10;x=-157630000;
#10;x=-157620000;
#10;x=-157610000;
#10;x=-157600000;
#10;x=-157590000;
#10;x=-157580000;
#10;x=-157570000;
#10;x=-157560000;
#10;x=-157550000;
#10;x=-157540000;
#10;x=-157530000;
#10;x=-157520000;
#10;x=-157510000;
#10;x=-157500000;
#10;x=-157490000;
#10;x=-157480000;
#10;x=-157470000;
#10;x=-157460000;
#10;x=-157450000;
#10;x=-157440000;
#10;x=-157430000;
#10;x=-157420000;
#10;x=-157410000;
#10;x=-157400000;
#10;x=-157390000;
#10;x=-157380000;
#10;x=-157370000;
#10;x=-157360000;
#10;x=-157350000;
#10;x=-157340000;
#10;x=-157330000;
#10;x=-157320000;
#10;x=-157310000;
#10;x=-157300000;
#10;x=-157290000;
#10;x=-157280000;
#10;x=-157270000;
#10;x=-157260000;
#10;x=-157250000;
#10;x=-157240000;
#10;x=-157230000;
#10;x=-157220000;
#10;x=-157210000;
#10;x=-157200000;
#10;x=-157190000;
#10;x=-157180000;
#10;x=-157170000;
#10;x=-157160000;
#10;x=-157150000;
#10;x=-157140000;
#10;x=-157130000;
#10;x=-157120000;
#10;x=-157110000;
#10;x=-157100000;
#10;x=-157090000;
#10;x=-157080000;
#10;x=-157070000;
#10;x=-157060000;
#10;x=-157050000;
#10;x=-157040000;
#10;x=-157030000;
#10;x=-157020000;
#10;x=-157010000;
#10;x=-157000000;
#10;x=-156990000;
#10;x=-156980000;
#10;x=-156970000;
#10;x=-156960000;
#10;x=-156950000;
#10;x=-156940000;
#10;x=-156930000;
#10;x=-156920000;
#10;x=-156910000;
#10;x=-156900000;
#10;x=-156890000;
#10;x=-156880000;
#10;x=-156870000;
#10;x=-156860000;
#10;x=-156850000;
#10;x=-156840000;
#10;x=-156830000;
#10;x=-156820000;
#10;x=-156810000;
#10;x=-156800000;
#10;x=-156790000;
#10;x=-156780000;
#10;x=-156770000;
#10;x=-156760000;
#10;x=-156750000;
#10;x=-156740000;
#10;x=-156730000;
#10;x=-156720000;
#10;x=-156710000;
#10;x=-156700000;
#10;x=-156690000;
#10;x=-156680000;
#10;x=-156670000;
#10;x=-156660000;
#10;x=-156650000;
#10;x=-156640000;
#10;x=-156630000;
#10;x=-156620000;
#10;x=-156610000;
#10;x=-156600000;
#10;x=-156590000;
#10;x=-156580000;
#10;x=-156570000;
#10;x=-156560000;
#10;x=-156550000;
#10;x=-156540000;
#10;x=-156530000;
#10;x=-156520000;
#10;x=-156510000;
#10;x=-156500000;
#10;x=-156490000;
#10;x=-156480000;
#10;x=-156470000;
#10;x=-156460000;
#10;x=-156450000;
#10;x=-156440000;
#10;x=-156430000;
#10;x=-156420000;
#10;x=-156410000;
#10;x=-156400000;
#10;x=-156390000;
#10;x=-156380000;
#10;x=-156370000;
#10;x=-156360000;
#10;x=-156350000;
#10;x=-156340000;
#10;x=-156330000;
#10;x=-156320000;
#10;x=-156310000;
#10;x=-156300000;
#10;x=-156290000;
#10;x=-156280000;
#10;x=-156270000;
#10;x=-156260000;
#10;x=-156250000;
#10;x=-156240000;
#10;x=-156230000;
#10;x=-156220000;
#10;x=-156210000;
#10;x=-156200000;
#10;x=-156190000;
#10;x=-156180000;
#10;x=-156170000;
#10;x=-156160000;
#10;x=-156150000;
#10;x=-156140000;
#10;x=-156130000;
#10;x=-156120000;
#10;x=-156110000;
#10;x=-156100000;
#10;x=-156090000;
#10;x=-156080000;
#10;x=-156070000;
#10;x=-156060000;
#10;x=-156050000;
#10;x=-156040000;
#10;x=-156030000;
#10;x=-156020000;
#10;x=-156010000;
#10;x=-156000000;
#10;x=-155990000;
#10;x=-155980000;
#10;x=-155970000;
#10;x=-155960000;
#10;x=-155950000;
#10;x=-155940000;
#10;x=-155930000;
#10;x=-155920000;
#10;x=-155910000;
#10;x=-155900000;
#10;x=-155890000;
#10;x=-155880000;
#10;x=-155870000;
#10;x=-155860000;
#10;x=-155850000;
#10;x=-155840000;
#10;x=-155830000;
#10;x=-155820000;
#10;x=-155810000;
#10;x=-155800000;
#10;x=-155790000;
#10;x=-155780000;
#10;x=-155770000;
#10;x=-155760000;
#10;x=-155750000;
#10;x=-155740000;
#10;x=-155730000;
#10;x=-155720000;
#10;x=-155710000;
#10;x=-155700000;
#10;x=-155690000;
#10;x=-155680000;
#10;x=-155670000;
#10;x=-155660000;
#10;x=-155650000;
#10;x=-155640000;
#10;x=-155630000;
#10;x=-155620000;
#10;x=-155610000;
#10;x=-155600000;
#10;x=-155590000;
#10;x=-155580000;
#10;x=-155570000;
#10;x=-155560000;
#10;x=-155550000;
#10;x=-155540000;
#10;x=-155530000;
#10;x=-155520000;
#10;x=-155510000;
#10;x=-155500000;
#10;x=-155490000;
#10;x=-155480000;
#10;x=-155470000;
#10;x=-155460000;
#10;x=-155450000;
#10;x=-155440000;
#10;x=-155430000;
#10;x=-155420000;
#10;x=-155410000;
#10;x=-155400000;
#10;x=-155390000;
#10;x=-155380000;
#10;x=-155370000;
#10;x=-155360000;
#10;x=-155350000;
#10;x=-155340000;
#10;x=-155330000;
#10;x=-155320000;
#10;x=-155310000;
#10;x=-155300000;
#10;x=-155290000;
#10;x=-155280000;
#10;x=-155270000;
#10;x=-155260000;
#10;x=-155250000;
#10;x=-155240000;
#10;x=-155230000;
#10;x=-155220000;
#10;x=-155210000;
#10;x=-155200000;
#10;x=-155190000;
#10;x=-155180000;
#10;x=-155170000;
#10;x=-155160000;
#10;x=-155150000;
#10;x=-155140000;
#10;x=-155130000;
#10;x=-155120000;
#10;x=-155110000;
#10;x=-155100000;
#10;x=-155090000;
#10;x=-155080000;
#10;x=-155070000;
#10;x=-155060000;
#10;x=-155050000;
#10;x=-155040000;
#10;x=-155030000;
#10;x=-155020000;
#10;x=-155010000;
#10;x=-155000000;
#10;x=-154990000;
#10;x=-154980000;
#10;x=-154970000;
#10;x=-154960000;
#10;x=-154950000;
#10;x=-154940000;
#10;x=-154930000;
#10;x=-154920000;
#10;x=-154910000;
#10;x=-154900000;
#10;x=-154890000;
#10;x=-154880000;
#10;x=-154870000;
#10;x=-154860000;
#10;x=-154850000;
#10;x=-154840000;
#10;x=-154830000;
#10;x=-154820000;
#10;x=-154810000;
#10;x=-154800000;
#10;x=-154790000;
#10;x=-154780000;
#10;x=-154770000;
#10;x=-154760000;
#10;x=-154750000;
#10;x=-154740000;
#10;x=-154730000;
#10;x=-154720000;
#10;x=-154710000;
#10;x=-154700000;
#10;x=-154690000;
#10;x=-154680000;
#10;x=-154670000;
#10;x=-154660000;
#10;x=-154650000;
#10;x=-154640000;
#10;x=-154630000;
#10;x=-154620000;
#10;x=-154610000;
#10;x=-154600000;
#10;x=-154590000;
#10;x=-154580000;
#10;x=-154570000;
#10;x=-154560000;
#10;x=-154550000;
#10;x=-154540000;
#10;x=-154530000;
#10;x=-154520000;
#10;x=-154510000;
#10;x=-154500000;
#10;x=-154490000;
#10;x=-154480000;
#10;x=-154470000;
#10;x=-154460000;
#10;x=-154450000;
#10;x=-154440000;
#10;x=-154430000;
#10;x=-154420000;
#10;x=-154410000;
#10;x=-154400000;
#10;x=-154390000;
#10;x=-154380000;
#10;x=-154370000;
#10;x=-154360000;
#10;x=-154350000;
#10;x=-154340000;
#10;x=-154330000;
#10;x=-154320000;
#10;x=-154310000;
#10;x=-154300000;
#10;x=-154290000;
#10;x=-154280000;
#10;x=-154270000;
#10;x=-154260000;
#10;x=-154250000;
#10;x=-154240000;
#10;x=-154230000;
#10;x=-154220000;
#10;x=-154210000;
#10;x=-154200000;
#10;x=-154190000;
#10;x=-154180000;
#10;x=-154170000;
#10;x=-154160000;
#10;x=-154150000;
#10;x=-154140000;
#10;x=-154130000;
#10;x=-154120000;
#10;x=-154110000;
#10;x=-154100000;
#10;x=-154090000;
#10;x=-154080000;
#10;x=-154070000;
#10;x=-154060000;
#10;x=-154050000;
#10;x=-154040000;
#10;x=-154030000;
#10;x=-154020000;
#10;x=-154010000;
#10;x=-154000000;
#10;x=-153990000;
#10;x=-153980000;
#10;x=-153970000;
#10;x=-153960000;
#10;x=-153950000;
#10;x=-153940000;
#10;x=-153930000;
#10;x=-153920000;
#10;x=-153910000;
#10;x=-153900000;
#10;x=-153890000;
#10;x=-153880000;
#10;x=-153870000;
#10;x=-153860000;
#10;x=-153850000;
#10;x=-153840000;
#10;x=-153830000;
#10;x=-153820000;
#10;x=-153810000;
#10;x=-153800000;
#10;x=-153790000;
#10;x=-153780000;
#10;x=-153770000;
#10;x=-153760000;
#10;x=-153750000;
#10;x=-153740000;
#10;x=-153730000;
#10;x=-153720000;
#10;x=-153710000;
#10;x=-153700000;
#10;x=-153690000;
#10;x=-153680000;
#10;x=-153670000;
#10;x=-153660000;
#10;x=-153650000;
#10;x=-153640000;
#10;x=-153630000;
#10;x=-153620000;
#10;x=-153610000;
#10;x=-153600000;
#10;x=-153590000;
#10;x=-153580000;
#10;x=-153570000;
#10;x=-153560000;
#10;x=-153550000;
#10;x=-153540000;
#10;x=-153530000;
#10;x=-153520000;
#10;x=-153510000;
#10;x=-153500000;
#10;x=-153490000;
#10;x=-153480000;
#10;x=-153470000;
#10;x=-153460000;
#10;x=-153450000;
#10;x=-153440000;
#10;x=-153430000;
#10;x=-153420000;
#10;x=-153410000;
#10;x=-153400000;
#10;x=-153390000;
#10;x=-153380000;
#10;x=-153370000;
#10;x=-153360000;
#10;x=-153350000;
#10;x=-153340000;
#10;x=-153330000;
#10;x=-153320000;
#10;x=-153310000;
#10;x=-153300000;
#10;x=-153290000;
#10;x=-153280000;
#10;x=-153270000;
#10;x=-153260000;
#10;x=-153250000;
#10;x=-153240000;
#10;x=-153230000;
#10;x=-153220000;
#10;x=-153210000;
#10;x=-153200000;
#10;x=-153190000;
#10;x=-153180000;
#10;x=-153170000;
#10;x=-153160000;
#10;x=-153150000;
#10;x=-153140000;
#10;x=-153130000;
#10;x=-153120000;
#10;x=-153110000;
#10;x=-153100000;
#10;x=-153090000;
#10;x=-153080000;
#10;x=-153070000;
#10;x=-153060000;
#10;x=-153050000;
#10;x=-153040000;
#10;x=-153030000;
#10;x=-153020000;
#10;x=-153010000;
#10;x=-153000000;
#10;x=-152990000;
#10;x=-152980000;
#10;x=-152970000;
#10;x=-152960000;
#10;x=-152950000;
#10;x=-152940000;
#10;x=-152930000;
#10;x=-152920000;
#10;x=-152910000;
#10;x=-152900000;
#10;x=-152890000;
#10;x=-152880000;
#10;x=-152870000;
#10;x=-152860000;
#10;x=-152850000;
#10;x=-152840000;
#10;x=-152830000;
#10;x=-152820000;
#10;x=-152810000;
#10;x=-152800000;
#10;x=-152790000;
#10;x=-152780000;
#10;x=-152770000;
#10;x=-152760000;
#10;x=-152750000;
#10;x=-152740000;
#10;x=-152730000;
#10;x=-152720000;
#10;x=-152710000;
#10;x=-152700000;
#10;x=-152690000;
#10;x=-152680000;
#10;x=-152670000;
#10;x=-152660000;
#10;x=-152650000;
#10;x=-152640000;
#10;x=-152630000;
#10;x=-152620000;
#10;x=-152610000;
#10;x=-152600000;
#10;x=-152590000;
#10;x=-152580000;
#10;x=-152570000;
#10;x=-152560000;
#10;x=-152550000;
#10;x=-152540000;
#10;x=-152530000;
#10;x=-152520000;
#10;x=-152510000;
#10;x=-152500000;
#10;x=-152490000;
#10;x=-152480000;
#10;x=-152470000;
#10;x=-152460000;
#10;x=-152450000;
#10;x=-152440000;
#10;x=-152430000;
#10;x=-152420000;
#10;x=-152410000;
#10;x=-152400000;
#10;x=-152390000;
#10;x=-152380000;
#10;x=-152370000;
#10;x=-152360000;
#10;x=-152350000;
#10;x=-152340000;
#10;x=-152330000;
#10;x=-152320000;
#10;x=-152310000;
#10;x=-152300000;
#10;x=-152290000;
#10;x=-152280000;
#10;x=-152270000;
#10;x=-152260000;
#10;x=-152250000;
#10;x=-152240000;
#10;x=-152230000;
#10;x=-152220000;
#10;x=-152210000;
#10;x=-152200000;
#10;x=-152190000;
#10;x=-152180000;
#10;x=-152170000;
#10;x=-152160000;
#10;x=-152150000;
#10;x=-152140000;
#10;x=-152130000;
#10;x=-152120000;
#10;x=-152110000;
#10;x=-152100000;
#10;x=-152090000;
#10;x=-152080000;
#10;x=-152070000;
#10;x=-152060000;
#10;x=-152050000;
#10;x=-152040000;
#10;x=-152030000;
#10;x=-152020000;
#10;x=-152010000;
#10;x=-152000000;
#10;x=-151990000;
#10;x=-151980000;
#10;x=-151970000;
#10;x=-151960000;
#10;x=-151950000;
#10;x=-151940000;
#10;x=-151930000;
#10;x=-151920000;
#10;x=-151910000;
#10;x=-151900000;
#10;x=-151890000;
#10;x=-151880000;
#10;x=-151870000;
#10;x=-151860000;
#10;x=-151850000;
#10;x=-151840000;
#10;x=-151830000;
#10;x=-151820000;
#10;x=-151810000;
#10;x=-151800000;
#10;x=-151790000;
#10;x=-151780000;
#10;x=-151770000;
#10;x=-151760000;
#10;x=-151750000;
#10;x=-151740000;
#10;x=-151730000;
#10;x=-151720000;
#10;x=-151710000;
#10;x=-151700000;
#10;x=-151690000;
#10;x=-151680000;
#10;x=-151670000;
#10;x=-151660000;
#10;x=-151650000;
#10;x=-151640000;
#10;x=-151630000;
#10;x=-151620000;
#10;x=-151610000;
#10;x=-151600000;
#10;x=-151590000;
#10;x=-151580000;
#10;x=-151570000;
#10;x=-151560000;
#10;x=-151550000;
#10;x=-151540000;
#10;x=-151530000;
#10;x=-151520000;
#10;x=-151510000;
#10;x=-151500000;
#10;x=-151490000;
#10;x=-151480000;
#10;x=-151470000;
#10;x=-151460000;
#10;x=-151450000;
#10;x=-151440000;
#10;x=-151430000;
#10;x=-151420000;
#10;x=-151410000;
#10;x=-151400000;
#10;x=-151390000;
#10;x=-151380000;
#10;x=-151370000;
#10;x=-151360000;
#10;x=-151350000;
#10;x=-151340000;
#10;x=-151330000;
#10;x=-151320000;
#10;x=-151310000;
#10;x=-151300000;
#10;x=-151290000;
#10;x=-151280000;
#10;x=-151270000;
#10;x=-151260000;
#10;x=-151250000;
#10;x=-151240000;
#10;x=-151230000;
#10;x=-151220000;
#10;x=-151210000;
#10;x=-151200000;
#10;x=-151190000;
#10;x=-151180000;
#10;x=-151170000;
#10;x=-151160000;
#10;x=-151150000;
#10;x=-151140000;
#10;x=-151130000;
#10;x=-151120000;
#10;x=-151110000;
#10;x=-151100000;
#10;x=-151090000;
#10;x=-151080000;
#10;x=-151070000;
#10;x=-151060000;
#10;x=-151050000;
#10;x=-151040000;
#10;x=-151030000;
#10;x=-151020000;
#10;x=-151010000;
#10;x=-151000000;
#10;x=-150990000;
#10;x=-150980000;
#10;x=-150970000;
#10;x=-150960000;
#10;x=-150950000;
#10;x=-150940000;
#10;x=-150930000;
#10;x=-150920000;
#10;x=-150910000;
#10;x=-150900000;
#10;x=-150890000;
#10;x=-150880000;
#10;x=-150870000;
#10;x=-150860000;
#10;x=-150850000;
#10;x=-150840000;
#10;x=-150830000;
#10;x=-150820000;
#10;x=-150810000;
#10;x=-150800000;
#10;x=-150790000;
#10;x=-150780000;
#10;x=-150770000;
#10;x=-150760000;
#10;x=-150750000;
#10;x=-150740000;
#10;x=-150730000;
#10;x=-150720000;
#10;x=-150710000;
#10;x=-150700000;
#10;x=-150690000;
#10;x=-150680000;
#10;x=-150670000;
#10;x=-150660000;
#10;x=-150650000;
#10;x=-150640000;
#10;x=-150630000;
#10;x=-150620000;
#10;x=-150610000;
#10;x=-150600000;
#10;x=-150590000;
#10;x=-150580000;
#10;x=-150570000;
#10;x=-150560000;
#10;x=-150550000;
#10;x=-150540000;
#10;x=-150530000;
#10;x=-150520000;
#10;x=-150510000;
#10;x=-150500000;
#10;x=-150490000;
#10;x=-150480000;
#10;x=-150470000;
#10;x=-150460000;
#10;x=-150450000;
#10;x=-150440000;
#10;x=-150430000;
#10;x=-150420000;
#10;x=-150410000;
#10;x=-150400000;
#10;x=-150390000;
#10;x=-150380000;
#10;x=-150370000;
#10;x=-150360000;
#10;x=-150350000;
#10;x=-150340000;
#10;x=-150330000;
#10;x=-150320000;
#10;x=-150310000;
#10;x=-150300000;
#10;x=-150290000;
#10;x=-150280000;
#10;x=-150270000;
#10;x=-150260000;
#10;x=-150250000;
#10;x=-150240000;
#10;x=-150230000;
#10;x=-150220000;
#10;x=-150210000;
#10;x=-150200000;
#10;x=-150190000;
#10;x=-150180000;
#10;x=-150170000;
#10;x=-150160000;
#10;x=-150150000;
#10;x=-150140000;
#10;x=-150130000;
#10;x=-150120000;
#10;x=-150110000;
#10;x=-150100000;
#10;x=-150090000;
#10;x=-150080000;
#10;x=-150070000;
#10;x=-150060000;
#10;x=-150050000;
#10;x=-150040000;
#10;x=-150030000;
#10;x=-150020000;
#10;x=-150010000;
#10;x=-150000000;
#10;x=-149990000;
#10;x=-149980000;
#10;x=-149970000;
#10;x=-149960000;
#10;x=-149950000;
#10;x=-149940000;
#10;x=-149930000;
#10;x=-149920000;
#10;x=-149910000;
#10;x=-149900000;
#10;x=-149890000;
#10;x=-149880000;
#10;x=-149870000;
#10;x=-149860000;
#10;x=-149850000;
#10;x=-149840000;
#10;x=-149830000;
#10;x=-149820000;
#10;x=-149810000;
#10;x=-149800000;
#10;x=-149790000;
#10;x=-149780000;
#10;x=-149770000;
#10;x=-149760000;
#10;x=-149750000;
#10;x=-149740000;
#10;x=-149730000;
#10;x=-149720000;
#10;x=-149710000;
#10;x=-149700000;
#10;x=-149690000;
#10;x=-149680000;
#10;x=-149670000;
#10;x=-149660000;
#10;x=-149650000;
#10;x=-149640000;
#10;x=-149630000;
#10;x=-149620000;
#10;x=-149610000;
#10;x=-149600000;
#10;x=-149590000;
#10;x=-149580000;
#10;x=-149570000;
#10;x=-149560000;
#10;x=-149550000;
#10;x=-149540000;
#10;x=-149530000;
#10;x=-149520000;
#10;x=-149510000;
#10;x=-149500000;
#10;x=-149490000;
#10;x=-149480000;
#10;x=-149470000;
#10;x=-149460000;
#10;x=-149450000;
#10;x=-149440000;
#10;x=-149430000;
#10;x=-149420000;
#10;x=-149410000;
#10;x=-149400000;
#10;x=-149390000;
#10;x=-149380000;
#10;x=-149370000;
#10;x=-149360000;
#10;x=-149350000;
#10;x=-149340000;
#10;x=-149330000;
#10;x=-149320000;
#10;x=-149310000;
#10;x=-149300000;
#10;x=-149290000;
#10;x=-149280000;
#10;x=-149270000;
#10;x=-149260000;
#10;x=-149250000;
#10;x=-149240000;
#10;x=-149230000;
#10;x=-149220000;
#10;x=-149210000;
#10;x=-149200000;
#10;x=-149190000;
#10;x=-149180000;
#10;x=-149170000;
#10;x=-149160000;
#10;x=-149150000;
#10;x=-149140000;
#10;x=-149130000;
#10;x=-149120000;
#10;x=-149110000;
#10;x=-149100000;
#10;x=-149090000;
#10;x=-149080000;
#10;x=-149070000;
#10;x=-149060000;
#10;x=-149050000;
#10;x=-149040000;
#10;x=-149030000;
#10;x=-149020000;
#10;x=-149010000;
#10;x=-149000000;
#10;x=-148990000;
#10;x=-148980000;
#10;x=-148970000;
#10;x=-148960000;
#10;x=-148950000;
#10;x=-148940000;
#10;x=-148930000;
#10;x=-148920000;
#10;x=-148910000;
#10;x=-148900000;
#10;x=-148890000;
#10;x=-148880000;
#10;x=-148870000;
#10;x=-148860000;
#10;x=-148850000;
#10;x=-148840000;
#10;x=-148830000;
#10;x=-148820000;
#10;x=-148810000;
#10;x=-148800000;
#10;x=-148790000;
#10;x=-148780000;
#10;x=-148770000;
#10;x=-148760000;
#10;x=-148750000;
#10;x=-148740000;
#10;x=-148730000;
#10;x=-148720000;
#10;x=-148710000;
#10;x=-148700000;
#10;x=-148690000;
#10;x=-148680000;
#10;x=-148670000;
#10;x=-148660000;
#10;x=-148650000;
#10;x=-148640000;
#10;x=-148630000;
#10;x=-148620000;
#10;x=-148610000;
#10;x=-148600000;
#10;x=-148590000;
#10;x=-148580000;
#10;x=-148570000;
#10;x=-148560000;
#10;x=-148550000;
#10;x=-148540000;
#10;x=-148530000;
#10;x=-148520000;
#10;x=-148510000;
#10;x=-148500000;
#10;x=-148490000;
#10;x=-148480000;
#10;x=-148470000;
#10;x=-148460000;
#10;x=-148450000;
#10;x=-148440000;
#10;x=-148430000;
#10;x=-148420000;
#10;x=-148410000;
#10;x=-148400000;
#10;x=-148390000;
#10;x=-148380000;
#10;x=-148370000;
#10;x=-148360000;
#10;x=-148350000;
#10;x=-148340000;
#10;x=-148330000;
#10;x=-148320000;
#10;x=-148310000;
#10;x=-148300000;
#10;x=-148290000;
#10;x=-148280000;
#10;x=-148270000;
#10;x=-148260000;
#10;x=-148250000;
#10;x=-148240000;
#10;x=-148230000;
#10;x=-148220000;
#10;x=-148210000;
#10;x=-148200000;
#10;x=-148190000;
#10;x=-148180000;
#10;x=-148170000;
#10;x=-148160000;
#10;x=-148150000;
#10;x=-148140000;
#10;x=-148130000;
#10;x=-148120000;
#10;x=-148110000;
#10;x=-148100000;
#10;x=-148090000;
#10;x=-148080000;
#10;x=-148070000;
#10;x=-148060000;
#10;x=-148050000;
#10;x=-148040000;
#10;x=-148030000;
#10;x=-148020000;
#10;x=-148010000;
#10;x=-148000000;
#10;x=-147990000;
#10;x=-147980000;
#10;x=-147970000;
#10;x=-147960000;
#10;x=-147950000;
#10;x=-147940000;
#10;x=-147930000;
#10;x=-147920000;
#10;x=-147910000;
#10;x=-147900000;
#10;x=-147890000;
#10;x=-147880000;
#10;x=-147870000;
#10;x=-147860000;
#10;x=-147850000;
#10;x=-147840000;
#10;x=-147830000;
#10;x=-147820000;
#10;x=-147810000;
#10;x=-147800000;
#10;x=-147790000;
#10;x=-147780000;
#10;x=-147770000;
#10;x=-147760000;
#10;x=-147750000;
#10;x=-147740000;
#10;x=-147730000;
#10;x=-147720000;
#10;x=-147710000;
#10;x=-147700000;
#10;x=-147690000;
#10;x=-147680000;
#10;x=-147670000;
#10;x=-147660000;
#10;x=-147650000;
#10;x=-147640000;
#10;x=-147630000;
#10;x=-147620000;
#10;x=-147610000;
#10;x=-147600000;
#10;x=-147590000;
#10;x=-147580000;
#10;x=-147570000;
#10;x=-147560000;
#10;x=-147550000;
#10;x=-147540000;
#10;x=-147530000;
#10;x=-147520000;
#10;x=-147510000;
#10;x=-147500000;
#10;x=-147490000;
#10;x=-147480000;
#10;x=-147470000;
#10;x=-147460000;
#10;x=-147450000;
#10;x=-147440000;
#10;x=-147430000;
#10;x=-147420000;
#10;x=-147410000;
#10;x=-147400000;
#10;x=-147390000;
#10;x=-147380000;
#10;x=-147370000;
#10;x=-147360000;
#10;x=-147350000;
#10;x=-147340000;
#10;x=-147330000;
#10;x=-147320000;
#10;x=-147310000;
#10;x=-147300000;
#10;x=-147290000;
#10;x=-147280000;
#10;x=-147270000;
#10;x=-147260000;
#10;x=-147250000;
#10;x=-147240000;
#10;x=-147230000;
#10;x=-147220000;
#10;x=-147210000;
#10;x=-147200000;
#10;x=-147190000;
#10;x=-147180000;
#10;x=-147170000;
#10;x=-147160000;
#10;x=-147150000;
#10;x=-147140000;
#10;x=-147130000;
#10;x=-147120000;
#10;x=-147110000;
#10;x=-147100000;
#10;x=-147090000;
#10;x=-147080000;
#10;x=-147070000;
#10;x=-147060000;
#10;x=-147050000;
#10;x=-147040000;
#10;x=-147030000;
#10;x=-147020000;
#10;x=-147010000;
#10;x=-147000000;
#10;x=-146990000;
#10;x=-146980000;
#10;x=-146970000;
#10;x=-146960000;
#10;x=-146950000;
#10;x=-146940000;
#10;x=-146930000;
#10;x=-146920000;
#10;x=-146910000;
#10;x=-146900000;
#10;x=-146890000;
#10;x=-146880000;
#10;x=-146870000;
#10;x=-146860000;
#10;x=-146850000;
#10;x=-146840000;
#10;x=-146830000;
#10;x=-146820000;
#10;x=-146810000;
#10;x=-146800000;
#10;x=-146790000;
#10;x=-146780000;
#10;x=-146770000;
#10;x=-146760000;
#10;x=-146750000;
#10;x=-146740000;
#10;x=-146730000;
#10;x=-146720000;
#10;x=-146710000;
#10;x=-146700000;
#10;x=-146690000;
#10;x=-146680000;
#10;x=-146670000;
#10;x=-146660000;
#10;x=-146650000;
#10;x=-146640000;
#10;x=-146630000;
#10;x=-146620000;
#10;x=-146610000;
#10;x=-146600000;
#10;x=-146590000;
#10;x=-146580000;
#10;x=-146570000;
#10;x=-146560000;
#10;x=-146550000;
#10;x=-146540000;
#10;x=-146530000;
#10;x=-146520000;
#10;x=-146510000;
#10;x=-146500000;
#10;x=-146490000;
#10;x=-146480000;
#10;x=-146470000;
#10;x=-146460000;
#10;x=-146450000;
#10;x=-146440000;
#10;x=-146430000;
#10;x=-146420000;
#10;x=-146410000;
#10;x=-146400000;
#10;x=-146390000;
#10;x=-146380000;
#10;x=-146370000;
#10;x=-146360000;
#10;x=-146350000;
#10;x=-146340000;
#10;x=-146330000;
#10;x=-146320000;
#10;x=-146310000;
#10;x=-146300000;
#10;x=-146290000;
#10;x=-146280000;
#10;x=-146270000;
#10;x=-146260000;
#10;x=-146250000;
#10;x=-146240000;
#10;x=-146230000;
#10;x=-146220000;
#10;x=-146210000;
#10;x=-146200000;
#10;x=-146190000;
#10;x=-146180000;
#10;x=-146170000;
#10;x=-146160000;
#10;x=-146150000;
#10;x=-146140000;
#10;x=-146130000;
#10;x=-146120000;
#10;x=-146110000;
#10;x=-146100000;
#10;x=-146090000;
#10;x=-146080000;
#10;x=-146070000;
#10;x=-146060000;
#10;x=-146050000;
#10;x=-146040000;
#10;x=-146030000;
#10;x=-146020000;
#10;x=-146010000;
#10;x=-146000000;
#10;x=-145990000;
#10;x=-145980000;
#10;x=-145970000;
#10;x=-145960000;
#10;x=-145950000;
#10;x=-145940000;
#10;x=-145930000;
#10;x=-145920000;
#10;x=-145910000;
#10;x=-145900000;
#10;x=-145890000;
#10;x=-145880000;
#10;x=-145870000;
#10;x=-145860000;
#10;x=-145850000;
#10;x=-145840000;
#10;x=-145830000;
#10;x=-145820000;
#10;x=-145810000;
#10;x=-145800000;
#10;x=-145790000;
#10;x=-145780000;
#10;x=-145770000;
#10;x=-145760000;
#10;x=-145750000;
#10;x=-145740000;
#10;x=-145730000;
#10;x=-145720000;
#10;x=-145710000;
#10;x=-145700000;
#10;x=-145690000;
#10;x=-145680000;
#10;x=-145670000;
#10;x=-145660000;
#10;x=-145650000;
#10;x=-145640000;
#10;x=-145630000;
#10;x=-145620000;
#10;x=-145610000;
#10;x=-145600000;
#10;x=-145590000;
#10;x=-145580000;
#10;x=-145570000;
#10;x=-145560000;
#10;x=-145550000;
#10;x=-145540000;
#10;x=-145530000;
#10;x=-145520000;
#10;x=-145510000;
#10;x=-145500000;
#10;x=-145490000;
#10;x=-145480000;
#10;x=-145470000;
#10;x=-145460000;
#10;x=-145450000;
#10;x=-145440000;
#10;x=-145430000;
#10;x=-145420000;
#10;x=-145410000;
#10;x=-145400000;
#10;x=-145390000;
#10;x=-145380000;
#10;x=-145370000;
#10;x=-145360000;
#10;x=-145350000;
#10;x=-145340000;
#10;x=-145330000;
#10;x=-145320000;
#10;x=-145310000;
#10;x=-145300000;
#10;x=-145290000;
#10;x=-145280000;
#10;x=-145270000;
#10;x=-145260000;
#10;x=-145250000;
#10;x=-145240000;
#10;x=-145230000;
#10;x=-145220000;
#10;x=-145210000;
#10;x=-145200000;
#10;x=-145190000;
#10;x=-145180000;
#10;x=-145170000;
#10;x=-145160000;
#10;x=-145150000;
#10;x=-145140000;
#10;x=-145130000;
#10;x=-145120000;
#10;x=-145110000;
#10;x=-145100000;
#10;x=-145090000;
#10;x=-145080000;
#10;x=-145070000;
#10;x=-145060000;
#10;x=-145050000;
#10;x=-145040000;
#10;x=-145030000;
#10;x=-145020000;
#10;x=-145010000;
#10;x=-145000000;
#10;x=-144990000;
#10;x=-144980000;
#10;x=-144970000;
#10;x=-144960000;
#10;x=-144950000;
#10;x=-144940000;
#10;x=-144930000;
#10;x=-144920000;
#10;x=-144910000;
#10;x=-144900000;
#10;x=-144890000;
#10;x=-144880000;
#10;x=-144870000;
#10;x=-144860000;
#10;x=-144850000;
#10;x=-144840000;
#10;x=-144830000;
#10;x=-144820000;
#10;x=-144810000;
#10;x=-144800000;
#10;x=-144790000;
#10;x=-144780000;
#10;x=-144770000;
#10;x=-144760000;
#10;x=-144750000;
#10;x=-144740000;
#10;x=-144730000;
#10;x=-144720000;
#10;x=-144710000;
#10;x=-144700000;
#10;x=-144690000;
#10;x=-144680000;
#10;x=-144670000;
#10;x=-144660000;
#10;x=-144650000;
#10;x=-144640000;
#10;x=-144630000;
#10;x=-144620000;
#10;x=-144610000;
#10;x=-144600000;
#10;x=-144590000;
#10;x=-144580000;
#10;x=-144570000;
#10;x=-144560000;
#10;x=-144550000;
#10;x=-144540000;
#10;x=-144530000;
#10;x=-144520000;
#10;x=-144510000;
#10;x=-144500000;
#10;x=-144490000;
#10;x=-144480000;
#10;x=-144470000;
#10;x=-144460000;
#10;x=-144450000;
#10;x=-144440000;
#10;x=-144430000;
#10;x=-144420000;
#10;x=-144410000;
#10;x=-144400000;
#10;x=-144390000;
#10;x=-144380000;
#10;x=-144370000;
#10;x=-144360000;
#10;x=-144350000;
#10;x=-144340000;
#10;x=-144330000;
#10;x=-144320000;
#10;x=-144310000;
#10;x=-144300000;
#10;x=-144290000;
#10;x=-144280000;
#10;x=-144270000;
#10;x=-144260000;
#10;x=-144250000;
#10;x=-144240000;
#10;x=-144230000;
#10;x=-144220000;
#10;x=-144210000;
#10;x=-144200000;
#10;x=-144190000;
#10;x=-144180000;
#10;x=-144170000;
#10;x=-144160000;
#10;x=-144150000;
#10;x=-144140000;
#10;x=-144130000;
#10;x=-144120000;
#10;x=-144110000;
#10;x=-144100000;
#10;x=-144090000;
#10;x=-144080000;
#10;x=-144070000;
#10;x=-144060000;
#10;x=-144050000;
#10;x=-144040000;
#10;x=-144030000;
#10;x=-144020000;
#10;x=-144010000;
#10;x=-144000000;
#10;x=-143990000;
#10;x=-143980000;
#10;x=-143970000;
#10;x=-143960000;
#10;x=-143950000;
#10;x=-143940000;
#10;x=-143930000;
#10;x=-143920000;
#10;x=-143910000;
#10;x=-143900000;
#10;x=-143890000;
#10;x=-143880000;
#10;x=-143870000;
#10;x=-143860000;
#10;x=-143850000;
#10;x=-143840000;
#10;x=-143830000;
#10;x=-143820000;
#10;x=-143810000;
#10;x=-143800000;
#10;x=-143790000;
#10;x=-143780000;
#10;x=-143770000;
#10;x=-143760000;
#10;x=-143750000;
#10;x=-143740000;
#10;x=-143730000;
#10;x=-143720000;
#10;x=-143710000;
#10;x=-143700000;
#10;x=-143690000;
#10;x=-143680000;
#10;x=-143670000;
#10;x=-143660000;
#10;x=-143650000;
#10;x=-143640000;
#10;x=-143630000;
#10;x=-143620000;
#10;x=-143610000;
#10;x=-143600000;
#10;x=-143590000;
#10;x=-143580000;
#10;x=-143570000;
#10;x=-143560000;
#10;x=-143550000;
#10;x=-143540000;
#10;x=-143530000;
#10;x=-143520000;
#10;x=-143510000;
#10;x=-143500000;
#10;x=-143490000;
#10;x=-143480000;
#10;x=-143470000;
#10;x=-143460000;
#10;x=-143450000;
#10;x=-143440000;
#10;x=-143430000;
#10;x=-143420000;
#10;x=-143410000;
#10;x=-143400000;
#10;x=-143390000;
#10;x=-143380000;
#10;x=-143370000;
#10;x=-143360000;
#10;x=-143350000;
#10;x=-143340000;
#10;x=-143330000;
#10;x=-143320000;
#10;x=-143310000;
#10;x=-143300000;
#10;x=-143290000;
#10;x=-143280000;
#10;x=-143270000;
#10;x=-143260000;
#10;x=-143250000;
#10;x=-143240000;
#10;x=-143230000;
#10;x=-143220000;
#10;x=-143210000;
#10;x=-143200000;
#10;x=-143190000;
#10;x=-143180000;
#10;x=-143170000;
#10;x=-143160000;
#10;x=-143150000;
#10;x=-143140000;
#10;x=-143130000;
#10;x=-143120000;
#10;x=-143110000;
#10;x=-143100000;
#10;x=-143090000;
#10;x=-143080000;
#10;x=-143070000;
#10;x=-143060000;
#10;x=-143050000;
#10;x=-143040000;
#10;x=-143030000;
#10;x=-143020000;
#10;x=-143010000;
#10;x=-143000000;
#10;x=-142990000;
#10;x=-142980000;
#10;x=-142970000;
#10;x=-142960000;
#10;x=-142950000;
#10;x=-142940000;
#10;x=-142930000;
#10;x=-142920000;
#10;x=-142910000;
#10;x=-142900000;
#10;x=-142890000;
#10;x=-142880000;
#10;x=-142870000;
#10;x=-142860000;
#10;x=-142850000;
#10;x=-142840000;
#10;x=-142830000;
#10;x=-142820000;
#10;x=-142810000;
#10;x=-142800000;
#10;x=-142790000;
#10;x=-142780000;
#10;x=-142770000;
#10;x=-142760000;
#10;x=-142750000;
#10;x=-142740000;
#10;x=-142730000;
#10;x=-142720000;
#10;x=-142710000;
#10;x=-142700000;
#10;x=-142690000;
#10;x=-142680000;
#10;x=-142670000;
#10;x=-142660000;
#10;x=-142650000;
#10;x=-142640000;
#10;x=-142630000;
#10;x=-142620000;
#10;x=-142610000;
#10;x=-142600000;
#10;x=-142590000;
#10;x=-142580000;
#10;x=-142570000;
#10;x=-142560000;
#10;x=-142550000;
#10;x=-142540000;
#10;x=-142530000;
#10;x=-142520000;
#10;x=-142510000;
#10;x=-142500000;
#10;x=-142490000;
#10;x=-142480000;
#10;x=-142470000;
#10;x=-142460000;
#10;x=-142450000;
#10;x=-142440000;
#10;x=-142430000;
#10;x=-142420000;
#10;x=-142410000;
#10;x=-142400000;
#10;x=-142390000;
#10;x=-142380000;
#10;x=-142370000;
#10;x=-142360000;
#10;x=-142350000;
#10;x=-142340000;
#10;x=-142330000;
#10;x=-142320000;
#10;x=-142310000;
#10;x=-142300000;
#10;x=-142290000;
#10;x=-142280000;
#10;x=-142270000;
#10;x=-142260000;
#10;x=-142250000;
#10;x=-142240000;
#10;x=-142230000;
#10;x=-142220000;
#10;x=-142210000;
#10;x=-142200000;
#10;x=-142190000;
#10;x=-142180000;
#10;x=-142170000;
#10;x=-142160000;
#10;x=-142150000;
#10;x=-142140000;
#10;x=-142130000;
#10;x=-142120000;
#10;x=-142110000;
#10;x=-142100000;
#10;x=-142090000;
#10;x=-142080000;
#10;x=-142070000;
#10;x=-142060000;
#10;x=-142050000;
#10;x=-142040000;
#10;x=-142030000;
#10;x=-142020000;
#10;x=-142010000;
#10;x=-142000000;
#10;x=-141990000;
#10;x=-141980000;
#10;x=-141970000;
#10;x=-141960000;
#10;x=-141950000;
#10;x=-141940000;
#10;x=-141930000;
#10;x=-141920000;
#10;x=-141910000;
#10;x=-141900000;
#10;x=-141890000;
#10;x=-141880000;
#10;x=-141870000;
#10;x=-141860000;
#10;x=-141850000;
#10;x=-141840000;
#10;x=-141830000;
#10;x=-141820000;
#10;x=-141810000;
#10;x=-141800000;
#10;x=-141790000;
#10;x=-141780000;
#10;x=-141770000;
#10;x=-141760000;
#10;x=-141750000;
#10;x=-141740000;
#10;x=-141730000;
#10;x=-141720000;
#10;x=-141710000;
#10;x=-141700000;
#10;x=-141690000;
#10;x=-141680000;
#10;x=-141670000;
#10;x=-141660000;
#10;x=-141650000;
#10;x=-141640000;
#10;x=-141630000;
#10;x=-141620000;
#10;x=-141610000;
#10;x=-141600000;
#10;x=-141590000;
#10;x=-141580000;
#10;x=-141570000;
#10;x=-141560000;
#10;x=-141550000;
#10;x=-141540000;
#10;x=-141530000;
#10;x=-141520000;
#10;x=-141510000;
#10;x=-141500000;
#10;x=-141490000;
#10;x=-141480000;
#10;x=-141470000;
#10;x=-141460000;
#10;x=-141450000;
#10;x=-141440000;
#10;x=-141430000;
#10;x=-141420000;
#10;x=-141410000;
#10;x=-141400000;
#10;x=-141390000;
#10;x=-141380000;
#10;x=-141370000;
#10;x=-141360000;
#10;x=-141350000;
#10;x=-141340000;
#10;x=-141330000;
#10;x=-141320000;
#10;x=-141310000;
#10;x=-141300000;
#10;x=-141290000;
#10;x=-141280000;
#10;x=-141270000;
#10;x=-141260000;
#10;x=-141250000;
#10;x=-141240000;
#10;x=-141230000;
#10;x=-141220000;
#10;x=-141210000;
#10;x=-141200000;
#10;x=-141190000;
#10;x=-141180000;
#10;x=-141170000;
#10;x=-141160000;
#10;x=-141150000;
#10;x=-141140000;
#10;x=-141130000;
#10;x=-141120000;
#10;x=-141110000;
#10;x=-141100000;
#10;x=-141090000;
#10;x=-141080000;
#10;x=-141070000;
#10;x=-141060000;
#10;x=-141050000;
#10;x=-141040000;
#10;x=-141030000;
#10;x=-141020000;
#10;x=-141010000;
#10;x=-141000000;
#10;x=-140990000;
#10;x=-140980000;
#10;x=-140970000;
#10;x=-140960000;
#10;x=-140950000;
#10;x=-140940000;
#10;x=-140930000;
#10;x=-140920000;
#10;x=-140910000;
#10;x=-140900000;
#10;x=-140890000;
#10;x=-140880000;
#10;x=-140870000;
#10;x=-140860000;
#10;x=-140850000;
#10;x=-140840000;
#10;x=-140830000;
#10;x=-140820000;
#10;x=-140810000;
#10;x=-140800000;
#10;x=-140790000;
#10;x=-140780000;
#10;x=-140770000;
#10;x=-140760000;
#10;x=-140750000;
#10;x=-140740000;
#10;x=-140730000;
#10;x=-140720000;
#10;x=-140710000;
#10;x=-140700000;
#10;x=-140690000;
#10;x=-140680000;
#10;x=-140670000;
#10;x=-140660000;
#10;x=-140650000;
#10;x=-140640000;
#10;x=-140630000;
#10;x=-140620000;
#10;x=-140610000;
#10;x=-140600000;
#10;x=-140590000;
#10;x=-140580000;
#10;x=-140570000;
#10;x=-140560000;
#10;x=-140550000;
#10;x=-140540000;
#10;x=-140530000;
#10;x=-140520000;
#10;x=-140510000;
#10;x=-140500000;
#10;x=-140490000;
#10;x=-140480000;
#10;x=-140470000;
#10;x=-140460000;
#10;x=-140450000;
#10;x=-140440000;
#10;x=-140430000;
#10;x=-140420000;
#10;x=-140410000;
#10;x=-140400000;
#10;x=-140390000;
#10;x=-140380000;
#10;x=-140370000;
#10;x=-140360000;
#10;x=-140350000;
#10;x=-140340000;
#10;x=-140330000;
#10;x=-140320000;
#10;x=-140310000;
#10;x=-140300000;
#10;x=-140290000;
#10;x=-140280000;
#10;x=-140270000;
#10;x=-140260000;
#10;x=-140250000;
#10;x=-140240000;
#10;x=-140230000;
#10;x=-140220000;
#10;x=-140210000;
#10;x=-140200000;
#10;x=-140190000;
#10;x=-140180000;
#10;x=-140170000;
#10;x=-140160000;
#10;x=-140150000;
#10;x=-140140000;
#10;x=-140130000;
#10;x=-140120000;
#10;x=-140110000;
#10;x=-140100000;
#10;x=-140090000;
#10;x=-140080000;
#10;x=-140070000;
#10;x=-140060000;
#10;x=-140050000;
#10;x=-140040000;
#10;x=-140030000;
#10;x=-140020000;
#10;x=-140010000;
#10;x=-140000000;
#10;x=-139990000;
#10;x=-139980000;
#10;x=-139970000;
#10;x=-139960000;
#10;x=-139950000;
#10;x=-139940000;
#10;x=-139930000;
#10;x=-139920000;
#10;x=-139910000;
#10;x=-139900000;
#10;x=-139890000;
#10;x=-139880000;
#10;x=-139870000;
#10;x=-139860000;
#10;x=-139850000;
#10;x=-139840000;
#10;x=-139830000;
#10;x=-139820000;
#10;x=-139810000;
#10;x=-139800000;
#10;x=-139790000;
#10;x=-139780000;
#10;x=-139770000;
#10;x=-139760000;
#10;x=-139750000;
#10;x=-139740000;
#10;x=-139730000;
#10;x=-139720000;
#10;x=-139710000;
#10;x=-139700000;
#10;x=-139690000;
#10;x=-139680000;
#10;x=-139670000;
#10;x=-139660000;
#10;x=-139650000;
#10;x=-139640000;
#10;x=-139630000;
#10;x=-139620000;
#10;x=-139610000;
#10;x=-139600000;
#10;x=-139590000;
#10;x=-139580000;
#10;x=-139570000;
#10;x=-139560000;
#10;x=-139550000;
#10;x=-139540000;
#10;x=-139530000;
#10;x=-139520000;
#10;x=-139510000;
#10;x=-139500000;
#10;x=-139490000;
#10;x=-139480000;
#10;x=-139470000;
#10;x=-139460000;
#10;x=-139450000;
#10;x=-139440000;
#10;x=-139430000;
#10;x=-139420000;
#10;x=-139410000;
#10;x=-139400000;
#10;x=-139390000;
#10;x=-139380000;
#10;x=-139370000;
#10;x=-139360000;
#10;x=-139350000;
#10;x=-139340000;
#10;x=-139330000;
#10;x=-139320000;
#10;x=-139310000;
#10;x=-139300000;
#10;x=-139290000;
#10;x=-139280000;
#10;x=-139270000;
#10;x=-139260000;
#10;x=-139250000;
#10;x=-139240000;
#10;x=-139230000;
#10;x=-139220000;
#10;x=-139210000;
#10;x=-139200000;
#10;x=-139190000;
#10;x=-139180000;
#10;x=-139170000;
#10;x=-139160000;
#10;x=-139150000;
#10;x=-139140000;
#10;x=-139130000;
#10;x=-139120000;
#10;x=-139110000;
#10;x=-139100000;
#10;x=-139090000;
#10;x=-139080000;
#10;x=-139070000;
#10;x=-139060000;
#10;x=-139050000;
#10;x=-139040000;
#10;x=-139030000;
#10;x=-139020000;
#10;x=-139010000;
#10;x=-139000000;
#10;x=-138990000;
#10;x=-138980000;
#10;x=-138970000;
#10;x=-138960000;
#10;x=-138950000;
#10;x=-138940000;
#10;x=-138930000;
#10;x=-138920000;
#10;x=-138910000;
#10;x=-138900000;
#10;x=-138890000;
#10;x=-138880000;
#10;x=-138870000;
#10;x=-138860000;
#10;x=-138850000;
#10;x=-138840000;
#10;x=-138830000;
#10;x=-138820000;
#10;x=-138810000;
#10;x=-138800000;
#10;x=-138790000;
#10;x=-138780000;
#10;x=-138770000;
#10;x=-138760000;
#10;x=-138750000;
#10;x=-138740000;
#10;x=-138730000;
#10;x=-138720000;
#10;x=-138710000;
#10;x=-138700000;
#10;x=-138690000;
#10;x=-138680000;
#10;x=-138670000;
#10;x=-138660000;
#10;x=-138650000;
#10;x=-138640000;
#10;x=-138630000;
#10;x=-138620000;
#10;x=-138610000;
#10;x=-138600000;
#10;x=-138590000;
#10;x=-138580000;
#10;x=-138570000;
#10;x=-138560000;
#10;x=-138550000;
#10;x=-138540000;
#10;x=-138530000;
#10;x=-138520000;
#10;x=-138510000;
#10;x=-138500000;
#10;x=-138490000;
#10;x=-138480000;
#10;x=-138470000;
#10;x=-138460000;
#10;x=-138450000;
#10;x=-138440000;
#10;x=-138430000;
#10;x=-138420000;
#10;x=-138410000;
#10;x=-138400000;
#10;x=-138390000;
#10;x=-138380000;
#10;x=-138370000;
#10;x=-138360000;
#10;x=-138350000;
#10;x=-138340000;
#10;x=-138330000;
#10;x=-138320000;
#10;x=-138310000;
#10;x=-138300000;
#10;x=-138290000;
#10;x=-138280000;
#10;x=-138270000;
#10;x=-138260000;
#10;x=-138250000;
#10;x=-138240000;
#10;x=-138230000;
#10;x=-138220000;
#10;x=-138210000;
#10;x=-138200000;
#10;x=-138190000;
#10;x=-138180000;
#10;x=-138170000;
#10;x=-138160000;
#10;x=-138150000;
#10;x=-138140000;
#10;x=-138130000;
#10;x=-138120000;
#10;x=-138110000;
#10;x=-138100000;
#10;x=-138090000;
#10;x=-138080000;
#10;x=-138070000;
#10;x=-138060000;
#10;x=-138050000;
#10;x=-138040000;
#10;x=-138030000;
#10;x=-138020000;
#10;x=-138010000;
#10;x=-138000000;
#10;x=-137990000;
#10;x=-137980000;
#10;x=-137970000;
#10;x=-137960000;
#10;x=-137950000;
#10;x=-137940000;
#10;x=-137930000;
#10;x=-137920000;
#10;x=-137910000;
#10;x=-137900000;
#10;x=-137890000;
#10;x=-137880000;
#10;x=-137870000;
#10;x=-137860000;
#10;x=-137850000;
#10;x=-137840000;
#10;x=-137830000;
#10;x=-137820000;
#10;x=-137810000;
#10;x=-137800000;
#10;x=-137790000;
#10;x=-137780000;
#10;x=-137770000;
#10;x=-137760000;
#10;x=-137750000;
#10;x=-137740000;
#10;x=-137730000;
#10;x=-137720000;
#10;x=-137710000;
#10;x=-137700000;
#10;x=-137690000;
#10;x=-137680000;
#10;x=-137670000;
#10;x=-137660000;
#10;x=-137650000;
#10;x=-137640000;
#10;x=-137630000;
#10;x=-137620000;
#10;x=-137610000;
#10;x=-137600000;
#10;x=-137590000;
#10;x=-137580000;
#10;x=-137570000;
#10;x=-137560000;
#10;x=-137550000;
#10;x=-137540000;
#10;x=-137530000;
#10;x=-137520000;
#10;x=-137510000;
#10;x=-137500000;
#10;x=-137490000;
#10;x=-137480000;
#10;x=-137470000;
#10;x=-137460000;
#10;x=-137450000;
#10;x=-137440000;
#10;x=-137430000;
#10;x=-137420000;
#10;x=-137410000;
#10;x=-137400000;
#10;x=-137390000;
#10;x=-137380000;
#10;x=-137370000;
#10;x=-137360000;
#10;x=-137350000;
#10;x=-137340000;
#10;x=-137330000;
#10;x=-137320000;
#10;x=-137310000;
#10;x=-137300000;
#10;x=-137290000;
#10;x=-137280000;
#10;x=-137270000;
#10;x=-137260000;
#10;x=-137250000;
#10;x=-137240000;
#10;x=-137230000;
#10;x=-137220000;
#10;x=-137210000;
#10;x=-137200000;
#10;x=-137190000;
#10;x=-137180000;
#10;x=-137170000;
#10;x=-137160000;
#10;x=-137150000;
#10;x=-137140000;
#10;x=-137130000;
#10;x=-137120000;
#10;x=-137110000;
#10;x=-137100000;
#10;x=-137090000;
#10;x=-137080000;
#10;x=-137070000;
#10;x=-137060000;
#10;x=-137050000;
#10;x=-137040000;
#10;x=-137030000;
#10;x=-137020000;
#10;x=-137010000;
#10;x=-137000000;
#10;x=-136990000;
#10;x=-136980000;
#10;x=-136970000;
#10;x=-136960000;
#10;x=-136950000;
#10;x=-136940000;
#10;x=-136930000;
#10;x=-136920000;
#10;x=-136910000;
#10;x=-136900000;
#10;x=-136890000;
#10;x=-136880000;
#10;x=-136870000;
#10;x=-136860000;
#10;x=-136850000;
#10;x=-136840000;
#10;x=-136830000;
#10;x=-136820000;
#10;x=-136810000;
#10;x=-136800000;
#10;x=-136790000;
#10;x=-136780000;
#10;x=-136770000;
#10;x=-136760000;
#10;x=-136750000;
#10;x=-136740000;
#10;x=-136730000;
#10;x=-136720000;
#10;x=-136710000;
#10;x=-136700000;
#10;x=-136690000;
#10;x=-136680000;
#10;x=-136670000;
#10;x=-136660000;
#10;x=-136650000;
#10;x=-136640000;
#10;x=-136630000;
#10;x=-136620000;
#10;x=-136610000;
#10;x=-136600000;
#10;x=-136590000;
#10;x=-136580000;
#10;x=-136570000;
#10;x=-136560000;
#10;x=-136550000;
#10;x=-136540000;
#10;x=-136530000;
#10;x=-136520000;
#10;x=-136510000;
#10;x=-136500000;
#10;x=-136490000;
#10;x=-136480000;
#10;x=-136470000;
#10;x=-136460000;
#10;x=-136450000;
#10;x=-136440000;
#10;x=-136430000;
#10;x=-136420000;
#10;x=-136410000;
#10;x=-136400000;
#10;x=-136390000;
#10;x=-136380000;
#10;x=-136370000;
#10;x=-136360000;
#10;x=-136350000;
#10;x=-136340000;
#10;x=-136330000;
#10;x=-136320000;
#10;x=-136310000;
#10;x=-136300000;
#10;x=-136290000;
#10;x=-136280000;
#10;x=-136270000;
#10;x=-136260000;
#10;x=-136250000;
#10;x=-136240000;
#10;x=-136230000;
#10;x=-136220000;
#10;x=-136210000;
#10;x=-136200000;
#10;x=-136190000;
#10;x=-136180000;
#10;x=-136170000;
#10;x=-136160000;
#10;x=-136150000;
#10;x=-136140000;
#10;x=-136130000;
#10;x=-136120000;
#10;x=-136110000;
#10;x=-136100000;
#10;x=-136090000;
#10;x=-136080000;
#10;x=-136070000;
#10;x=-136060000;
#10;x=-136050000;
#10;x=-136040000;
#10;x=-136030000;
#10;x=-136020000;
#10;x=-136010000;
#10;x=-136000000;
#10;x=-135990000;
#10;x=-135980000;
#10;x=-135970000;
#10;x=-135960000;
#10;x=-135950000;
#10;x=-135940000;
#10;x=-135930000;
#10;x=-135920000;
#10;x=-135910000;
#10;x=-135900000;
#10;x=-135890000;
#10;x=-135880000;
#10;x=-135870000;
#10;x=-135860000;
#10;x=-135850000;
#10;x=-135840000;
#10;x=-135830000;
#10;x=-135820000;
#10;x=-135810000;
#10;x=-135800000;
#10;x=-135790000;
#10;x=-135780000;
#10;x=-135770000;
#10;x=-135760000;
#10;x=-135750000;
#10;x=-135740000;
#10;x=-135730000;
#10;x=-135720000;
#10;x=-135710000;
#10;x=-135700000;
#10;x=-135690000;
#10;x=-135680000;
#10;x=-135670000;
#10;x=-135660000;
#10;x=-135650000;
#10;x=-135640000;
#10;x=-135630000;
#10;x=-135620000;
#10;x=-135610000;
#10;x=-135600000;
#10;x=-135590000;
#10;x=-135580000;
#10;x=-135570000;
#10;x=-135560000;
#10;x=-135550000;
#10;x=-135540000;
#10;x=-135530000;
#10;x=-135520000;
#10;x=-135510000;
#10;x=-135500000;
#10;x=-135490000;
#10;x=-135480000;
#10;x=-135470000;
#10;x=-135460000;
#10;x=-135450000;
#10;x=-135440000;
#10;x=-135430000;
#10;x=-135420000;
#10;x=-135410000;
#10;x=-135400000;
#10;x=-135390000;
#10;x=-135380000;
#10;x=-135370000;
#10;x=-135360000;
#10;x=-135350000;
#10;x=-135340000;
#10;x=-135330000;
#10;x=-135320000;
#10;x=-135310000;
#10;x=-135300000;
#10;x=-135290000;
#10;x=-135280000;
#10;x=-135270000;
#10;x=-135260000;
#10;x=-135250000;
#10;x=-135240000;
#10;x=-135230000;
#10;x=-135220000;
#10;x=-135210000;
#10;x=-135200000;
#10;x=-135190000;
#10;x=-135180000;
#10;x=-135170000;
#10;x=-135160000;
#10;x=-135150000;
#10;x=-135140000;
#10;x=-135130000;
#10;x=-135120000;
#10;x=-135110000;
#10;x=-135100000;
#10;x=-135090000;
#10;x=-135080000;
#10;x=-135070000;
#10;x=-135060000;
#10;x=-135050000;
#10;x=-135040000;
#10;x=-135030000;
#10;x=-135020000;
#10;x=-135010000;
#10;x=-135000000;
#10;x=-134990000;
#10;x=-134980000;
#10;x=-134970000;
#10;x=-134960000;
#10;x=-134950000;
#10;x=-134940000;
#10;x=-134930000;
#10;x=-134920000;
#10;x=-134910000;
#10;x=-134900000;
#10;x=-134890000;
#10;x=-134880000;
#10;x=-134870000;
#10;x=-134860000;
#10;x=-134850000;
#10;x=-134840000;
#10;x=-134830000;
#10;x=-134820000;
#10;x=-134810000;
#10;x=-134800000;
#10;x=-134790000;
#10;x=-134780000;
#10;x=-134770000;
#10;x=-134760000;
#10;x=-134750000;
#10;x=-134740000;
#10;x=-134730000;
#10;x=-134720000;
#10;x=-134710000;
#10;x=-134700000;
#10;x=-134690000;
#10;x=-134680000;
#10;x=-134670000;
#10;x=-134660000;
#10;x=-134650000;
#10;x=-134640000;
#10;x=-134630000;
#10;x=-134620000;
#10;x=-134610000;
#10;x=-134600000;
#10;x=-134590000;
#10;x=-134580000;
#10;x=-134570000;
#10;x=-134560000;
#10;x=-134550000;
#10;x=-134540000;
#10;x=-134530000;
#10;x=-134520000;
#10;x=-134510000;
#10;x=-134500000;
#10;x=-134490000;
#10;x=-134480000;
#10;x=-134470000;
#10;x=-134460000;
#10;x=-134450000;
#10;x=-134440000;
#10;x=-134430000;
#10;x=-134420000;
#10;x=-134410000;
#10;x=-134400000;
#10;x=-134390000;
#10;x=-134380000;
#10;x=-134370000;
#10;x=-134360000;
#10;x=-134350000;
#10;x=-134340000;
#10;x=-134330000;
#10;x=-134320000;
#10;x=-134310000;
#10;x=-134300000;
#10;x=-134290000;
#10;x=-134280000;
#10;x=-134270000;
#10;x=-134260000;
#10;x=-134250000;
#10;x=-134240000;
#10;x=-134230000;
#10;x=-134220000;
#10;x=-134210000;
#10;x=-134200000;
#10;x=-134190000;
#10;x=-134180000;
#10;x=-134170000;
#10;x=-134160000;
#10;x=-134150000;
#10;x=-134140000;
#10;x=-134130000;
#10;x=-134120000;
#10;x=-134110000;
#10;x=-134100000;
#10;x=-134090000;
#10;x=-134080000;
#10;x=-134070000;
#10;x=-134060000;
#10;x=-134050000;
#10;x=-134040000;
#10;x=-134030000;
#10;x=-134020000;
#10;x=-134010000;
#10;x=-134000000;
#10;x=-133990000;
#10;x=-133980000;
#10;x=-133970000;
#10;x=-133960000;
#10;x=-133950000;
#10;x=-133940000;
#10;x=-133930000;
#10;x=-133920000;
#10;x=-133910000;
#10;x=-133900000;
#10;x=-133890000;
#10;x=-133880000;
#10;x=-133870000;
#10;x=-133860000;
#10;x=-133850000;
#10;x=-133840000;
#10;x=-133830000;
#10;x=-133820000;
#10;x=-133810000;
#10;x=-133800000;
#10;x=-133790000;
#10;x=-133780000;
#10;x=-133770000;
#10;x=-133760000;
#10;x=-133750000;
#10;x=-133740000;
#10;x=-133730000;
#10;x=-133720000;
#10;x=-133710000;
#10;x=-133700000;
#10;x=-133690000;
#10;x=-133680000;
#10;x=-133670000;
#10;x=-133660000;
#10;x=-133650000;
#10;x=-133640000;
#10;x=-133630000;
#10;x=-133620000;
#10;x=-133610000;
#10;x=-133600000;
#10;x=-133590000;
#10;x=-133580000;
#10;x=-133570000;
#10;x=-133560000;
#10;x=-133550000;
#10;x=-133540000;
#10;x=-133530000;
#10;x=-133520000;
#10;x=-133510000;
#10;x=-133500000;
#10;x=-133490000;
#10;x=-133480000;
#10;x=-133470000;
#10;x=-133460000;
#10;x=-133450000;
#10;x=-133440000;
#10;x=-133430000;
#10;x=-133420000;
#10;x=-133410000;
#10;x=-133400000;
#10;x=-133390000;
#10;x=-133380000;
#10;x=-133370000;
#10;x=-133360000;
#10;x=-133350000;
#10;x=-133340000;
#10;x=-133330000;
#10;x=-133320000;
#10;x=-133310000;
#10;x=-133300000;
#10;x=-133290000;
#10;x=-133280000;
#10;x=-133270000;
#10;x=-133260000;
#10;x=-133250000;
#10;x=-133240000;
#10;x=-133230000;
#10;x=-133220000;
#10;x=-133210000;
#10;x=-133200000;
#10;x=-133190000;
#10;x=-133180000;
#10;x=-133170000;
#10;x=-133160000;
#10;x=-133150000;
#10;x=-133140000;
#10;x=-133130000;
#10;x=-133120000;
#10;x=-133110000;
#10;x=-133100000;
#10;x=-133090000;
#10;x=-133080000;
#10;x=-133070000;
#10;x=-133060000;
#10;x=-133050000;
#10;x=-133040000;
#10;x=-133030000;
#10;x=-133020000;
#10;x=-133010000;
#10;x=-133000000;
#10;x=-132990000;
#10;x=-132980000;
#10;x=-132970000;
#10;x=-132960000;
#10;x=-132950000;
#10;x=-132940000;
#10;x=-132930000;
#10;x=-132920000;
#10;x=-132910000;
#10;x=-132900000;
#10;x=-132890000;
#10;x=-132880000;
#10;x=-132870000;
#10;x=-132860000;
#10;x=-132850000;
#10;x=-132840000;
#10;x=-132830000;
#10;x=-132820000;
#10;x=-132810000;
#10;x=-132800000;
#10;x=-132790000;
#10;x=-132780000;
#10;x=-132770000;
#10;x=-132760000;
#10;x=-132750000;
#10;x=-132740000;
#10;x=-132730000;
#10;x=-132720000;
#10;x=-132710000;
#10;x=-132700000;
#10;x=-132690000;
#10;x=-132680000;
#10;x=-132670000;
#10;x=-132660000;
#10;x=-132650000;
#10;x=-132640000;
#10;x=-132630000;
#10;x=-132620000;
#10;x=-132610000;
#10;x=-132600000;
#10;x=-132590000;
#10;x=-132580000;
#10;x=-132570000;
#10;x=-132560000;
#10;x=-132550000;
#10;x=-132540000;
#10;x=-132530000;
#10;x=-132520000;
#10;x=-132510000;
#10;x=-132500000;
#10;x=-132490000;
#10;x=-132480000;
#10;x=-132470000;
#10;x=-132460000;
#10;x=-132450000;
#10;x=-132440000;
#10;x=-132430000;
#10;x=-132420000;
#10;x=-132410000;
#10;x=-132400000;
#10;x=-132390000;
#10;x=-132380000;
#10;x=-132370000;
#10;x=-132360000;
#10;x=-132350000;
#10;x=-132340000;
#10;x=-132330000;
#10;x=-132320000;
#10;x=-132310000;
#10;x=-132300000;
#10;x=-132290000;
#10;x=-132280000;
#10;x=-132270000;
#10;x=-132260000;
#10;x=-132250000;
#10;x=-132240000;
#10;x=-132230000;
#10;x=-132220000;
#10;x=-132210000;
#10;x=-132200000;
#10;x=-132190000;
#10;x=-132180000;
#10;x=-132170000;
#10;x=-132160000;
#10;x=-132150000;
#10;x=-132140000;
#10;x=-132130000;
#10;x=-132120000;
#10;x=-132110000;
#10;x=-132100000;
#10;x=-132090000;
#10;x=-132080000;
#10;x=-132070000;
#10;x=-132060000;
#10;x=-132050000;
#10;x=-132040000;
#10;x=-132030000;
#10;x=-132020000;
#10;x=-132010000;
#10;x=-132000000;
#10;x=-131990000;
#10;x=-131980000;
#10;x=-131970000;
#10;x=-131960000;
#10;x=-131950000;
#10;x=-131940000;
#10;x=-131930000;
#10;x=-131920000;
#10;x=-131910000;
#10;x=-131900000;
#10;x=-131890000;
#10;x=-131880000;
#10;x=-131870000;
#10;x=-131860000;
#10;x=-131850000;
#10;x=-131840000;
#10;x=-131830000;
#10;x=-131820000;
#10;x=-131810000;
#10;x=-131800000;
#10;x=-131790000;
#10;x=-131780000;
#10;x=-131770000;
#10;x=-131760000;
#10;x=-131750000;
#10;x=-131740000;
#10;x=-131730000;
#10;x=-131720000;
#10;x=-131710000;
#10;x=-131700000;
#10;x=-131690000;
#10;x=-131680000;
#10;x=-131670000;
#10;x=-131660000;
#10;x=-131650000;
#10;x=-131640000;
#10;x=-131630000;
#10;x=-131620000;
#10;x=-131610000;
#10;x=-131600000;
#10;x=-131590000;
#10;x=-131580000;
#10;x=-131570000;
#10;x=-131560000;
#10;x=-131550000;
#10;x=-131540000;
#10;x=-131530000;
#10;x=-131520000;
#10;x=-131510000;
#10;x=-131500000;
#10;x=-131490000;
#10;x=-131480000;
#10;x=-131470000;
#10;x=-131460000;
#10;x=-131450000;
#10;x=-131440000;
#10;x=-131430000;
#10;x=-131420000;
#10;x=-131410000;
#10;x=-131400000;
#10;x=-131390000;
#10;x=-131380000;
#10;x=-131370000;
#10;x=-131360000;
#10;x=-131350000;
#10;x=-131340000;
#10;x=-131330000;
#10;x=-131320000;
#10;x=-131310000;
#10;x=-131300000;
#10;x=-131290000;
#10;x=-131280000;
#10;x=-131270000;
#10;x=-131260000;
#10;x=-131250000;
#10;x=-131240000;
#10;x=-131230000;
#10;x=-131220000;
#10;x=-131210000;
#10;x=-131200000;
#10;x=-131190000;
#10;x=-131180000;
#10;x=-131170000;
#10;x=-131160000;
#10;x=-131150000;
#10;x=-131140000;
#10;x=-131130000;
#10;x=-131120000;
#10;x=-131110000;
#10;x=-131100000;
#10;x=-131090000;
#10;x=-131080000;
#10;x=-131070000;
#10;x=-131060000;
#10;x=-131050000;
#10;x=-131040000;
#10;x=-131030000;
#10;x=-131020000;
#10;x=-131010000;
#10;x=-131000000;
#10;x=-130990000;
#10;x=-130980000;
#10;x=-130970000;
#10;x=-130960000;
#10;x=-130950000;
#10;x=-130940000;
#10;x=-130930000;
#10;x=-130920000;
#10;x=-130910000;
#10;x=-130900000;
#10;x=-130890000;
#10;x=-130880000;
#10;x=-130870000;
#10;x=-130860000;
#10;x=-130850000;
#10;x=-130840000;
#10;x=-130830000;
#10;x=-130820000;
#10;x=-130810000;
#10;x=-130800000;
#10;x=-130790000;
#10;x=-130780000;
#10;x=-130770000;
#10;x=-130760000;
#10;x=-130750000;
#10;x=-130740000;
#10;x=-130730000;
#10;x=-130720000;
#10;x=-130710000;
#10;x=-130700000;
#10;x=-130690000;
#10;x=-130680000;
#10;x=-130670000;
#10;x=-130660000;
#10;x=-130650000;
#10;x=-130640000;
#10;x=-130630000;
#10;x=-130620000;
#10;x=-130610000;
#10;x=-130600000;
#10;x=-130590000;
#10;x=-130580000;
#10;x=-130570000;
#10;x=-130560000;
#10;x=-130550000;
#10;x=-130540000;
#10;x=-130530000;
#10;x=-130520000;
#10;x=-130510000;
#10;x=-130500000;
#10;x=-130490000;
#10;x=-130480000;
#10;x=-130470000;
#10;x=-130460000;
#10;x=-130450000;
#10;x=-130440000;
#10;x=-130430000;
#10;x=-130420000;
#10;x=-130410000;
#10;x=-130400000;
#10;x=-130390000;
#10;x=-130380000;
#10;x=-130370000;
#10;x=-130360000;
#10;x=-130350000;
#10;x=-130340000;
#10;x=-130330000;
#10;x=-130320000;
#10;x=-130310000;
#10;x=-130300000;
#10;x=-130290000;
#10;x=-130280000;
#10;x=-130270000;
#10;x=-130260000;
#10;x=-130250000;
#10;x=-130240000;
#10;x=-130230000;
#10;x=-130220000;
#10;x=-130210000;
#10;x=-130200000;
#10;x=-130190000;
#10;x=-130180000;
#10;x=-130170000;
#10;x=-130160000;
#10;x=-130150000;
#10;x=-130140000;
#10;x=-130130000;
#10;x=-130120000;
#10;x=-130110000;
#10;x=-130100000;
#10;x=-130090000;
#10;x=-130080000;
#10;x=-130070000;
#10;x=-130060000;
#10;x=-130050000;
#10;x=-130040000;
#10;x=-130030000;
#10;x=-130020000;
#10;x=-130010000;
#10;x=-130000000;
#10;x=-129990000;
#10;x=-129980000;
#10;x=-129970000;
#10;x=-129960000;
#10;x=-129950000;
#10;x=-129940000;
#10;x=-129930000;
#10;x=-129920000;
#10;x=-129910000;
#10;x=-129900000;
#10;x=-129890000;
#10;x=-129880000;
#10;x=-129870000;
#10;x=-129860000;
#10;x=-129850000;
#10;x=-129840000;
#10;x=-129830000;
#10;x=-129820000;
#10;x=-129810000;
#10;x=-129800000;
#10;x=-129790000;
#10;x=-129780000;
#10;x=-129770000;
#10;x=-129760000;
#10;x=-129750000;
#10;x=-129740000;
#10;x=-129730000;
#10;x=-129720000;
#10;x=-129710000;
#10;x=-129700000;
#10;x=-129690000;
#10;x=-129680000;
#10;x=-129670000;
#10;x=-129660000;
#10;x=-129650000;
#10;x=-129640000;
#10;x=-129630000;
#10;x=-129620000;
#10;x=-129610000;
#10;x=-129600000;
#10;x=-129590000;
#10;x=-129580000;
#10;x=-129570000;
#10;x=-129560000;
#10;x=-129550000;
#10;x=-129540000;
#10;x=-129530000;
#10;x=-129520000;
#10;x=-129510000;
#10;x=-129500000;
#10;x=-129490000;
#10;x=-129480000;
#10;x=-129470000;
#10;x=-129460000;
#10;x=-129450000;
#10;x=-129440000;
#10;x=-129430000;
#10;x=-129420000;
#10;x=-129410000;
#10;x=-129400000;
#10;x=-129390000;
#10;x=-129380000;
#10;x=-129370000;
#10;x=-129360000;
#10;x=-129350000;
#10;x=-129340000;
#10;x=-129330000;
#10;x=-129320000;
#10;x=-129310000;
#10;x=-129300000;
#10;x=-129290000;
#10;x=-129280000;
#10;x=-129270000;
#10;x=-129260000;
#10;x=-129250000;
#10;x=-129240000;
#10;x=-129230000;
#10;x=-129220000;
#10;x=-129210000;
#10;x=-129200000;
#10;x=-129190000;
#10;x=-129180000;
#10;x=-129170000;
#10;x=-129160000;
#10;x=-129150000;
#10;x=-129140000;
#10;x=-129130000;
#10;x=-129120000;
#10;x=-129110000;
#10;x=-129100000;
#10;x=-129090000;
#10;x=-129080000;
#10;x=-129070000;
#10;x=-129060000;
#10;x=-129050000;
#10;x=-129040000;
#10;x=-129030000;
#10;x=-129020000;
#10;x=-129010000;
#10;x=-129000000;
#10;x=-128990000;
#10;x=-128980000;
#10;x=-128970000;
#10;x=-128960000;
#10;x=-128950000;
#10;x=-128940000;
#10;x=-128930000;
#10;x=-128920000;
#10;x=-128910000;
#10;x=-128900000;
#10;x=-128890000;
#10;x=-128880000;
#10;x=-128870000;
#10;x=-128860000;
#10;x=-128850000;
#10;x=-128840000;
#10;x=-128830000;
#10;x=-128820000;
#10;x=-128810000;
#10;x=-128800000;
#10;x=-128790000;
#10;x=-128780000;
#10;x=-128770000;
#10;x=-128760000;
#10;x=-128750000;
#10;x=-128740000;
#10;x=-128730000;
#10;x=-128720000;
#10;x=-128710000;
#10;x=-128700000;
#10;x=-128690000;
#10;x=-128680000;
#10;x=-128670000;
#10;x=-128660000;
#10;x=-128650000;
#10;x=-128640000;
#10;x=-128630000;
#10;x=-128620000;
#10;x=-128610000;
#10;x=-128600000;
#10;x=-128590000;
#10;x=-128580000;
#10;x=-128570000;
#10;x=-128560000;
#10;x=-128550000;
#10;x=-128540000;
#10;x=-128530000;
#10;x=-128520000;
#10;x=-128510000;
#10;x=-128500000;
#10;x=-128490000;
#10;x=-128480000;
#10;x=-128470000;
#10;x=-128460000;
#10;x=-128450000;
#10;x=-128440000;
#10;x=-128430000;
#10;x=-128420000;
#10;x=-128410000;
#10;x=-128400000;
#10;x=-128390000;
#10;x=-128380000;
#10;x=-128370000;
#10;x=-128360000;
#10;x=-128350000;
#10;x=-128340000;
#10;x=-128330000;
#10;x=-128320000;
#10;x=-128310000;
#10;x=-128300000;
#10;x=-128290000;
#10;x=-128280000;
#10;x=-128270000;
#10;x=-128260000;
#10;x=-128250000;
#10;x=-128240000;
#10;x=-128230000;
#10;x=-128220000;
#10;x=-128210000;
#10;x=-128200000;
#10;x=-128190000;
#10;x=-128180000;
#10;x=-128170000;
#10;x=-128160000;
#10;x=-128150000;
#10;x=-128140000;
#10;x=-128130000;
#10;x=-128120000;
#10;x=-128110000;
#10;x=-128100000;
#10;x=-128090000;
#10;x=-128080000;
#10;x=-128070000;
#10;x=-128060000;
#10;x=-128050000;
#10;x=-128040000;
#10;x=-128030000;
#10;x=-128020000;
#10;x=-128010000;
#10;x=-128000000;
#10;x=-127990000;
#10;x=-127980000;
#10;x=-127970000;
#10;x=-127960000;
#10;x=-127950000;
#10;x=-127940000;
#10;x=-127930000;
#10;x=-127920000;
#10;x=-127910000;
#10;x=-127900000;
#10;x=-127890000;
#10;x=-127880000;
#10;x=-127870000;
#10;x=-127860000;
#10;x=-127850000;
#10;x=-127840000;
#10;x=-127830000;
#10;x=-127820000;
#10;x=-127810000;
#10;x=-127800000;
#10;x=-127790000;
#10;x=-127780000;
#10;x=-127770000;
#10;x=-127760000;
#10;x=-127750000;
#10;x=-127740000;
#10;x=-127730000;
#10;x=-127720000;
#10;x=-127710000;
#10;x=-127700000;
#10;x=-127690000;
#10;x=-127680000;
#10;x=-127670000;
#10;x=-127660000;
#10;x=-127650000;
#10;x=-127640000;
#10;x=-127630000;
#10;x=-127620000;
#10;x=-127610000;
#10;x=-127600000;
#10;x=-127590000;
#10;x=-127580000;
#10;x=-127570000;
#10;x=-127560000;
#10;x=-127550000;
#10;x=-127540000;
#10;x=-127530000;
#10;x=-127520000;
#10;x=-127510000;
#10;x=-127500000;
#10;x=-127490000;
#10;x=-127480000;
#10;x=-127470000;
#10;x=-127460000;
#10;x=-127450000;
#10;x=-127440000;
#10;x=-127430000;
#10;x=-127420000;
#10;x=-127410000;
#10;x=-127400000;
#10;x=-127390000;
#10;x=-127380000;
#10;x=-127370000;
#10;x=-127360000;
#10;x=-127350000;
#10;x=-127340000;
#10;x=-127330000;
#10;x=-127320000;
#10;x=-127310000;
#10;x=-127300000;
#10;x=-127290000;
#10;x=-127280000;
#10;x=-127270000;
#10;x=-127260000;
#10;x=-127250000;
#10;x=-127240000;
#10;x=-127230000;
#10;x=-127220000;
#10;x=-127210000;
#10;x=-127200000;
#10;x=-127190000;
#10;x=-127180000;
#10;x=-127170000;
#10;x=-127160000;
#10;x=-127150000;
#10;x=-127140000;
#10;x=-127130000;
#10;x=-127120000;
#10;x=-127110000;
#10;x=-127100000;
#10;x=-127090000;
#10;x=-127080000;
#10;x=-127070000;
#10;x=-127060000;
#10;x=-127050000;
#10;x=-127040000;
#10;x=-127030000;
#10;x=-127020000;
#10;x=-127010000;
#10;x=-127000000;
#10;x=-126990000;
#10;x=-126980000;
#10;x=-126970000;
#10;x=-126960000;
#10;x=-126950000;
#10;x=-126940000;
#10;x=-126930000;
#10;x=-126920000;
#10;x=-126910000;
#10;x=-126900000;
#10;x=-126890000;
#10;x=-126880000;
#10;x=-126870000;
#10;x=-126860000;
#10;x=-126850000;
#10;x=-126840000;
#10;x=-126830000;
#10;x=-126820000;
#10;x=-126810000;
#10;x=-126800000;
#10;x=-126790000;
#10;x=-126780000;
#10;x=-126770000;
#10;x=-126760000;
#10;x=-126750000;
#10;x=-126740000;
#10;x=-126730000;
#10;x=-126720000;
#10;x=-126710000;
#10;x=-126700000;
#10;x=-126690000;
#10;x=-126680000;
#10;x=-126670000;
#10;x=-126660000;
#10;x=-126650000;
#10;x=-126640000;
#10;x=-126630000;
#10;x=-126620000;
#10;x=-126610000;
#10;x=-126600000;
#10;x=-126590000;
#10;x=-126580000;
#10;x=-126570000;
#10;x=-126560000;
#10;x=-126550000;
#10;x=-126540000;
#10;x=-126530000;
#10;x=-126520000;
#10;x=-126510000;
#10;x=-126500000;
#10;x=-126490000;
#10;x=-126480000;
#10;x=-126470000;
#10;x=-126460000;
#10;x=-126450000;
#10;x=-126440000;
#10;x=-126430000;
#10;x=-126420000;
#10;x=-126410000;
#10;x=-126400000;
#10;x=-126390000;
#10;x=-126380000;
#10;x=-126370000;
#10;x=-126360000;
#10;x=-126350000;
#10;x=-126340000;
#10;x=-126330000;
#10;x=-126320000;
#10;x=-126310000;
#10;x=-126300000;
#10;x=-126290000;
#10;x=-126280000;
#10;x=-126270000;
#10;x=-126260000;
#10;x=-126250000;
#10;x=-126240000;
#10;x=-126230000;
#10;x=-126220000;
#10;x=-126210000;
#10;x=-126200000;
#10;x=-126190000;
#10;x=-126180000;
#10;x=-126170000;
#10;x=-126160000;
#10;x=-126150000;
#10;x=-126140000;
#10;x=-126130000;
#10;x=-126120000;
#10;x=-126110000;
#10;x=-126100000;
#10;x=-126090000;
#10;x=-126080000;
#10;x=-126070000;
#10;x=-126060000;
#10;x=-126050000;
#10;x=-126040000;
#10;x=-126030000;
#10;x=-126020000;
#10;x=-126010000;
#10;x=-126000000;
#10;x=-125990000;
#10;x=-125980000;
#10;x=-125970000;
#10;x=-125960000;
#10;x=-125950000;
#10;x=-125940000;
#10;x=-125930000;
#10;x=-125920000;
#10;x=-125910000;
#10;x=-125900000;
#10;x=-125890000;
#10;x=-125880000;
#10;x=-125870000;
#10;x=-125860000;
#10;x=-125850000;
#10;x=-125840000;
#10;x=-125830000;
#10;x=-125820000;
#10;x=-125810000;
#10;x=-125800000;
#10;x=-125790000;
#10;x=-125780000;
#10;x=-125770000;
#10;x=-125760000;
#10;x=-125750000;
#10;x=-125740000;
#10;x=-125730000;
#10;x=-125720000;
#10;x=-125710000;
#10;x=-125700000;
#10;x=-125690000;
#10;x=-125680000;
#10;x=-125670000;
#10;x=-125660000;
#10;x=-125650000;
#10;x=-125640000;
#10;x=-125630000;
#10;x=-125620000;
#10;x=-125610000;
#10;x=-125600000;
#10;x=-125590000;
#10;x=-125580000;
#10;x=-125570000;
#10;x=-125560000;
#10;x=-125550000;
#10;x=-125540000;
#10;x=-125530000;
#10;x=-125520000;
#10;x=-125510000;
#10;x=-125500000;
#10;x=-125490000;
#10;x=-125480000;
#10;x=-125470000;
#10;x=-125460000;
#10;x=-125450000;
#10;x=-125440000;
#10;x=-125430000;
#10;x=-125420000;
#10;x=-125410000;
#10;x=-125400000;
#10;x=-125390000;
#10;x=-125380000;
#10;x=-125370000;
#10;x=-125360000;
#10;x=-125350000;
#10;x=-125340000;
#10;x=-125330000;
#10;x=-125320000;
#10;x=-125310000;
#10;x=-125300000;
#10;x=-125290000;
#10;x=-125280000;
#10;x=-125270000;
#10;x=-125260000;
#10;x=-125250000;
#10;x=-125240000;
#10;x=-125230000;
#10;x=-125220000;
#10;x=-125210000;
#10;x=-125200000;
#10;x=-125190000;
#10;x=-125180000;
#10;x=-125170000;
#10;x=-125160000;
#10;x=-125150000;
#10;x=-125140000;
#10;x=-125130000;
#10;x=-125120000;
#10;x=-125110000;
#10;x=-125100000;
#10;x=-125090000;
#10;x=-125080000;
#10;x=-125070000;
#10;x=-125060000;
#10;x=-125050000;
#10;x=-125040000;
#10;x=-125030000;
#10;x=-125020000;
#10;x=-125010000;
#10;x=-125000000;
#10;x=-124990000;
#10;x=-124980000;
#10;x=-124970000;
#10;x=-124960000;
#10;x=-124950000;
#10;x=-124940000;
#10;x=-124930000;
#10;x=-124920000;
#10;x=-124910000;
#10;x=-124900000;
#10;x=-124890000;
#10;x=-124880000;
#10;x=-124870000;
#10;x=-124860000;
#10;x=-124850000;
#10;x=-124840000;
#10;x=-124830000;
#10;x=-124820000;
#10;x=-124810000;
#10;x=-124800000;
#10;x=-124790000;
#10;x=-124780000;
#10;x=-124770000;
#10;x=-124760000;
#10;x=-124750000;
#10;x=-124740000;
#10;x=-124730000;
#10;x=-124720000;
#10;x=-124710000;
#10;x=-124700000;
#10;x=-124690000;
#10;x=-124680000;
#10;x=-124670000;
#10;x=-124660000;
#10;x=-124650000;
#10;x=-124640000;
#10;x=-124630000;
#10;x=-124620000;
#10;x=-124610000;
#10;x=-124600000;
#10;x=-124590000;
#10;x=-124580000;
#10;x=-124570000;
#10;x=-124560000;
#10;x=-124550000;
#10;x=-124540000;
#10;x=-124530000;
#10;x=-124520000;
#10;x=-124510000;
#10;x=-124500000;
#10;x=-124490000;
#10;x=-124480000;
#10;x=-124470000;
#10;x=-124460000;
#10;x=-124450000;
#10;x=-124440000;
#10;x=-124430000;
#10;x=-124420000;
#10;x=-124410000;
#10;x=-124400000;
#10;x=-124390000;
#10;x=-124380000;
#10;x=-124370000;
#10;x=-124360000;
#10;x=-124350000;
#10;x=-124340000;
#10;x=-124330000;
#10;x=-124320000;
#10;x=-124310000;
#10;x=-124300000;
#10;x=-124290000;
#10;x=-124280000;
#10;x=-124270000;
#10;x=-124260000;
#10;x=-124250000;
#10;x=-124240000;
#10;x=-124230000;
#10;x=-124220000;
#10;x=-124210000;
#10;x=-124200000;
#10;x=-124190000;
#10;x=-124180000;
#10;x=-124170000;
#10;x=-124160000;
#10;x=-124150000;
#10;x=-124140000;
#10;x=-124130000;
#10;x=-124120000;
#10;x=-124110000;
#10;x=-124100000;
#10;x=-124090000;
#10;x=-124080000;
#10;x=-124070000;
#10;x=-124060000;
#10;x=-124050000;
#10;x=-124040000;
#10;x=-124030000;
#10;x=-124020000;
#10;x=-124010000;
#10;x=-124000000;
#10;x=-123990000;
#10;x=-123980000;
#10;x=-123970000;
#10;x=-123960000;
#10;x=-123950000;
#10;x=-123940000;
#10;x=-123930000;
#10;x=-123920000;
#10;x=-123910000;
#10;x=-123900000;
#10;x=-123890000;
#10;x=-123880000;
#10;x=-123870000;
#10;x=-123860000;
#10;x=-123850000;
#10;x=-123840000;
#10;x=-123830000;
#10;x=-123820000;
#10;x=-123810000;
#10;x=-123800000;
#10;x=-123790000;
#10;x=-123780000;
#10;x=-123770000;
#10;x=-123760000;
#10;x=-123750000;
#10;x=-123740000;
#10;x=-123730000;
#10;x=-123720000;
#10;x=-123710000;
#10;x=-123700000;
#10;x=-123690000;
#10;x=-123680000;
#10;x=-123670000;
#10;x=-123660000;
#10;x=-123650000;
#10;x=-123640000;
#10;x=-123630000;
#10;x=-123620000;
#10;x=-123610000;
#10;x=-123600000;
#10;x=-123590000;
#10;x=-123580000;
#10;x=-123570000;
#10;x=-123560000;
#10;x=-123550000;
#10;x=-123540000;
#10;x=-123530000;
#10;x=-123520000;
#10;x=-123510000;
#10;x=-123500000;
#10;x=-123490000;
#10;x=-123480000;
#10;x=-123470000;
#10;x=-123460000;
#10;x=-123450000;
#10;x=-123440000;
#10;x=-123430000;
#10;x=-123420000;
#10;x=-123410000;
#10;x=-123400000;
#10;x=-123390000;
#10;x=-123380000;
#10;x=-123370000;
#10;x=-123360000;
#10;x=-123350000;
#10;x=-123340000;
#10;x=-123330000;
#10;x=-123320000;
#10;x=-123310000;
#10;x=-123300000;
#10;x=-123290000;
#10;x=-123280000;
#10;x=-123270000;
#10;x=-123260000;
#10;x=-123250000;
#10;x=-123240000;
#10;x=-123230000;
#10;x=-123220000;
#10;x=-123210000;
#10;x=-123200000;
#10;x=-123190000;
#10;x=-123180000;
#10;x=-123170000;
#10;x=-123160000;
#10;x=-123150000;
#10;x=-123140000;
#10;x=-123130000;
#10;x=-123120000;
#10;x=-123110000;
#10;x=-123100000;
#10;x=-123090000;
#10;x=-123080000;
#10;x=-123070000;
#10;x=-123060000;
#10;x=-123050000;
#10;x=-123040000;
#10;x=-123030000;
#10;x=-123020000;
#10;x=-123010000;
#10;x=-123000000;
#10;x=-122990000;
#10;x=-122980000;
#10;x=-122970000;
#10;x=-122960000;
#10;x=-122950000;
#10;x=-122940000;
#10;x=-122930000;
#10;x=-122920000;
#10;x=-122910000;
#10;x=-122900000;
#10;x=-122890000;
#10;x=-122880000;
#10;x=-122870000;
#10;x=-122860000;
#10;x=-122850000;
#10;x=-122840000;
#10;x=-122830000;
#10;x=-122820000;
#10;x=-122810000;
#10;x=-122800000;
#10;x=-122790000;
#10;x=-122780000;
#10;x=-122770000;
#10;x=-122760000;
#10;x=-122750000;
#10;x=-122740000;
#10;x=-122730000;
#10;x=-122720000;
#10;x=-122710000;
#10;x=-122700000;
#10;x=-122690000;
#10;x=-122680000;
#10;x=-122670000;
#10;x=-122660000;
#10;x=-122650000;
#10;x=-122640000;
#10;x=-122630000;
#10;x=-122620000;
#10;x=-122610000;
#10;x=-122600000;
#10;x=-122590000;
#10;x=-122580000;
#10;x=-122570000;
#10;x=-122560000;
#10;x=-122550000;
#10;x=-122540000;
#10;x=-122530000;
#10;x=-122520000;
#10;x=-122510000;
#10;x=-122500000;
#10;x=-122490000;
#10;x=-122480000;
#10;x=-122470000;
#10;x=-122460000;
#10;x=-122450000;
#10;x=-122440000;
#10;x=-122430000;
#10;x=-122420000;
#10;x=-122410000;
#10;x=-122400000;
#10;x=-122390000;
#10;x=-122380000;
#10;x=-122370000;
#10;x=-122360000;
#10;x=-122350000;
#10;x=-122340000;
#10;x=-122330000;
#10;x=-122320000;
#10;x=-122310000;
#10;x=-122300000;
#10;x=-122290000;
#10;x=-122280000;
#10;x=-122270000;
#10;x=-122260000;
#10;x=-122250000;
#10;x=-122240000;
#10;x=-122230000;
#10;x=-122220000;
#10;x=-122210000;
#10;x=-122200000;
#10;x=-122190000;
#10;x=-122180000;
#10;x=-122170000;
#10;x=-122160000;
#10;x=-122150000;
#10;x=-122140000;
#10;x=-122130000;
#10;x=-122120000;
#10;x=-122110000;
#10;x=-122100000;
#10;x=-122090000;
#10;x=-122080000;
#10;x=-122070000;
#10;x=-122060000;
#10;x=-122050000;
#10;x=-122040000;
#10;x=-122030000;
#10;x=-122020000;
#10;x=-122010000;
#10;x=-122000000;
#10;x=-121990000;
#10;x=-121980000;
#10;x=-121970000;
#10;x=-121960000;
#10;x=-121950000;
#10;x=-121940000;
#10;x=-121930000;
#10;x=-121920000;
#10;x=-121910000;
#10;x=-121900000;
#10;x=-121890000;
#10;x=-121880000;
#10;x=-121870000;
#10;x=-121860000;
#10;x=-121850000;
#10;x=-121840000;
#10;x=-121830000;
#10;x=-121820000;
#10;x=-121810000;
#10;x=-121800000;
#10;x=-121790000;
#10;x=-121780000;
#10;x=-121770000;
#10;x=-121760000;
#10;x=-121750000;
#10;x=-121740000;
#10;x=-121730000;
#10;x=-121720000;
#10;x=-121710000;
#10;x=-121700000;
#10;x=-121690000;
#10;x=-121680000;
#10;x=-121670000;
#10;x=-121660000;
#10;x=-121650000;
#10;x=-121640000;
#10;x=-121630000;
#10;x=-121620000;
#10;x=-121610000;
#10;x=-121600000;
#10;x=-121590000;
#10;x=-121580000;
#10;x=-121570000;
#10;x=-121560000;
#10;x=-121550000;
#10;x=-121540000;
#10;x=-121530000;
#10;x=-121520000;
#10;x=-121510000;
#10;x=-121500000;
#10;x=-121490000;
#10;x=-121480000;
#10;x=-121470000;
#10;x=-121460000;
#10;x=-121450000;
#10;x=-121440000;
#10;x=-121430000;
#10;x=-121420000;
#10;x=-121410000;
#10;x=-121400000;
#10;x=-121390000;
#10;x=-121380000;
#10;x=-121370000;
#10;x=-121360000;
#10;x=-121350000;
#10;x=-121340000;
#10;x=-121330000;
#10;x=-121320000;
#10;x=-121310000;
#10;x=-121300000;
#10;x=-121290000;
#10;x=-121280000;
#10;x=-121270000;
#10;x=-121260000;
#10;x=-121250000;
#10;x=-121240000;
#10;x=-121230000;
#10;x=-121220000;
#10;x=-121210000;
#10;x=-121200000;
#10;x=-121190000;
#10;x=-121180000;
#10;x=-121170000;
#10;x=-121160000;
#10;x=-121150000;
#10;x=-121140000;
#10;x=-121130000;
#10;x=-121120000;
#10;x=-121110000;
#10;x=-121100000;
#10;x=-121090000;
#10;x=-121080000;
#10;x=-121070000;
#10;x=-121060000;
#10;x=-121050000;
#10;x=-121040000;
#10;x=-121030000;
#10;x=-121020000;
#10;x=-121010000;
#10;x=-121000000;
#10;x=-120990000;
#10;x=-120980000;
#10;x=-120970000;
#10;x=-120960000;
#10;x=-120950000;
#10;x=-120940000;
#10;x=-120930000;
#10;x=-120920000;
#10;x=-120910000;
#10;x=-120900000;
#10;x=-120890000;
#10;x=-120880000;
#10;x=-120870000;
#10;x=-120860000;
#10;x=-120850000;
#10;x=-120840000;
#10;x=-120830000;
#10;x=-120820000;
#10;x=-120810000;
#10;x=-120800000;
#10;x=-120790000;
#10;x=-120780000;
#10;x=-120770000;
#10;x=-120760000;
#10;x=-120750000;
#10;x=-120740000;
#10;x=-120730000;
#10;x=-120720000;
#10;x=-120710000;
#10;x=-120700000;
#10;x=-120690000;
#10;x=-120680000;
#10;x=-120670000;
#10;x=-120660000;
#10;x=-120650000;
#10;x=-120640000;
#10;x=-120630000;
#10;x=-120620000;
#10;x=-120610000;
#10;x=-120600000;
#10;x=-120590000;
#10;x=-120580000;
#10;x=-120570000;
#10;x=-120560000;
#10;x=-120550000;
#10;x=-120540000;
#10;x=-120530000;
#10;x=-120520000;
#10;x=-120510000;
#10;x=-120500000;
#10;x=-120490000;
#10;x=-120480000;
#10;x=-120470000;
#10;x=-120460000;
#10;x=-120450000;
#10;x=-120440000;
#10;x=-120430000;
#10;x=-120420000;
#10;x=-120410000;
#10;x=-120400000;
#10;x=-120390000;
#10;x=-120380000;
#10;x=-120370000;
#10;x=-120360000;
#10;x=-120350000;
#10;x=-120340000;
#10;x=-120330000;
#10;x=-120320000;
#10;x=-120310000;
#10;x=-120300000;
#10;x=-120290000;
#10;x=-120280000;
#10;x=-120270000;
#10;x=-120260000;
#10;x=-120250000;
#10;x=-120240000;
#10;x=-120230000;
#10;x=-120220000;
#10;x=-120210000;
#10;x=-120200000;
#10;x=-120190000;
#10;x=-120180000;
#10;x=-120170000;
#10;x=-120160000;
#10;x=-120150000;
#10;x=-120140000;
#10;x=-120130000;
#10;x=-120120000;
#10;x=-120110000;
#10;x=-120100000;
#10;x=-120090000;
#10;x=-120080000;
#10;x=-120070000;
#10;x=-120060000;
#10;x=-120050000;
#10;x=-120040000;
#10;x=-120030000;
#10;x=-120020000;
#10;x=-120010000;
#10;x=-120000000;
#10;x=-119990000;
#10;x=-119980000;
#10;x=-119970000;
#10;x=-119960000;
#10;x=-119950000;
#10;x=-119940000;
#10;x=-119930000;
#10;x=-119920000;
#10;x=-119910000;
#10;x=-119900000;
#10;x=-119890000;
#10;x=-119880000;
#10;x=-119870000;
#10;x=-119860000;
#10;x=-119850000;
#10;x=-119840000;
#10;x=-119830000;
#10;x=-119820000;
#10;x=-119810000;
#10;x=-119800000;
#10;x=-119790000;
#10;x=-119780000;
#10;x=-119770000;
#10;x=-119760000;
#10;x=-119750000;
#10;x=-119740000;
#10;x=-119730000;
#10;x=-119720000;
#10;x=-119710000;
#10;x=-119700000;
#10;x=-119690000;
#10;x=-119680000;
#10;x=-119670000;
#10;x=-119660000;
#10;x=-119650000;
#10;x=-119640000;
#10;x=-119630000;
#10;x=-119620000;
#10;x=-119610000;
#10;x=-119600000;
#10;x=-119590000;
#10;x=-119580000;
#10;x=-119570000;
#10;x=-119560000;
#10;x=-119550000;
#10;x=-119540000;
#10;x=-119530000;
#10;x=-119520000;
#10;x=-119510000;
#10;x=-119500000;
#10;x=-119490000;
#10;x=-119480000;
#10;x=-119470000;
#10;x=-119460000;
#10;x=-119450000;
#10;x=-119440000;
#10;x=-119430000;
#10;x=-119420000;
#10;x=-119410000;
#10;x=-119400000;
#10;x=-119390000;
#10;x=-119380000;
#10;x=-119370000;
#10;x=-119360000;
#10;x=-119350000;
#10;x=-119340000;
#10;x=-119330000;
#10;x=-119320000;
#10;x=-119310000;
#10;x=-119300000;
#10;x=-119290000;
#10;x=-119280000;
#10;x=-119270000;
#10;x=-119260000;
#10;x=-119250000;
#10;x=-119240000;
#10;x=-119230000;
#10;x=-119220000;
#10;x=-119210000;
#10;x=-119200000;
#10;x=-119190000;
#10;x=-119180000;
#10;x=-119170000;
#10;x=-119160000;
#10;x=-119150000;
#10;x=-119140000;
#10;x=-119130000;
#10;x=-119120000;
#10;x=-119110000;
#10;x=-119100000;
#10;x=-119090000;
#10;x=-119080000;
#10;x=-119070000;
#10;x=-119060000;
#10;x=-119050000;
#10;x=-119040000;
#10;x=-119030000;
#10;x=-119020000;
#10;x=-119010000;
#10;x=-119000000;
#10;x=-118990000;
#10;x=-118980000;
#10;x=-118970000;
#10;x=-118960000;
#10;x=-118950000;
#10;x=-118940000;
#10;x=-118930000;
#10;x=-118920000;
#10;x=-118910000;
#10;x=-118900000;
#10;x=-118890000;
#10;x=-118880000;
#10;x=-118870000;
#10;x=-118860000;
#10;x=-118850000;
#10;x=-118840000;
#10;x=-118830000;
#10;x=-118820000;
#10;x=-118810000;
#10;x=-118800000;
#10;x=-118790000;
#10;x=-118780000;
#10;x=-118770000;
#10;x=-118760000;
#10;x=-118750000;
#10;x=-118740000;
#10;x=-118730000;
#10;x=-118720000;
#10;x=-118710000;
#10;x=-118700000;
#10;x=-118690000;
#10;x=-118680000;
#10;x=-118670000;
#10;x=-118660000;
#10;x=-118650000;
#10;x=-118640000;
#10;x=-118630000;
#10;x=-118620000;
#10;x=-118610000;
#10;x=-118600000;
#10;x=-118590000;
#10;x=-118580000;
#10;x=-118570000;
#10;x=-118560000;
#10;x=-118550000;
#10;x=-118540000;
#10;x=-118530000;
#10;x=-118520000;
#10;x=-118510000;
#10;x=-118500000;
#10;x=-118490000;
#10;x=-118480000;
#10;x=-118470000;
#10;x=-118460000;
#10;x=-118450000;
#10;x=-118440000;
#10;x=-118430000;
#10;x=-118420000;
#10;x=-118410000;
#10;x=-118400000;
#10;x=-118390000;
#10;x=-118380000;
#10;x=-118370000;
#10;x=-118360000;
#10;x=-118350000;
#10;x=-118340000;
#10;x=-118330000;
#10;x=-118320000;
#10;x=-118310000;
#10;x=-118300000;
#10;x=-118290000;
#10;x=-118280000;
#10;x=-118270000;
#10;x=-118260000;
#10;x=-118250000;
#10;x=-118240000;
#10;x=-118230000;
#10;x=-118220000;
#10;x=-118210000;
#10;x=-118200000;
#10;x=-118190000;
#10;x=-118180000;
#10;x=-118170000;
#10;x=-118160000;
#10;x=-118150000;
#10;x=-118140000;
#10;x=-118130000;
#10;x=-118120000;
#10;x=-118110000;
#10;x=-118100000;
#10;x=-118090000;
#10;x=-118080000;
#10;x=-118070000;
#10;x=-118060000;
#10;x=-118050000;
#10;x=-118040000;
#10;x=-118030000;
#10;x=-118020000;
#10;x=-118010000;
#10;x=-118000000;
#10;x=-117990000;
#10;x=-117980000;
#10;x=-117970000;
#10;x=-117960000;
#10;x=-117950000;
#10;x=-117940000;
#10;x=-117930000;
#10;x=-117920000;
#10;x=-117910000;
#10;x=-117900000;
#10;x=-117890000;
#10;x=-117880000;
#10;x=-117870000;
#10;x=-117860000;
#10;x=-117850000;
#10;x=-117840000;
#10;x=-117830000;
#10;x=-117820000;
#10;x=-117810000;
#10;x=-117800000;
#10;x=-117790000;
#10;x=-117780000;
#10;x=-117770000;
#10;x=-117760000;
#10;x=-117750000;
#10;x=-117740000;
#10;x=-117730000;
#10;x=-117720000;
#10;x=-117710000;
#10;x=-117700000;
#10;x=-117690000;
#10;x=-117680000;
#10;x=-117670000;
#10;x=-117660000;
#10;x=-117650000;
#10;x=-117640000;
#10;x=-117630000;
#10;x=-117620000;
#10;x=-117610000;
#10;x=-117600000;
#10;x=-117590000;
#10;x=-117580000;
#10;x=-117570000;
#10;x=-117560000;
#10;x=-117550000;
#10;x=-117540000;
#10;x=-117530000;
#10;x=-117520000;
#10;x=-117510000;
#10;x=-117500000;
#10;x=-117490000;
#10;x=-117480000;
#10;x=-117470000;
#10;x=-117460000;
#10;x=-117450000;
#10;x=-117440000;
#10;x=-117430000;
#10;x=-117420000;
#10;x=-117410000;
#10;x=-117400000;
#10;x=-117390000;
#10;x=-117380000;
#10;x=-117370000;
#10;x=-117360000;
#10;x=-117350000;
#10;x=-117340000;
#10;x=-117330000;
#10;x=-117320000;
#10;x=-117310000;
#10;x=-117300000;
#10;x=-117290000;
#10;x=-117280000;
#10;x=-117270000;
#10;x=-117260000;
#10;x=-117250000;
#10;x=-117240000;
#10;x=-117230000;
#10;x=-117220000;
#10;x=-117210000;
#10;x=-117200000;
#10;x=-117190000;
#10;x=-117180000;
#10;x=-117170000;
#10;x=-117160000;
#10;x=-117150000;
#10;x=-117140000;
#10;x=-117130000;
#10;x=-117120000;
#10;x=-117110000;
#10;x=-117100000;
#10;x=-117090000;
#10;x=-117080000;
#10;x=-117070000;
#10;x=-117060000;
#10;x=-117050000;
#10;x=-117040000;
#10;x=-117030000;
#10;x=-117020000;
#10;x=-117010000;
#10;x=-117000000;
#10;x=-116990000;
#10;x=-116980000;
#10;x=-116970000;
#10;x=-116960000;
#10;x=-116950000;
#10;x=-116940000;
#10;x=-116930000;
#10;x=-116920000;
#10;x=-116910000;
#10;x=-116900000;
#10;x=-116890000;
#10;x=-116880000;
#10;x=-116870000;
#10;x=-116860000;
#10;x=-116850000;
#10;x=-116840000;
#10;x=-116830000;
#10;x=-116820000;
#10;x=-116810000;
#10;x=-116800000;
#10;x=-116790000;
#10;x=-116780000;
#10;x=-116770000;
#10;x=-116760000;
#10;x=-116750000;
#10;x=-116740000;
#10;x=-116730000;
#10;x=-116720000;
#10;x=-116710000;
#10;x=-116700000;
#10;x=-116690000;
#10;x=-116680000;
#10;x=-116670000;
#10;x=-116660000;
#10;x=-116650000;
#10;x=-116640000;
#10;x=-116630000;
#10;x=-116620000;
#10;x=-116610000;
#10;x=-116600000;
#10;x=-116590000;
#10;x=-116580000;
#10;x=-116570000;
#10;x=-116560000;
#10;x=-116550000;
#10;x=-116540000;
#10;x=-116530000;
#10;x=-116520000;
#10;x=-116510000;
#10;x=-116500000;
#10;x=-116490000;
#10;x=-116480000;
#10;x=-116470000;
#10;x=-116460000;
#10;x=-116450000;
#10;x=-116440000;
#10;x=-116430000;
#10;x=-116420000;
#10;x=-116410000;
#10;x=-116400000;
#10;x=-116390000;
#10;x=-116380000;
#10;x=-116370000;
#10;x=-116360000;
#10;x=-116350000;
#10;x=-116340000;
#10;x=-116330000;
#10;x=-116320000;
#10;x=-116310000;
#10;x=-116300000;
#10;x=-116290000;
#10;x=-116280000;
#10;x=-116270000;
#10;x=-116260000;
#10;x=-116250000;
#10;x=-116240000;
#10;x=-116230000;
#10;x=-116220000;
#10;x=-116210000;
#10;x=-116200000;
#10;x=-116190000;
#10;x=-116180000;
#10;x=-116170000;
#10;x=-116160000;
#10;x=-116150000;
#10;x=-116140000;
#10;x=-116130000;
#10;x=-116120000;
#10;x=-116110000;
#10;x=-116100000;
#10;x=-116090000;
#10;x=-116080000;
#10;x=-116070000;
#10;x=-116060000;
#10;x=-116050000;
#10;x=-116040000;
#10;x=-116030000;
#10;x=-116020000;
#10;x=-116010000;
#10;x=-116000000;
#10;x=-115990000;
#10;x=-115980000;
#10;x=-115970000;
#10;x=-115960000;
#10;x=-115950000;
#10;x=-115940000;
#10;x=-115930000;
#10;x=-115920000;
#10;x=-115910000;
#10;x=-115900000;
#10;x=-115890000;
#10;x=-115880000;
#10;x=-115870000;
#10;x=-115860000;
#10;x=-115850000;
#10;x=-115840000;
#10;x=-115830000;
#10;x=-115820000;
#10;x=-115810000;
#10;x=-115800000;
#10;x=-115790000;
#10;x=-115780000;
#10;x=-115770000;
#10;x=-115760000;
#10;x=-115750000;
#10;x=-115740000;
#10;x=-115730000;
#10;x=-115720000;
#10;x=-115710000;
#10;x=-115700000;
#10;x=-115690000;
#10;x=-115680000;
#10;x=-115670000;
#10;x=-115660000;
#10;x=-115650000;
#10;x=-115640000;
#10;x=-115630000;
#10;x=-115620000;
#10;x=-115610000;
#10;x=-115600000;
#10;x=-115590000;
#10;x=-115580000;
#10;x=-115570000;
#10;x=-115560000;
#10;x=-115550000;
#10;x=-115540000;
#10;x=-115530000;
#10;x=-115520000;
#10;x=-115510000;
#10;x=-115500000;
#10;x=-115490000;
#10;x=-115480000;
#10;x=-115470000;
#10;x=-115460000;
#10;x=-115450000;
#10;x=-115440000;
#10;x=-115430000;
#10;x=-115420000;
#10;x=-115410000;
#10;x=-115400000;
#10;x=-115390000;
#10;x=-115380000;
#10;x=-115370000;
#10;x=-115360000;
#10;x=-115350000;
#10;x=-115340000;
#10;x=-115330000;
#10;x=-115320000;
#10;x=-115310000;
#10;x=-115300000;
#10;x=-115290000;
#10;x=-115280000;
#10;x=-115270000;
#10;x=-115260000;
#10;x=-115250000;
#10;x=-115240000;
#10;x=-115230000;
#10;x=-115220000;
#10;x=-115210000;
#10;x=-115200000;
#10;x=-115190000;
#10;x=-115180000;
#10;x=-115170000;
#10;x=-115160000;
#10;x=-115150000;
#10;x=-115140000;
#10;x=-115130000;
#10;x=-115120000;
#10;x=-115110000;
#10;x=-115100000;
#10;x=-115090000;
#10;x=-115080000;
#10;x=-115070000;
#10;x=-115060000;
#10;x=-115050000;
#10;x=-115040000;
#10;x=-115030000;
#10;x=-115020000;
#10;x=-115010000;
#10;x=-115000000;
#10;x=-114990000;
#10;x=-114980000;
#10;x=-114970000;
#10;x=-114960000;
#10;x=-114950000;
#10;x=-114940000;
#10;x=-114930000;
#10;x=-114920000;
#10;x=-114910000;
#10;x=-114900000;
#10;x=-114890000;
#10;x=-114880000;
#10;x=-114870000;
#10;x=-114860000;
#10;x=-114850000;
#10;x=-114840000;
#10;x=-114830000;
#10;x=-114820000;
#10;x=-114810000;
#10;x=-114800000;
#10;x=-114790000;
#10;x=-114780000;
#10;x=-114770000;
#10;x=-114760000;
#10;x=-114750000;
#10;x=-114740000;
#10;x=-114730000;
#10;x=-114720000;
#10;x=-114710000;
#10;x=-114700000;
#10;x=-114690000;
#10;x=-114680000;
#10;x=-114670000;
#10;x=-114660000;
#10;x=-114650000;
#10;x=-114640000;
#10;x=-114630000;
#10;x=-114620000;
#10;x=-114610000;
#10;x=-114600000;
#10;x=-114590000;
#10;x=-114580000;
#10;x=-114570000;
#10;x=-114560000;
#10;x=-114550000;
#10;x=-114540000;
#10;x=-114530000;
#10;x=-114520000;
#10;x=-114510000;
#10;x=-114500000;
#10;x=-114490000;
#10;x=-114480000;
#10;x=-114470000;
#10;x=-114460000;
#10;x=-114450000;
#10;x=-114440000;
#10;x=-114430000;
#10;x=-114420000;
#10;x=-114410000;
#10;x=-114400000;
#10;x=-114390000;
#10;x=-114380000;
#10;x=-114370000;
#10;x=-114360000;
#10;x=-114350000;
#10;x=-114340000;
#10;x=-114330000;
#10;x=-114320000;
#10;x=-114310000;
#10;x=-114300000;
#10;x=-114290000;
#10;x=-114280000;
#10;x=-114270000;
#10;x=-114260000;
#10;x=-114250000;
#10;x=-114240000;
#10;x=-114230000;
#10;x=-114220000;
#10;x=-114210000;
#10;x=-114200000;
#10;x=-114190000;
#10;x=-114180000;
#10;x=-114170000;
#10;x=-114160000;
#10;x=-114150000;
#10;x=-114140000;
#10;x=-114130000;
#10;x=-114120000;
#10;x=-114110000;
#10;x=-114100000;
#10;x=-114090000;
#10;x=-114080000;
#10;x=-114070000;
#10;x=-114060000;
#10;x=-114050000;
#10;x=-114040000;
#10;x=-114030000;
#10;x=-114020000;
#10;x=-114010000;
#10;x=-114000000;
#10;x=-113990000;
#10;x=-113980000;
#10;x=-113970000;
#10;x=-113960000;
#10;x=-113950000;
#10;x=-113940000;
#10;x=-113930000;
#10;x=-113920000;
#10;x=-113910000;
#10;x=-113900000;
#10;x=-113890000;
#10;x=-113880000;
#10;x=-113870000;
#10;x=-113860000;
#10;x=-113850000;
#10;x=-113840000;
#10;x=-113830000;
#10;x=-113820000;
#10;x=-113810000;
#10;x=-113800000;
#10;x=-113790000;
#10;x=-113780000;
#10;x=-113770000;
#10;x=-113760000;
#10;x=-113750000;
#10;x=-113740000;
#10;x=-113730000;
#10;x=-113720000;
#10;x=-113710000;
#10;x=-113700000;
#10;x=-113690000;
#10;x=-113680000;
#10;x=-113670000;
#10;x=-113660000;
#10;x=-113650000;
#10;x=-113640000;
#10;x=-113630000;
#10;x=-113620000;
#10;x=-113610000;
#10;x=-113600000;
#10;x=-113590000;
#10;x=-113580000;
#10;x=-113570000;
#10;x=-113560000;
#10;x=-113550000;
#10;x=-113540000;
#10;x=-113530000;
#10;x=-113520000;
#10;x=-113510000;
#10;x=-113500000;
#10;x=-113490000;
#10;x=-113480000;
#10;x=-113470000;
#10;x=-113460000;
#10;x=-113450000;
#10;x=-113440000;
#10;x=-113430000;
#10;x=-113420000;
#10;x=-113410000;
#10;x=-113400000;
#10;x=-113390000;
#10;x=-113380000;
#10;x=-113370000;
#10;x=-113360000;
#10;x=-113350000;
#10;x=-113340000;
#10;x=-113330000;
#10;x=-113320000;
#10;x=-113310000;
#10;x=-113300000;
#10;x=-113290000;
#10;x=-113280000;
#10;x=-113270000;
#10;x=-113260000;
#10;x=-113250000;
#10;x=-113240000;
#10;x=-113230000;
#10;x=-113220000;
#10;x=-113210000;
#10;x=-113200000;
#10;x=-113190000;
#10;x=-113180000;
#10;x=-113170000;
#10;x=-113160000;
#10;x=-113150000;
#10;x=-113140000;
#10;x=-113130000;
#10;x=-113120000;
#10;x=-113110000;
#10;x=-113100000;
#10;x=-113090000;
#10;x=-113080000;
#10;x=-113070000;
#10;x=-113060000;
#10;x=-113050000;
#10;x=-113040000;
#10;x=-113030000;
#10;x=-113020000;
#10;x=-113010000;
#10;x=-113000000;
#10;x=-112990000;
#10;x=-112980000;
#10;x=-112970000;
#10;x=-112960000;
#10;x=-112950000;
#10;x=-112940000;
#10;x=-112930000;
#10;x=-112920000;
#10;x=-112910000;
#10;x=-112900000;
#10;x=-112890000;
#10;x=-112880000;
#10;x=-112870000;
#10;x=-112860000;
#10;x=-112850000;
#10;x=-112840000;
#10;x=-112830000;
#10;x=-112820000;
#10;x=-112810000;
#10;x=-112800000;
#10;x=-112790000;
#10;x=-112780000;
#10;x=-112770000;
#10;x=-112760000;
#10;x=-112750000;
#10;x=-112740000;
#10;x=-112730000;
#10;x=-112720000;
#10;x=-112710000;
#10;x=-112700000;
#10;x=-112690000;
#10;x=-112680000;
#10;x=-112670000;
#10;x=-112660000;
#10;x=-112650000;
#10;x=-112640000;
#10;x=-112630000;
#10;x=-112620000;
#10;x=-112610000;
#10;x=-112600000;
#10;x=-112590000;
#10;x=-112580000;
#10;x=-112570000;
#10;x=-112560000;
#10;x=-112550000;
#10;x=-112540000;
#10;x=-112530000;
#10;x=-112520000;
#10;x=-112510000;
#10;x=-112500000;
#10;x=-112490000;
#10;x=-112480000;
#10;x=-112470000;
#10;x=-112460000;
#10;x=-112450000;
#10;x=-112440000;
#10;x=-112430000;
#10;x=-112420000;
#10;x=-112410000;
#10;x=-112400000;
#10;x=-112390000;
#10;x=-112380000;
#10;x=-112370000;
#10;x=-112360000;
#10;x=-112350000;
#10;x=-112340000;
#10;x=-112330000;
#10;x=-112320000;
#10;x=-112310000;
#10;x=-112300000;
#10;x=-112290000;
#10;x=-112280000;
#10;x=-112270000;
#10;x=-112260000;
#10;x=-112250000;
#10;x=-112240000;
#10;x=-112230000;
#10;x=-112220000;
#10;x=-112210000;
#10;x=-112200000;
#10;x=-112190000;
#10;x=-112180000;
#10;x=-112170000;
#10;x=-112160000;
#10;x=-112150000;
#10;x=-112140000;
#10;x=-112130000;
#10;x=-112120000;
#10;x=-112110000;
#10;x=-112100000;
#10;x=-112090000;
#10;x=-112080000;
#10;x=-112070000;
#10;x=-112060000;
#10;x=-112050000;
#10;x=-112040000;
#10;x=-112030000;
#10;x=-112020000;
#10;x=-112010000;
#10;x=-112000000;
#10;x=-111990000;
#10;x=-111980000;
#10;x=-111970000;
#10;x=-111960000;
#10;x=-111950000;
#10;x=-111940000;
#10;x=-111930000;
#10;x=-111920000;
#10;x=-111910000;
#10;x=-111900000;
#10;x=-111890000;
#10;x=-111880000;
#10;x=-111870000;
#10;x=-111860000;
#10;x=-111850000;
#10;x=-111840000;
#10;x=-111830000;
#10;x=-111820000;
#10;x=-111810000;
#10;x=-111800000;
#10;x=-111790000;
#10;x=-111780000;
#10;x=-111770000;
#10;x=-111760000;
#10;x=-111750000;
#10;x=-111740000;
#10;x=-111730000;
#10;x=-111720000;
#10;x=-111710000;
#10;x=-111700000;
#10;x=-111690000;
#10;x=-111680000;
#10;x=-111670000;
#10;x=-111660000;
#10;x=-111650000;
#10;x=-111640000;
#10;x=-111630000;
#10;x=-111620000;
#10;x=-111610000;
#10;x=-111600000;
#10;x=-111590000;
#10;x=-111580000;
#10;x=-111570000;
#10;x=-111560000;
#10;x=-111550000;
#10;x=-111540000;
#10;x=-111530000;
#10;x=-111520000;
#10;x=-111510000;
#10;x=-111500000;
#10;x=-111490000;
#10;x=-111480000;
#10;x=-111470000;
#10;x=-111460000;
#10;x=-111450000;
#10;x=-111440000;
#10;x=-111430000;
#10;x=-111420000;
#10;x=-111410000;
#10;x=-111400000;
#10;x=-111390000;
#10;x=-111380000;
#10;x=-111370000;
#10;x=-111360000;
#10;x=-111350000;
#10;x=-111340000;
#10;x=-111330000;
#10;x=-111320000;
#10;x=-111310000;
#10;x=-111300000;
#10;x=-111290000;
#10;x=-111280000;
#10;x=-111270000;
#10;x=-111260000;
#10;x=-111250000;
#10;x=-111240000;
#10;x=-111230000;
#10;x=-111220000;
#10;x=-111210000;
#10;x=-111200000;
#10;x=-111190000;
#10;x=-111180000;
#10;x=-111170000;
#10;x=-111160000;
#10;x=-111150000;
#10;x=-111140000;
#10;x=-111130000;
#10;x=-111120000;
#10;x=-111110000;
#10;x=-111100000;
#10;x=-111090000;
#10;x=-111080000;
#10;x=-111070000;
#10;x=-111060000;
#10;x=-111050000;
#10;x=-111040000;
#10;x=-111030000;
#10;x=-111020000;
#10;x=-111010000;
#10;x=-111000000;
#10;x=-110990000;
#10;x=-110980000;
#10;x=-110970000;
#10;x=-110960000;
#10;x=-110950000;
#10;x=-110940000;
#10;x=-110930000;
#10;x=-110920000;
#10;x=-110910000;
#10;x=-110900000;
#10;x=-110890000;
#10;x=-110880000;
#10;x=-110870000;
#10;x=-110860000;
#10;x=-110850000;
#10;x=-110840000;
#10;x=-110830000;
#10;x=-110820000;
#10;x=-110810000;
#10;x=-110800000;
#10;x=-110790000;
#10;x=-110780000;
#10;x=-110770000;
#10;x=-110760000;
#10;x=-110750000;
#10;x=-110740000;
#10;x=-110730000;
#10;x=-110720000;
#10;x=-110710000;
#10;x=-110700000;
#10;x=-110690000;
#10;x=-110680000;
#10;x=-110670000;
#10;x=-110660000;
#10;x=-110650000;
#10;x=-110640000;
#10;x=-110630000;
#10;x=-110620000;
#10;x=-110610000;
#10;x=-110600000;
#10;x=-110590000;
#10;x=-110580000;
#10;x=-110570000;
#10;x=-110560000;
#10;x=-110550000;
#10;x=-110540000;
#10;x=-110530000;
#10;x=-110520000;
#10;x=-110510000;
#10;x=-110500000;
#10;x=-110490000;
#10;x=-110480000;
#10;x=-110470000;
#10;x=-110460000;
#10;x=-110450000;
#10;x=-110440000;
#10;x=-110430000;
#10;x=-110420000;
#10;x=-110410000;
#10;x=-110400000;
#10;x=-110390000;
#10;x=-110380000;
#10;x=-110370000;
#10;x=-110360000;
#10;x=-110350000;
#10;x=-110340000;
#10;x=-110330000;
#10;x=-110320000;
#10;x=-110310000;
#10;x=-110300000;
#10;x=-110290000;
#10;x=-110280000;
#10;x=-110270000;
#10;x=-110260000;
#10;x=-110250000;
#10;x=-110240000;
#10;x=-110230000;
#10;x=-110220000;
#10;x=-110210000;
#10;x=-110200000;
#10;x=-110190000;
#10;x=-110180000;
#10;x=-110170000;
#10;x=-110160000;
#10;x=-110150000;
#10;x=-110140000;
#10;x=-110130000;
#10;x=-110120000;
#10;x=-110110000;
#10;x=-110100000;
#10;x=-110090000;
#10;x=-110080000;
#10;x=-110070000;
#10;x=-110060000;
#10;x=-110050000;
#10;x=-110040000;
#10;x=-110030000;
#10;x=-110020000;
#10;x=-110010000;
#10;x=-110000000;
#10;x=-109990000;
#10;x=-109980000;
#10;x=-109970000;
#10;x=-109960000;
#10;x=-109950000;
#10;x=-109940000;
#10;x=-109930000;
#10;x=-109920000;
#10;x=-109910000;
#10;x=-109900000;
#10;x=-109890000;
#10;x=-109880000;
#10;x=-109870000;
#10;x=-109860000;
#10;x=-109850000;
#10;x=-109840000;
#10;x=-109830000;
#10;x=-109820000;
#10;x=-109810000;
#10;x=-109800000;
#10;x=-109790000;
#10;x=-109780000;
#10;x=-109770000;
#10;x=-109760000;
#10;x=-109750000;
#10;x=-109740000;
#10;x=-109730000;
#10;x=-109720000;
#10;x=-109710000;
#10;x=-109700000;
#10;x=-109690000;
#10;x=-109680000;
#10;x=-109670000;
#10;x=-109660000;
#10;x=-109650000;
#10;x=-109640000;
#10;x=-109630000;
#10;x=-109620000;
#10;x=-109610000;
#10;x=-109600000;
#10;x=-109590000;
#10;x=-109580000;
#10;x=-109570000;
#10;x=-109560000;
#10;x=-109550000;
#10;x=-109540000;
#10;x=-109530000;
#10;x=-109520000;
#10;x=-109510000;
#10;x=-109500000;
#10;x=-109490000;
#10;x=-109480000;
#10;x=-109470000;
#10;x=-109460000;
#10;x=-109450000;
#10;x=-109440000;
#10;x=-109430000;
#10;x=-109420000;
#10;x=-109410000;
#10;x=-109400000;
#10;x=-109390000;
#10;x=-109380000;
#10;x=-109370000;
#10;x=-109360000;
#10;x=-109350000;
#10;x=-109340000;
#10;x=-109330000;
#10;x=-109320000;
#10;x=-109310000;
#10;x=-109300000;
#10;x=-109290000;
#10;x=-109280000;
#10;x=-109270000;
#10;x=-109260000;
#10;x=-109250000;
#10;x=-109240000;
#10;x=-109230000;
#10;x=-109220000;
#10;x=-109210000;
#10;x=-109200000;
#10;x=-109190000;
#10;x=-109180000;
#10;x=-109170000;
#10;x=-109160000;
#10;x=-109150000;
#10;x=-109140000;
#10;x=-109130000;
#10;x=-109120000;
#10;x=-109110000;
#10;x=-109100000;
#10;x=-109090000;
#10;x=-109080000;
#10;x=-109070000;
#10;x=-109060000;
#10;x=-109050000;
#10;x=-109040000;
#10;x=-109030000;
#10;x=-109020000;
#10;x=-109010000;
#10;x=-109000000;
#10;x=-108990000;
#10;x=-108980000;
#10;x=-108970000;
#10;x=-108960000;
#10;x=-108950000;
#10;x=-108940000;
#10;x=-108930000;
#10;x=-108920000;
#10;x=-108910000;
#10;x=-108900000;
#10;x=-108890000;
#10;x=-108880000;
#10;x=-108870000;
#10;x=-108860000;
#10;x=-108850000;
#10;x=-108840000;
#10;x=-108830000;
#10;x=-108820000;
#10;x=-108810000;
#10;x=-108800000;
#10;x=-108790000;
#10;x=-108780000;
#10;x=-108770000;
#10;x=-108760000;
#10;x=-108750000;
#10;x=-108740000;
#10;x=-108730000;
#10;x=-108720000;
#10;x=-108710000;
#10;x=-108700000;
#10;x=-108690000;
#10;x=-108680000;
#10;x=-108670000;
#10;x=-108660000;
#10;x=-108650000;
#10;x=-108640000;
#10;x=-108630000;
#10;x=-108620000;
#10;x=-108610000;
#10;x=-108600000;
#10;x=-108590000;
#10;x=-108580000;
#10;x=-108570000;
#10;x=-108560000;
#10;x=-108550000;
#10;x=-108540000;
#10;x=-108530000;
#10;x=-108520000;
#10;x=-108510000;
#10;x=-108500000;
#10;x=-108490000;
#10;x=-108480000;
#10;x=-108470000;
#10;x=-108460000;
#10;x=-108450000;
#10;x=-108440000;
#10;x=-108430000;
#10;x=-108420000;
#10;x=-108410000;
#10;x=-108400000;
#10;x=-108390000;
#10;x=-108380000;
#10;x=-108370000;
#10;x=-108360000;
#10;x=-108350000;
#10;x=-108340000;
#10;x=-108330000;
#10;x=-108320000;
#10;x=-108310000;
#10;x=-108300000;
#10;x=-108290000;
#10;x=-108280000;
#10;x=-108270000;
#10;x=-108260000;
#10;x=-108250000;
#10;x=-108240000;
#10;x=-108230000;
#10;x=-108220000;
#10;x=-108210000;
#10;x=-108200000;
#10;x=-108190000;
#10;x=-108180000;
#10;x=-108170000;
#10;x=-108160000;
#10;x=-108150000;
#10;x=-108140000;
#10;x=-108130000;
#10;x=-108120000;
#10;x=-108110000;
#10;x=-108100000;
#10;x=-108090000;
#10;x=-108080000;
#10;x=-108070000;
#10;x=-108060000;
#10;x=-108050000;
#10;x=-108040000;
#10;x=-108030000;
#10;x=-108020000;
#10;x=-108010000;
#10;x=-108000000;
#10;x=-107990000;
#10;x=-107980000;
#10;x=-107970000;
#10;x=-107960000;
#10;x=-107950000;
#10;x=-107940000;
#10;x=-107930000;
#10;x=-107920000;
#10;x=-107910000;
#10;x=-107900000;
#10;x=-107890000;
#10;x=-107880000;
#10;x=-107870000;
#10;x=-107860000;
#10;x=-107850000;
#10;x=-107840000;
#10;x=-107830000;
#10;x=-107820000;
#10;x=-107810000;
#10;x=-107800000;
#10;x=-107790000;
#10;x=-107780000;
#10;x=-107770000;
#10;x=-107760000;
#10;x=-107750000;
#10;x=-107740000;
#10;x=-107730000;
#10;x=-107720000;
#10;x=-107710000;
#10;x=-107700000;
#10;x=-107690000;
#10;x=-107680000;
#10;x=-107670000;
#10;x=-107660000;
#10;x=-107650000;
#10;x=-107640000;
#10;x=-107630000;
#10;x=-107620000;
#10;x=-107610000;
#10;x=-107600000;
#10;x=-107590000;
#10;x=-107580000;
#10;x=-107570000;
#10;x=-107560000;
#10;x=-107550000;
#10;x=-107540000;
#10;x=-107530000;
#10;x=-107520000;
#10;x=-107510000;
#10;x=-107500000;
#10;x=-107490000;
#10;x=-107480000;
#10;x=-107470000;
#10;x=-107460000;
#10;x=-107450000;
#10;x=-107440000;
#10;x=-107430000;
#10;x=-107420000;
#10;x=-107410000;
#10;x=-107400000;
#10;x=-107390000;
#10;x=-107380000;
#10;x=-107370000;
#10;x=-107360000;
#10;x=-107350000;
#10;x=-107340000;
#10;x=-107330000;
#10;x=-107320000;
#10;x=-107310000;
#10;x=-107300000;
#10;x=-107290000;
#10;x=-107280000;
#10;x=-107270000;
#10;x=-107260000;
#10;x=-107250000;
#10;x=-107240000;
#10;x=-107230000;
#10;x=-107220000;
#10;x=-107210000;
#10;x=-107200000;
#10;x=-107190000;
#10;x=-107180000;
#10;x=-107170000;
#10;x=-107160000;
#10;x=-107150000;
#10;x=-107140000;
#10;x=-107130000;
#10;x=-107120000;
#10;x=-107110000;
#10;x=-107100000;
#10;x=-107090000;
#10;x=-107080000;
#10;x=-107070000;
#10;x=-107060000;
#10;x=-107050000;
#10;x=-107040000;
#10;x=-107030000;
#10;x=-107020000;
#10;x=-107010000;
#10;x=-107000000;
#10;x=-106990000;
#10;x=-106980000;
#10;x=-106970000;
#10;x=-106960000;
#10;x=-106950000;
#10;x=-106940000;
#10;x=-106930000;
#10;x=-106920000;
#10;x=-106910000;
#10;x=-106900000;
#10;x=-106890000;
#10;x=-106880000;
#10;x=-106870000;
#10;x=-106860000;
#10;x=-106850000;
#10;x=-106840000;
#10;x=-106830000;
#10;x=-106820000;
#10;x=-106810000;
#10;x=-106800000;
#10;x=-106790000;
#10;x=-106780000;
#10;x=-106770000;
#10;x=-106760000;
#10;x=-106750000;
#10;x=-106740000;
#10;x=-106730000;
#10;x=-106720000;
#10;x=-106710000;
#10;x=-106700000;
#10;x=-106690000;
#10;x=-106680000;
#10;x=-106670000;
#10;x=-106660000;
#10;x=-106650000;
#10;x=-106640000;
#10;x=-106630000;
#10;x=-106620000;
#10;x=-106610000;
#10;x=-106600000;
#10;x=-106590000;
#10;x=-106580000;
#10;x=-106570000;
#10;x=-106560000;
#10;x=-106550000;
#10;x=-106540000;
#10;x=-106530000;
#10;x=-106520000;
#10;x=-106510000;
#10;x=-106500000;
#10;x=-106490000;
#10;x=-106480000;
#10;x=-106470000;
#10;x=-106460000;
#10;x=-106450000;
#10;x=-106440000;
#10;x=-106430000;
#10;x=-106420000;
#10;x=-106410000;
#10;x=-106400000;
#10;x=-106390000;
#10;x=-106380000;
#10;x=-106370000;
#10;x=-106360000;
#10;x=-106350000;
#10;x=-106340000;
#10;x=-106330000;
#10;x=-106320000;
#10;x=-106310000;
#10;x=-106300000;
#10;x=-106290000;
#10;x=-106280000;
#10;x=-106270000;
#10;x=-106260000;
#10;x=-106250000;
#10;x=-106240000;
#10;x=-106230000;
#10;x=-106220000;
#10;x=-106210000;
#10;x=-106200000;
#10;x=-106190000;
#10;x=-106180000;
#10;x=-106170000;
#10;x=-106160000;
#10;x=-106150000;
#10;x=-106140000;
#10;x=-106130000;
#10;x=-106120000;
#10;x=-106110000;
#10;x=-106100000;
#10;x=-106090000;
#10;x=-106080000;
#10;x=-106070000;
#10;x=-106060000;
#10;x=-106050000;
#10;x=-106040000;
#10;x=-106030000;
#10;x=-106020000;
#10;x=-106010000;
#10;x=-106000000;
#10;x=-105990000;
#10;x=-105980000;
#10;x=-105970000;
#10;x=-105960000;
#10;x=-105950000;
#10;x=-105940000;
#10;x=-105930000;
#10;x=-105920000;
#10;x=-105910000;
#10;x=-105900000;
#10;x=-105890000;
#10;x=-105880000;
#10;x=-105870000;
#10;x=-105860000;
#10;x=-105850000;
#10;x=-105840000;
#10;x=-105830000;
#10;x=-105820000;
#10;x=-105810000;
#10;x=-105800000;
#10;x=-105790000;
#10;x=-105780000;
#10;x=-105770000;
#10;x=-105760000;
#10;x=-105750000;
#10;x=-105740000;
#10;x=-105730000;
#10;x=-105720000;
#10;x=-105710000;
#10;x=-105700000;
#10;x=-105690000;
#10;x=-105680000;
#10;x=-105670000;
#10;x=-105660000;
#10;x=-105650000;
#10;x=-105640000;
#10;x=-105630000;
#10;x=-105620000;
#10;x=-105610000;
#10;x=-105600000;
#10;x=-105590000;
#10;x=-105580000;
#10;x=-105570000;
#10;x=-105560000;
#10;x=-105550000;
#10;x=-105540000;
#10;x=-105530000;
#10;x=-105520000;
#10;x=-105510000;
#10;x=-105500000;
#10;x=-105490000;
#10;x=-105480000;
#10;x=-105470000;
#10;x=-105460000;
#10;x=-105450000;
#10;x=-105440000;
#10;x=-105430000;
#10;x=-105420000;
#10;x=-105410000;
#10;x=-105400000;
#10;x=-105390000;
#10;x=-105380000;
#10;x=-105370000;
#10;x=-105360000;
#10;x=-105350000;
#10;x=-105340000;
#10;x=-105330000;
#10;x=-105320000;
#10;x=-105310000;
#10;x=-105300000;
#10;x=-105290000;
#10;x=-105280000;
#10;x=-105270000;
#10;x=-105260000;
#10;x=-105250000;
#10;x=-105240000;
#10;x=-105230000;
#10;x=-105220000;
#10;x=-105210000;
#10;x=-105200000;
#10;x=-105190000;
#10;x=-105180000;
#10;x=-105170000;
#10;x=-105160000;
#10;x=-105150000;
#10;x=-105140000;
#10;x=-105130000;
#10;x=-105120000;
#10;x=-105110000;
#10;x=-105100000;
#10;x=-105090000;
#10;x=-105080000;
#10;x=-105070000;
#10;x=-105060000;
#10;x=-105050000;
#10;x=-105040000;
#10;x=-105030000;
#10;x=-105020000;
#10;x=-105010000;
#10;x=-105000000;
#10;x=-104990000;
#10;x=-104980000;
#10;x=-104970000;
#10;x=-104960000;
#10;x=-104950000;
#10;x=-104940000;
#10;x=-104930000;
#10;x=-104920000;
#10;x=-104910000;
#10;x=-104900000;
#10;x=-104890000;
#10;x=-104880000;
#10;x=-104870000;
#10;x=-104860000;
#10;x=-104850000;
#10;x=-104840000;
#10;x=-104830000;
#10;x=-104820000;
#10;x=-104810000;
#10;x=-104800000;
#10;x=-104790000;
#10;x=-104780000;
#10;x=-104770000;
#10;x=-104760000;
#10;x=-104750000;
#10;x=-104740000;
#10;x=-104730000;
#10;x=-104720000;
#10;x=-104710000;
#10;x=-104700000;
#10;x=-104690000;
#10;x=-104680000;
#10;x=-104670000;
#10;x=-104660000;
#10;x=-104650000;
#10;x=-104640000;
#10;x=-104630000;
#10;x=-104620000;
#10;x=-104610000;
#10;x=-104600000;
#10;x=-104590000;
#10;x=-104580000;
#10;x=-104570000;
#10;x=-104560000;
#10;x=-104550000;
#10;x=-104540000;
#10;x=-104530000;
#10;x=-104520000;
#10;x=-104510000;
#10;x=-104500000;
#10;x=-104490000;
#10;x=-104480000;
#10;x=-104470000;
#10;x=-104460000;
#10;x=-104450000;
#10;x=-104440000;
#10;x=-104430000;
#10;x=-104420000;
#10;x=-104410000;
#10;x=-104400000;
#10;x=-104390000;
#10;x=-104380000;
#10;x=-104370000;
#10;x=-104360000;
#10;x=-104350000;
#10;x=-104340000;
#10;x=-104330000;
#10;x=-104320000;
#10;x=-104310000;
#10;x=-104300000;
#10;x=-104290000;
#10;x=-104280000;
#10;x=-104270000;
#10;x=-104260000;
#10;x=-104250000;
#10;x=-104240000;
#10;x=-104230000;
#10;x=-104220000;
#10;x=-104210000;
#10;x=-104200000;
#10;x=-104190000;
#10;x=-104180000;
#10;x=-104170000;
#10;x=-104160000;
#10;x=-104150000;
#10;x=-104140000;
#10;x=-104130000;
#10;x=-104120000;
#10;x=-104110000;
#10;x=-104100000;
#10;x=-104090000;
#10;x=-104080000;
#10;x=-104070000;
#10;x=-104060000;
#10;x=-104050000;
#10;x=-104040000;
#10;x=-104030000;
#10;x=-104020000;
#10;x=-104010000;
#10;x=-104000000;
#10;x=-103990000;
#10;x=-103980000;
#10;x=-103970000;
#10;x=-103960000;
#10;x=-103950000;
#10;x=-103940000;
#10;x=-103930000;
#10;x=-103920000;
#10;x=-103910000;
#10;x=-103900000;
#10;x=-103890000;
#10;x=-103880000;
#10;x=-103870000;
#10;x=-103860000;
#10;x=-103850000;
#10;x=-103840000;
#10;x=-103830000;
#10;x=-103820000;
#10;x=-103810000;
#10;x=-103800000;
#10;x=-103790000;
#10;x=-103780000;
#10;x=-103770000;
#10;x=-103760000;
#10;x=-103750000;
#10;x=-103740000;
#10;x=-103730000;
#10;x=-103720000;
#10;x=-103710000;
#10;x=-103700000;
#10;x=-103690000;
#10;x=-103680000;
#10;x=-103670000;
#10;x=-103660000;
#10;x=-103650000;
#10;x=-103640000;
#10;x=-103630000;
#10;x=-103620000;
#10;x=-103610000;
#10;x=-103600000;
#10;x=-103590000;
#10;x=-103580000;
#10;x=-103570000;
#10;x=-103560000;
#10;x=-103550000;
#10;x=-103540000;
#10;x=-103530000;
#10;x=-103520000;
#10;x=-103510000;
#10;x=-103500000;
#10;x=-103490000;
#10;x=-103480000;
#10;x=-103470000;
#10;x=-103460000;
#10;x=-103450000;
#10;x=-103440000;
#10;x=-103430000;
#10;x=-103420000;
#10;x=-103410000;
#10;x=-103400000;
#10;x=-103390000;
#10;x=-103380000;
#10;x=-103370000;
#10;x=-103360000;
#10;x=-103350000;
#10;x=-103340000;
#10;x=-103330000;
#10;x=-103320000;
#10;x=-103310000;
#10;x=-103300000;
#10;x=-103290000;
#10;x=-103280000;
#10;x=-103270000;
#10;x=-103260000;
#10;x=-103250000;
#10;x=-103240000;
#10;x=-103230000;
#10;x=-103220000;
#10;x=-103210000;
#10;x=-103200000;
#10;x=-103190000;
#10;x=-103180000;
#10;x=-103170000;
#10;x=-103160000;
#10;x=-103150000;
#10;x=-103140000;
#10;x=-103130000;
#10;x=-103120000;
#10;x=-103110000;
#10;x=-103100000;
#10;x=-103090000;
#10;x=-103080000;
#10;x=-103070000;
#10;x=-103060000;
#10;x=-103050000;
#10;x=-103040000;
#10;x=-103030000;
#10;x=-103020000;
#10;x=-103010000;
#10;x=-103000000;
#10;x=-102990000;
#10;x=-102980000;
#10;x=-102970000;
#10;x=-102960000;
#10;x=-102950000;
#10;x=-102940000;
#10;x=-102930000;
#10;x=-102920000;
#10;x=-102910000;
#10;x=-102900000;
#10;x=-102890000;
#10;x=-102880000;
#10;x=-102870000;
#10;x=-102860000;
#10;x=-102850000;
#10;x=-102840000;
#10;x=-102830000;
#10;x=-102820000;
#10;x=-102810000;
#10;x=-102800000;
#10;x=-102790000;
#10;x=-102780000;
#10;x=-102770000;
#10;x=-102760000;
#10;x=-102750000;
#10;x=-102740000;
#10;x=-102730000;
#10;x=-102720000;
#10;x=-102710000;
#10;x=-102700000;
#10;x=-102690000;
#10;x=-102680000;
#10;x=-102670000;
#10;x=-102660000;
#10;x=-102650000;
#10;x=-102640000;
#10;x=-102630000;
#10;x=-102620000;
#10;x=-102610000;
#10;x=-102600000;
#10;x=-102590000;
#10;x=-102580000;
#10;x=-102570000;
#10;x=-102560000;
#10;x=-102550000;
#10;x=-102540000;
#10;x=-102530000;
#10;x=-102520000;
#10;x=-102510000;
#10;x=-102500000;
#10;x=-102490000;
#10;x=-102480000;
#10;x=-102470000;
#10;x=-102460000;
#10;x=-102450000;
#10;x=-102440000;
#10;x=-102430000;
#10;x=-102420000;
#10;x=-102410000;
#10;x=-102400000;
#10;x=-102390000;
#10;x=-102380000;
#10;x=-102370000;
#10;x=-102360000;
#10;x=-102350000;
#10;x=-102340000;
#10;x=-102330000;
#10;x=-102320000;
#10;x=-102310000;
#10;x=-102300000;
#10;x=-102290000;
#10;x=-102280000;
#10;x=-102270000;
#10;x=-102260000;
#10;x=-102250000;
#10;x=-102240000;
#10;x=-102230000;
#10;x=-102220000;
#10;x=-102210000;
#10;x=-102200000;
#10;x=-102190000;
#10;x=-102180000;
#10;x=-102170000;
#10;x=-102160000;
#10;x=-102150000;
#10;x=-102140000;
#10;x=-102130000;
#10;x=-102120000;
#10;x=-102110000;
#10;x=-102100000;
#10;x=-102090000;
#10;x=-102080000;
#10;x=-102070000;
#10;x=-102060000;
#10;x=-102050000;
#10;x=-102040000;
#10;x=-102030000;
#10;x=-102020000;
#10;x=-102010000;
#10;x=-102000000;
#10;x=-101990000;
#10;x=-101980000;
#10;x=-101970000;
#10;x=-101960000;
#10;x=-101950000;
#10;x=-101940000;
#10;x=-101930000;
#10;x=-101920000;
#10;x=-101910000;
#10;x=-101900000;
#10;x=-101890000;
#10;x=-101880000;
#10;x=-101870000;
#10;x=-101860000;
#10;x=-101850000;
#10;x=-101840000;
#10;x=-101830000;
#10;x=-101820000;
#10;x=-101810000;
#10;x=-101800000;
#10;x=-101790000;
#10;x=-101780000;
#10;x=-101770000;
#10;x=-101760000;
#10;x=-101750000;
#10;x=-101740000;
#10;x=-101730000;
#10;x=-101720000;
#10;x=-101710000;
#10;x=-101700000;
#10;x=-101690000;
#10;x=-101680000;
#10;x=-101670000;
#10;x=-101660000;
#10;x=-101650000;
#10;x=-101640000;
#10;x=-101630000;
#10;x=-101620000;
#10;x=-101610000;
#10;x=-101600000;
#10;x=-101590000;
#10;x=-101580000;
#10;x=-101570000;
#10;x=-101560000;
#10;x=-101550000;
#10;x=-101540000;
#10;x=-101530000;
#10;x=-101520000;
#10;x=-101510000;
#10;x=-101500000;
#10;x=-101490000;
#10;x=-101480000;
#10;x=-101470000;
#10;x=-101460000;
#10;x=-101450000;
#10;x=-101440000;
#10;x=-101430000;
#10;x=-101420000;
#10;x=-101410000;
#10;x=-101400000;
#10;x=-101390000;
#10;x=-101380000;
#10;x=-101370000;
#10;x=-101360000;
#10;x=-101350000;
#10;x=-101340000;
#10;x=-101330000;
#10;x=-101320000;
#10;x=-101310000;
#10;x=-101300000;
#10;x=-101290000;
#10;x=-101280000;
#10;x=-101270000;
#10;x=-101260000;
#10;x=-101250000;
#10;x=-101240000;
#10;x=-101230000;
#10;x=-101220000;
#10;x=-101210000;
#10;x=-101200000;
#10;x=-101190000;
#10;x=-101180000;
#10;x=-101170000;
#10;x=-101160000;
#10;x=-101150000;
#10;x=-101140000;
#10;x=-101130000;
#10;x=-101120000;
#10;x=-101110000;
#10;x=-101100000;
#10;x=-101090000;
#10;x=-101080000;
#10;x=-101070000;
#10;x=-101060000;
#10;x=-101050000;
#10;x=-101040000;
#10;x=-101030000;
#10;x=-101020000;
#10;x=-101010000;
#10;x=-101000000;
#10;x=-100990000;
#10;x=-100980000;
#10;x=-100970000;
#10;x=-100960000;
#10;x=-100950000;
#10;x=-100940000;
#10;x=-100930000;
#10;x=-100920000;
#10;x=-100910000;
#10;x=-100900000;
#10;x=-100890000;
#10;x=-100880000;
#10;x=-100870000;
#10;x=-100860000;
#10;x=-100850000;
#10;x=-100840000;
#10;x=-100830000;
#10;x=-100820000;
#10;x=-100810000;
#10;x=-100800000;
#10;x=-100790000;
#10;x=-100780000;
#10;x=-100770000;
#10;x=-100760000;
#10;x=-100750000;
#10;x=-100740000;
#10;x=-100730000;
#10;x=-100720000;
#10;x=-100710000;
#10;x=-100700000;
#10;x=-100690000;
#10;x=-100680000;
#10;x=-100670000;
#10;x=-100660000;
#10;x=-100650000;
#10;x=-100640000;
#10;x=-100630000;
#10;x=-100620000;
#10;x=-100610000;
#10;x=-100600000;
#10;x=-100590000;
#10;x=-100580000;
#10;x=-100570000;
#10;x=-100560000;
#10;x=-100550000;
#10;x=-100540000;
#10;x=-100530000;
#10;x=-100520000;
#10;x=-100510000;
#10;x=-100500000;
#10;x=-100490000;
#10;x=-100480000;
#10;x=-100470000;
#10;x=-100460000;
#10;x=-100450000;
#10;x=-100440000;
#10;x=-100430000;
#10;x=-100420000;
#10;x=-100410000;
#10;x=-100400000;
#10;x=-100390000;
#10;x=-100380000;
#10;x=-100370000;
#10;x=-100360000;
#10;x=-100350000;
#10;x=-100340000;
#10;x=-100330000;
#10;x=-100320000;
#10;x=-100310000;
#10;x=-100300000;
#10;x=-100290000;
#10;x=-100280000;
#10;x=-100270000;
#10;x=-100260000;
#10;x=-100250000;
#10;x=-100240000;
#10;x=-100230000;
#10;x=-100220000;
#10;x=-100210000;
#10;x=-100200000;
#10;x=-100190000;
#10;x=-100180000;
#10;x=-100170000;
#10;x=-100160000;
#10;x=-100150000;
#10;x=-100140000;
#10;x=-100130000;
#10;x=-100120000;
#10;x=-100110000;
#10;x=-100100000;
#10;x=-100090000;
#10;x=-100080000;
#10;x=-100070000;
#10;x=-100060000;
#10;x=-100050000;
#10;x=-100040000;
#10;x=-100030000;
#10;x=-100020000;
#10;x=-100010000;
#10;x=-100000000;
#10;x=-99990000;
#10;x=-99980000;
#10;x=-99970000;
#10;x=-99960000;
#10;x=-99950000;
#10;x=-99940000;
#10;x=-99930000;
#10;x=-99920000;
#10;x=-99910000;
#10;x=-99900000;
#10;x=-99890000;
#10;x=-99880000;
#10;x=-99870000;
#10;x=-99860000;
#10;x=-99850000;
#10;x=-99840000;
#10;x=-99830000;
#10;x=-99820000;
#10;x=-99810000;
#10;x=-99800000;
#10;x=-99790000;
#10;x=-99780000;
#10;x=-99770000;
#10;x=-99760000;
#10;x=-99750000;
#10;x=-99740000;
#10;x=-99730000;
#10;x=-99720000;
#10;x=-99710000;
#10;x=-99700000;
#10;x=-99690000;
#10;x=-99680000;
#10;x=-99670000;
#10;x=-99660000;
#10;x=-99650000;
#10;x=-99640000;
#10;x=-99630000;
#10;x=-99620000;
#10;x=-99610000;
#10;x=-99600000;
#10;x=-99590000;
#10;x=-99580000;
#10;x=-99570000;
#10;x=-99560000;
#10;x=-99550000;
#10;x=-99540000;
#10;x=-99530000;
#10;x=-99520000;
#10;x=-99510000;
#10;x=-99500000;
#10;x=-99490000;
#10;x=-99480000;
#10;x=-99470000;
#10;x=-99460000;
#10;x=-99450000;
#10;x=-99440000;
#10;x=-99430000;
#10;x=-99420000;
#10;x=-99410000;
#10;x=-99400000;
#10;x=-99390000;
#10;x=-99380000;
#10;x=-99370000;
#10;x=-99360000;
#10;x=-99350000;
#10;x=-99340000;
#10;x=-99330000;
#10;x=-99320000;
#10;x=-99310000;
#10;x=-99300000;
#10;x=-99290000;
#10;x=-99280000;
#10;x=-99270000;
#10;x=-99260000;
#10;x=-99250000;
#10;x=-99240000;
#10;x=-99230000;
#10;x=-99220000;
#10;x=-99210000;
#10;x=-99200000;
#10;x=-99190000;
#10;x=-99180000;
#10;x=-99170000;
#10;x=-99160000;
#10;x=-99150000;
#10;x=-99140000;
#10;x=-99130000;
#10;x=-99120000;
#10;x=-99110000;
#10;x=-99100000;
#10;x=-99090000;
#10;x=-99080000;
#10;x=-99070000;
#10;x=-99060000;
#10;x=-99050000;
#10;x=-99040000;
#10;x=-99030000;
#10;x=-99020000;
#10;x=-99010000;
#10;x=-99000000;
#10;x=-98990000;
#10;x=-98980000;
#10;x=-98970000;
#10;x=-98960000;
#10;x=-98950000;
#10;x=-98940000;
#10;x=-98930000;
#10;x=-98920000;
#10;x=-98910000;
#10;x=-98900000;
#10;x=-98890000;
#10;x=-98880000;
#10;x=-98870000;
#10;x=-98860000;
#10;x=-98850000;
#10;x=-98840000;
#10;x=-98830000;
#10;x=-98820000;
#10;x=-98810000;
#10;x=-98800000;
#10;x=-98790000;
#10;x=-98780000;
#10;x=-98770000;
#10;x=-98760000;
#10;x=-98750000;
#10;x=-98740000;
#10;x=-98730000;
#10;x=-98720000;
#10;x=-98710000;
#10;x=-98700000;
#10;x=-98690000;
#10;x=-98680000;
#10;x=-98670000;
#10;x=-98660000;
#10;x=-98650000;
#10;x=-98640000;
#10;x=-98630000;
#10;x=-98620000;
#10;x=-98610000;
#10;x=-98600000;
#10;x=-98590000;
#10;x=-98580000;
#10;x=-98570000;
#10;x=-98560000;
#10;x=-98550000;
#10;x=-98540000;
#10;x=-98530000;
#10;x=-98520000;
#10;x=-98510000;
#10;x=-98500000;
#10;x=-98490000;
#10;x=-98480000;
#10;x=-98470000;
#10;x=-98460000;
#10;x=-98450000;
#10;x=-98440000;
#10;x=-98430000;
#10;x=-98420000;
#10;x=-98410000;
#10;x=-98400000;
#10;x=-98390000;
#10;x=-98380000;
#10;x=-98370000;
#10;x=-98360000;
#10;x=-98350000;
#10;x=-98340000;
#10;x=-98330000;
#10;x=-98320000;
#10;x=-98310000;
#10;x=-98300000;
#10;x=-98290000;
#10;x=-98280000;
#10;x=-98270000;
#10;x=-98260000;
#10;x=-98250000;
#10;x=-98240000;
#10;x=-98230000;
#10;x=-98220000;
#10;x=-98210000;
#10;x=-98200000;
#10;x=-98190000;
#10;x=-98180000;
#10;x=-98170000;
#10;x=-98160000;
#10;x=-98150000;
#10;x=-98140000;
#10;x=-98130000;
#10;x=-98120000;
#10;x=-98110000;
#10;x=-98100000;
#10;x=-98090000;
#10;x=-98080000;
#10;x=-98070000;
#10;x=-98060000;
#10;x=-98050000;
#10;x=-98040000;
#10;x=-98030000;
#10;x=-98020000;
#10;x=-98010000;
#10;x=-98000000;
#10;x=-97990000;
#10;x=-97980000;
#10;x=-97970000;
#10;x=-97960000;
#10;x=-97950000;
#10;x=-97940000;
#10;x=-97930000;
#10;x=-97920000;
#10;x=-97910000;
#10;x=-97900000;
#10;x=-97890000;
#10;x=-97880000;
#10;x=-97870000;
#10;x=-97860000;
#10;x=-97850000;
#10;x=-97840000;
#10;x=-97830000;
#10;x=-97820000;
#10;x=-97810000;
#10;x=-97800000;
#10;x=-97790000;
#10;x=-97780000;
#10;x=-97770000;
#10;x=-97760000;
#10;x=-97750000;
#10;x=-97740000;
#10;x=-97730000;
#10;x=-97720000;
#10;x=-97710000;
#10;x=-97700000;
#10;x=-97690000;
#10;x=-97680000;
#10;x=-97670000;
#10;x=-97660000;
#10;x=-97650000;
#10;x=-97640000;
#10;x=-97630000;
#10;x=-97620000;
#10;x=-97610000;
#10;x=-97600000;
#10;x=-97590000;
#10;x=-97580000;
#10;x=-97570000;
#10;x=-97560000;
#10;x=-97550000;
#10;x=-97540000;
#10;x=-97530000;
#10;x=-97520000;
#10;x=-97510000;
#10;x=-97500000;
#10;x=-97490000;
#10;x=-97480000;
#10;x=-97470000;
#10;x=-97460000;
#10;x=-97450000;
#10;x=-97440000;
#10;x=-97430000;
#10;x=-97420000;
#10;x=-97410000;
#10;x=-97400000;
#10;x=-97390000;
#10;x=-97380000;
#10;x=-97370000;
#10;x=-97360000;
#10;x=-97350000;
#10;x=-97340000;
#10;x=-97330000;
#10;x=-97320000;
#10;x=-97310000;
#10;x=-97300000;
#10;x=-97290000;
#10;x=-97280000;
#10;x=-97270000;
#10;x=-97260000;
#10;x=-97250000;
#10;x=-97240000;
#10;x=-97230000;
#10;x=-97220000;
#10;x=-97210000;
#10;x=-97200000;
#10;x=-97190000;
#10;x=-97180000;
#10;x=-97170000;
#10;x=-97160000;
#10;x=-97150000;
#10;x=-97140000;
#10;x=-97130000;
#10;x=-97120000;
#10;x=-97110000;
#10;x=-97100000;
#10;x=-97090000;
#10;x=-97080000;
#10;x=-97070000;
#10;x=-97060000;
#10;x=-97050000;
#10;x=-97040000;
#10;x=-97030000;
#10;x=-97020000;
#10;x=-97010000;
#10;x=-97000000;
#10;x=-96990000;
#10;x=-96980000;
#10;x=-96970000;
#10;x=-96960000;
#10;x=-96950000;
#10;x=-96940000;
#10;x=-96930000;
#10;x=-96920000;
#10;x=-96910000;
#10;x=-96900000;
#10;x=-96890000;
#10;x=-96880000;
#10;x=-96870000;
#10;x=-96860000;
#10;x=-96850000;
#10;x=-96840000;
#10;x=-96830000;
#10;x=-96820000;
#10;x=-96810000;
#10;x=-96800000;
#10;x=-96790000;
#10;x=-96780000;
#10;x=-96770000;
#10;x=-96760000;
#10;x=-96750000;
#10;x=-96740000;
#10;x=-96730000;
#10;x=-96720000;
#10;x=-96710000;
#10;x=-96700000;
#10;x=-96690000;
#10;x=-96680000;
#10;x=-96670000;
#10;x=-96660000;
#10;x=-96650000;
#10;x=-96640000;
#10;x=-96630000;
#10;x=-96620000;
#10;x=-96610000;
#10;x=-96600000;
#10;x=-96590000;
#10;x=-96580000;
#10;x=-96570000;
#10;x=-96560000;
#10;x=-96550000;
#10;x=-96540000;
#10;x=-96530000;
#10;x=-96520000;
#10;x=-96510000;
#10;x=-96500000;
#10;x=-96490000;
#10;x=-96480000;
#10;x=-96470000;
#10;x=-96460000;
#10;x=-96450000;
#10;x=-96440000;
#10;x=-96430000;
#10;x=-96420000;
#10;x=-96410000;
#10;x=-96400000;
#10;x=-96390000;
#10;x=-96380000;
#10;x=-96370000;
#10;x=-96360000;
#10;x=-96350000;
#10;x=-96340000;
#10;x=-96330000;
#10;x=-96320000;
#10;x=-96310000;
#10;x=-96300000;
#10;x=-96290000;
#10;x=-96280000;
#10;x=-96270000;
#10;x=-96260000;
#10;x=-96250000;
#10;x=-96240000;
#10;x=-96230000;
#10;x=-96220000;
#10;x=-96210000;
#10;x=-96200000;
#10;x=-96190000;
#10;x=-96180000;
#10;x=-96170000;
#10;x=-96160000;
#10;x=-96150000;
#10;x=-96140000;
#10;x=-96130000;
#10;x=-96120000;
#10;x=-96110000;
#10;x=-96100000;
#10;x=-96090000;
#10;x=-96080000;
#10;x=-96070000;
#10;x=-96060000;
#10;x=-96050000;
#10;x=-96040000;
#10;x=-96030000;
#10;x=-96020000;
#10;x=-96010000;
#10;x=-96000000;
#10;x=-95990000;
#10;x=-95980000;
#10;x=-95970000;
#10;x=-95960000;
#10;x=-95950000;
#10;x=-95940000;
#10;x=-95930000;
#10;x=-95920000;
#10;x=-95910000;
#10;x=-95900000;
#10;x=-95890000;
#10;x=-95880000;
#10;x=-95870000;
#10;x=-95860000;
#10;x=-95850000;
#10;x=-95840000;
#10;x=-95830000;
#10;x=-95820000;
#10;x=-95810000;
#10;x=-95800000;
#10;x=-95790000;
#10;x=-95780000;
#10;x=-95770000;
#10;x=-95760000;
#10;x=-95750000;
#10;x=-95740000;
#10;x=-95730000;
#10;x=-95720000;
#10;x=-95710000;
#10;x=-95700000;
#10;x=-95690000;
#10;x=-95680000;
#10;x=-95670000;
#10;x=-95660000;
#10;x=-95650000;
#10;x=-95640000;
#10;x=-95630000;
#10;x=-95620000;
#10;x=-95610000;
#10;x=-95600000;
#10;x=-95590000;
#10;x=-95580000;
#10;x=-95570000;
#10;x=-95560000;
#10;x=-95550000;
#10;x=-95540000;
#10;x=-95530000;
#10;x=-95520000;
#10;x=-95510000;
#10;x=-95500000;
#10;x=-95490000;
#10;x=-95480000;
#10;x=-95470000;
#10;x=-95460000;
#10;x=-95450000;
#10;x=-95440000;
#10;x=-95430000;
#10;x=-95420000;
#10;x=-95410000;
#10;x=-95400000;
#10;x=-95390000;
#10;x=-95380000;
#10;x=-95370000;
#10;x=-95360000;
#10;x=-95350000;
#10;x=-95340000;
#10;x=-95330000;
#10;x=-95320000;
#10;x=-95310000;
#10;x=-95300000;
#10;x=-95290000;
#10;x=-95280000;
#10;x=-95270000;
#10;x=-95260000;
#10;x=-95250000;
#10;x=-95240000;
#10;x=-95230000;
#10;x=-95220000;
#10;x=-95210000;
#10;x=-95200000;
#10;x=-95190000;
#10;x=-95180000;
#10;x=-95170000;
#10;x=-95160000;
#10;x=-95150000;
#10;x=-95140000;
#10;x=-95130000;
#10;x=-95120000;
#10;x=-95110000;
#10;x=-95100000;
#10;x=-95090000;
#10;x=-95080000;
#10;x=-95070000;
#10;x=-95060000;
#10;x=-95050000;
#10;x=-95040000;
#10;x=-95030000;
#10;x=-95020000;
#10;x=-95010000;
#10;x=-95000000;
#10;x=-94990000;
#10;x=-94980000;
#10;x=-94970000;
#10;x=-94960000;
#10;x=-94950000;
#10;x=-94940000;
#10;x=-94930000;
#10;x=-94920000;
#10;x=-94910000;
#10;x=-94900000;
#10;x=-94890000;
#10;x=-94880000;
#10;x=-94870000;
#10;x=-94860000;
#10;x=-94850000;
#10;x=-94840000;
#10;x=-94830000;
#10;x=-94820000;
#10;x=-94810000;
#10;x=-94800000;
#10;x=-94790000;
#10;x=-94780000;
#10;x=-94770000;
#10;x=-94760000;
#10;x=-94750000;
#10;x=-94740000;
#10;x=-94730000;
#10;x=-94720000;
#10;x=-94710000;
#10;x=-94700000;
#10;x=-94690000;
#10;x=-94680000;
#10;x=-94670000;
#10;x=-94660000;
#10;x=-94650000;
#10;x=-94640000;
#10;x=-94630000;
#10;x=-94620000;
#10;x=-94610000;
#10;x=-94600000;
#10;x=-94590000;
#10;x=-94580000;
#10;x=-94570000;
#10;x=-94560000;
#10;x=-94550000;
#10;x=-94540000;
#10;x=-94530000;
#10;x=-94520000;
#10;x=-94510000;
#10;x=-94500000;
#10;x=-94490000;
#10;x=-94480000;
#10;x=-94470000;
#10;x=-94460000;
#10;x=-94450000;
#10;x=-94440000;
#10;x=-94430000;
#10;x=-94420000;
#10;x=-94410000;
#10;x=-94400000;
#10;x=-94390000;
#10;x=-94380000;
#10;x=-94370000;
#10;x=-94360000;
#10;x=-94350000;
#10;x=-94340000;
#10;x=-94330000;
#10;x=-94320000;
#10;x=-94310000;
#10;x=-94300000;
#10;x=-94290000;
#10;x=-94280000;
#10;x=-94270000;
#10;x=-94260000;
#10;x=-94250000;
#10;x=-94240000;
#10;x=-94230000;
#10;x=-94220000;
#10;x=-94210000;
#10;x=-94200000;
#10;x=-94190000;
#10;x=-94180000;
#10;x=-94170000;
#10;x=-94160000;
#10;x=-94150000;
#10;x=-94140000;
#10;x=-94130000;
#10;x=-94120000;
#10;x=-94110000;
#10;x=-94100000;
#10;x=-94090000;
#10;x=-94080000;
#10;x=-94070000;
#10;x=-94060000;
#10;x=-94050000;
#10;x=-94040000;
#10;x=-94030000;
#10;x=-94020000;
#10;x=-94010000;
#10;x=-94000000;
#10;x=-93990000;
#10;x=-93980000;
#10;x=-93970000;
#10;x=-93960000;
#10;x=-93950000;
#10;x=-93940000;
#10;x=-93930000;
#10;x=-93920000;
#10;x=-93910000;
#10;x=-93900000;
#10;x=-93890000;
#10;x=-93880000;
#10;x=-93870000;
#10;x=-93860000;
#10;x=-93850000;
#10;x=-93840000;
#10;x=-93830000;
#10;x=-93820000;
#10;x=-93810000;
#10;x=-93800000;
#10;x=-93790000;
#10;x=-93780000;
#10;x=-93770000;
#10;x=-93760000;
#10;x=-93750000;
#10;x=-93740000;
#10;x=-93730000;
#10;x=-93720000;
#10;x=-93710000;
#10;x=-93700000;
#10;x=-93690000;
#10;x=-93680000;
#10;x=-93670000;
#10;x=-93660000;
#10;x=-93650000;
#10;x=-93640000;
#10;x=-93630000;
#10;x=-93620000;
#10;x=-93610000;
#10;x=-93600000;
#10;x=-93590000;
#10;x=-93580000;
#10;x=-93570000;
#10;x=-93560000;
#10;x=-93550000;
#10;x=-93540000;
#10;x=-93530000;
#10;x=-93520000;
#10;x=-93510000;
#10;x=-93500000;
#10;x=-93490000;
#10;x=-93480000;
#10;x=-93470000;
#10;x=-93460000;
#10;x=-93450000;
#10;x=-93440000;
#10;x=-93430000;
#10;x=-93420000;
#10;x=-93410000;
#10;x=-93400000;
#10;x=-93390000;
#10;x=-93380000;
#10;x=-93370000;
#10;x=-93360000;
#10;x=-93350000;
#10;x=-93340000;
#10;x=-93330000;
#10;x=-93320000;
#10;x=-93310000;
#10;x=-93300000;
#10;x=-93290000;
#10;x=-93280000;
#10;x=-93270000;
#10;x=-93260000;
#10;x=-93250000;
#10;x=-93240000;
#10;x=-93230000;
#10;x=-93220000;
#10;x=-93210000;
#10;x=-93200000;
#10;x=-93190000;
#10;x=-93180000;
#10;x=-93170000;
#10;x=-93160000;
#10;x=-93150000;
#10;x=-93140000;
#10;x=-93130000;
#10;x=-93120000;
#10;x=-93110000;
#10;x=-93100000;
#10;x=-93090000;
#10;x=-93080000;
#10;x=-93070000;
#10;x=-93060000;
#10;x=-93050000;
#10;x=-93040000;
#10;x=-93030000;
#10;x=-93020000;
#10;x=-93010000;
#10;x=-93000000;
#10;x=-92990000;
#10;x=-92980000;
#10;x=-92970000;
#10;x=-92960000;
#10;x=-92950000;
#10;x=-92940000;
#10;x=-92930000;
#10;x=-92920000;
#10;x=-92910000;
#10;x=-92900000;
#10;x=-92890000;
#10;x=-92880000;
#10;x=-92870000;
#10;x=-92860000;
#10;x=-92850000;
#10;x=-92840000;
#10;x=-92830000;
#10;x=-92820000;
#10;x=-92810000;
#10;x=-92800000;
#10;x=-92790000;
#10;x=-92780000;
#10;x=-92770000;
#10;x=-92760000;
#10;x=-92750000;
#10;x=-92740000;
#10;x=-92730000;
#10;x=-92720000;
#10;x=-92710000;
#10;x=-92700000;
#10;x=-92690000;
#10;x=-92680000;
#10;x=-92670000;
#10;x=-92660000;
#10;x=-92650000;
#10;x=-92640000;
#10;x=-92630000;
#10;x=-92620000;
#10;x=-92610000;
#10;x=-92600000;
#10;x=-92590000;
#10;x=-92580000;
#10;x=-92570000;
#10;x=-92560000;
#10;x=-92550000;
#10;x=-92540000;
#10;x=-92530000;
#10;x=-92520000;
#10;x=-92510000;
#10;x=-92500000;
#10;x=-92490000;
#10;x=-92480000;
#10;x=-92470000;
#10;x=-92460000;
#10;x=-92450000;
#10;x=-92440000;
#10;x=-92430000;
#10;x=-92420000;
#10;x=-92410000;
#10;x=-92400000;
#10;x=-92390000;
#10;x=-92380000;
#10;x=-92370000;
#10;x=-92360000;
#10;x=-92350000;
#10;x=-92340000;
#10;x=-92330000;
#10;x=-92320000;
#10;x=-92310000;
#10;x=-92300000;
#10;x=-92290000;
#10;x=-92280000;
#10;x=-92270000;
#10;x=-92260000;
#10;x=-92250000;
#10;x=-92240000;
#10;x=-92230000;
#10;x=-92220000;
#10;x=-92210000;
#10;x=-92200000;
#10;x=-92190000;
#10;x=-92180000;
#10;x=-92170000;
#10;x=-92160000;
#10;x=-92150000;
#10;x=-92140000;
#10;x=-92130000;
#10;x=-92120000;
#10;x=-92110000;
#10;x=-92100000;
#10;x=-92090000;
#10;x=-92080000;
#10;x=-92070000;
#10;x=-92060000;
#10;x=-92050000;
#10;x=-92040000;
#10;x=-92030000;
#10;x=-92020000;
#10;x=-92010000;
#10;x=-92000000;
#10;x=-91990000;
#10;x=-91980000;
#10;x=-91970000;
#10;x=-91960000;
#10;x=-91950000;
#10;x=-91940000;
#10;x=-91930000;
#10;x=-91920000;
#10;x=-91910000;
#10;x=-91900000;
#10;x=-91890000;
#10;x=-91880000;
#10;x=-91870000;
#10;x=-91860000;
#10;x=-91850000;
#10;x=-91840000;
#10;x=-91830000;
#10;x=-91820000;
#10;x=-91810000;
#10;x=-91800000;
#10;x=-91790000;
#10;x=-91780000;
#10;x=-91770000;
#10;x=-91760000;
#10;x=-91750000;
#10;x=-91740000;
#10;x=-91730000;
#10;x=-91720000;
#10;x=-91710000;
#10;x=-91700000;
#10;x=-91690000;
#10;x=-91680000;
#10;x=-91670000;
#10;x=-91660000;
#10;x=-91650000;
#10;x=-91640000;
#10;x=-91630000;
#10;x=-91620000;
#10;x=-91610000;
#10;x=-91600000;
#10;x=-91590000;
#10;x=-91580000;
#10;x=-91570000;
#10;x=-91560000;
#10;x=-91550000;
#10;x=-91540000;
#10;x=-91530000;
#10;x=-91520000;
#10;x=-91510000;
#10;x=-91500000;
#10;x=-91490000;
#10;x=-91480000;
#10;x=-91470000;
#10;x=-91460000;
#10;x=-91450000;
#10;x=-91440000;
#10;x=-91430000;
#10;x=-91420000;
#10;x=-91410000;
#10;x=-91400000;
#10;x=-91390000;
#10;x=-91380000;
#10;x=-91370000;
#10;x=-91360000;
#10;x=-91350000;
#10;x=-91340000;
#10;x=-91330000;
#10;x=-91320000;
#10;x=-91310000;
#10;x=-91300000;
#10;x=-91290000;
#10;x=-91280000;
#10;x=-91270000;
#10;x=-91260000;
#10;x=-91250000;
#10;x=-91240000;
#10;x=-91230000;
#10;x=-91220000;
#10;x=-91210000;
#10;x=-91200000;
#10;x=-91190000;
#10;x=-91180000;
#10;x=-91170000;
#10;x=-91160000;
#10;x=-91150000;
#10;x=-91140000;
#10;x=-91130000;
#10;x=-91120000;
#10;x=-91110000;
#10;x=-91100000;
#10;x=-91090000;
#10;x=-91080000;
#10;x=-91070000;
#10;x=-91060000;
#10;x=-91050000;
#10;x=-91040000;
#10;x=-91030000;
#10;x=-91020000;
#10;x=-91010000;
#10;x=-91000000;
#10;x=-90990000;
#10;x=-90980000;
#10;x=-90970000;
#10;x=-90960000;
#10;x=-90950000;
#10;x=-90940000;
#10;x=-90930000;
#10;x=-90920000;
#10;x=-90910000;
#10;x=-90900000;
#10;x=-90890000;
#10;x=-90880000;
#10;x=-90870000;
#10;x=-90860000;
#10;x=-90850000;
#10;x=-90840000;
#10;x=-90830000;
#10;x=-90820000;
#10;x=-90810000;
#10;x=-90800000;
#10;x=-90790000;
#10;x=-90780000;
#10;x=-90770000;
#10;x=-90760000;
#10;x=-90750000;
#10;x=-90740000;
#10;x=-90730000;
#10;x=-90720000;
#10;x=-90710000;
#10;x=-90700000;
#10;x=-90690000;
#10;x=-90680000;
#10;x=-90670000;
#10;x=-90660000;
#10;x=-90650000;
#10;x=-90640000;
#10;x=-90630000;
#10;x=-90620000;
#10;x=-90610000;
#10;x=-90600000;
#10;x=-90590000;
#10;x=-90580000;
#10;x=-90570000;
#10;x=-90560000;
#10;x=-90550000;
#10;x=-90540000;
#10;x=-90530000;
#10;x=-90520000;
#10;x=-90510000;
#10;x=-90500000;
#10;x=-90490000;
#10;x=-90480000;
#10;x=-90470000;
#10;x=-90460000;
#10;x=-90450000;
#10;x=-90440000;
#10;x=-90430000;
#10;x=-90420000;
#10;x=-90410000;
#10;x=-90400000;
#10;x=-90390000;
#10;x=-90380000;
#10;x=-90370000;
#10;x=-90360000;
#10;x=-90350000;
#10;x=-90340000;
#10;x=-90330000;
#10;x=-90320000;
#10;x=-90310000;
#10;x=-90300000;
#10;x=-90290000;
#10;x=-90280000;
#10;x=-90270000;
#10;x=-90260000;
#10;x=-90250000;
#10;x=-90240000;
#10;x=-90230000;
#10;x=-90220000;
#10;x=-90210000;
#10;x=-90200000;
#10;x=-90190000;
#10;x=-90180000;
#10;x=-90170000;
#10;x=-90160000;
#10;x=-90150000;
#10;x=-90140000;
#10;x=-90130000;
#10;x=-90120000;
#10;x=-90110000;
#10;x=-90100000;
#10;x=-90090000;
#10;x=-90080000;
#10;x=-90070000;
#10;x=-90060000;
#10;x=-90050000;
#10;x=-90040000;
#10;x=-90030000;
#10;x=-90020000;
#10;x=-90010000;
#10;x=-90000000;
#10;x=-89990000;
#10;x=-89980000;
#10;x=-89970000;
#10;x=-89960000;
#10;x=-89950000;
#10;x=-89940000;
#10;x=-89930000;
#10;x=-89920000;
#10;x=-89910000;
#10;x=-89900000;
#10;x=-89890000;
#10;x=-89880000;
#10;x=-89870000;
#10;x=-89860000;
#10;x=-89850000;
#10;x=-89840000;
#10;x=-89830000;
#10;x=-89820000;
#10;x=-89810000;
#10;x=-89800000;
#10;x=-89790000;
#10;x=-89780000;
#10;x=-89770000;
#10;x=-89760000;
#10;x=-89750000;
#10;x=-89740000;
#10;x=-89730000;
#10;x=-89720000;
#10;x=-89710000;
#10;x=-89700000;
#10;x=-89690000;
#10;x=-89680000;
#10;x=-89670000;
#10;x=-89660000;
#10;x=-89650000;
#10;x=-89640000;
#10;x=-89630000;
#10;x=-89620000;
#10;x=-89610000;
#10;x=-89600000;
#10;x=-89590000;
#10;x=-89580000;
#10;x=-89570000;
#10;x=-89560000;
#10;x=-89550000;
#10;x=-89540000;
#10;x=-89530000;
#10;x=-89520000;
#10;x=-89510000;
#10;x=-89500000;
#10;x=-89490000;
#10;x=-89480000;
#10;x=-89470000;
#10;x=-89460000;
#10;x=-89450000;
#10;x=-89440000;
#10;x=-89430000;
#10;x=-89420000;
#10;x=-89410000;
#10;x=-89400000;
#10;x=-89390000;
#10;x=-89380000;
#10;x=-89370000;
#10;x=-89360000;
#10;x=-89350000;
#10;x=-89340000;
#10;x=-89330000;
#10;x=-89320000;
#10;x=-89310000;
#10;x=-89300000;
#10;x=-89290000;
#10;x=-89280000;
#10;x=-89270000;
#10;x=-89260000;
#10;x=-89250000;
#10;x=-89240000;
#10;x=-89230000;
#10;x=-89220000;
#10;x=-89210000;
#10;x=-89200000;
#10;x=-89190000;
#10;x=-89180000;
#10;x=-89170000;
#10;x=-89160000;
#10;x=-89150000;
#10;x=-89140000;
#10;x=-89130000;
#10;x=-89120000;
#10;x=-89110000;
#10;x=-89100000;
#10;x=-89090000;
#10;x=-89080000;
#10;x=-89070000;
#10;x=-89060000;
#10;x=-89050000;
#10;x=-89040000;
#10;x=-89030000;
#10;x=-89020000;
#10;x=-89010000;
#10;x=-89000000;
#10;x=-88990000;
#10;x=-88980000;
#10;x=-88970000;
#10;x=-88960000;
#10;x=-88950000;
#10;x=-88940000;
#10;x=-88930000;
#10;x=-88920000;
#10;x=-88910000;
#10;x=-88900000;
#10;x=-88890000;
#10;x=-88880000;
#10;x=-88870000;
#10;x=-88860000;
#10;x=-88850000;
#10;x=-88840000;
#10;x=-88830000;
#10;x=-88820000;
#10;x=-88810000;
#10;x=-88800000;
#10;x=-88790000;
#10;x=-88780000;
#10;x=-88770000;
#10;x=-88760000;
#10;x=-88750000;
#10;x=-88740000;
#10;x=-88730000;
#10;x=-88720000;
#10;x=-88710000;
#10;x=-88700000;
#10;x=-88690000;
#10;x=-88680000;
#10;x=-88670000;
#10;x=-88660000;
#10;x=-88650000;
#10;x=-88640000;
#10;x=-88630000;
#10;x=-88620000;
#10;x=-88610000;
#10;x=-88600000;
#10;x=-88590000;
#10;x=-88580000;
#10;x=-88570000;
#10;x=-88560000;
#10;x=-88550000;
#10;x=-88540000;
#10;x=-88530000;
#10;x=-88520000;
#10;x=-88510000;
#10;x=-88500000;
#10;x=-88490000;
#10;x=-88480000;
#10;x=-88470000;
#10;x=-88460000;
#10;x=-88450000;
#10;x=-88440000;
#10;x=-88430000;
#10;x=-88420000;
#10;x=-88410000;
#10;x=-88400000;
#10;x=-88390000;
#10;x=-88380000;
#10;x=-88370000;
#10;x=-88360000;
#10;x=-88350000;
#10;x=-88340000;
#10;x=-88330000;
#10;x=-88320000;
#10;x=-88310000;
#10;x=-88300000;
#10;x=-88290000;
#10;x=-88280000;
#10;x=-88270000;
#10;x=-88260000;
#10;x=-88250000;
#10;x=-88240000;
#10;x=-88230000;
#10;x=-88220000;
#10;x=-88210000;
#10;x=-88200000;
#10;x=-88190000;
#10;x=-88180000;
#10;x=-88170000;
#10;x=-88160000;
#10;x=-88150000;
#10;x=-88140000;
#10;x=-88130000;
#10;x=-88120000;
#10;x=-88110000;
#10;x=-88100000;
#10;x=-88090000;
#10;x=-88080000;
#10;x=-88070000;
#10;x=-88060000;
#10;x=-88050000;
#10;x=-88040000;
#10;x=-88030000;
#10;x=-88020000;
#10;x=-88010000;
#10;x=-88000000;
#10;x=-87990000;
#10;x=-87980000;
#10;x=-87970000;
#10;x=-87960000;
#10;x=-87950000;
#10;x=-87940000;
#10;x=-87930000;
#10;x=-87920000;
#10;x=-87910000;
#10;x=-87900000;
#10;x=-87890000;
#10;x=-87880000;
#10;x=-87870000;
#10;x=-87860000;
#10;x=-87850000;
#10;x=-87840000;
#10;x=-87830000;
#10;x=-87820000;
#10;x=-87810000;
#10;x=-87800000;
#10;x=-87790000;
#10;x=-87780000;
#10;x=-87770000;
#10;x=-87760000;
#10;x=-87750000;
#10;x=-87740000;
#10;x=-87730000;
#10;x=-87720000;
#10;x=-87710000;
#10;x=-87700000;
#10;x=-87690000;
#10;x=-87680000;
#10;x=-87670000;
#10;x=-87660000;
#10;x=-87650000;
#10;x=-87640000;
#10;x=-87630000;
#10;x=-87620000;
#10;x=-87610000;
#10;x=-87600000;
#10;x=-87590000;
#10;x=-87580000;
#10;x=-87570000;
#10;x=-87560000;
#10;x=-87550000;
#10;x=-87540000;
#10;x=-87530000;
#10;x=-87520000;
#10;x=-87510000;
#10;x=-87500000;
#10;x=-87490000;
#10;x=-87480000;
#10;x=-87470000;
#10;x=-87460000;
#10;x=-87450000;
#10;x=-87440000;
#10;x=-87430000;
#10;x=-87420000;
#10;x=-87410000;
#10;x=-87400000;
#10;x=-87390000;
#10;x=-87380000;
#10;x=-87370000;
#10;x=-87360000;
#10;x=-87350000;
#10;x=-87340000;
#10;x=-87330000;
#10;x=-87320000;
#10;x=-87310000;
#10;x=-87300000;
#10;x=-87290000;
#10;x=-87280000;
#10;x=-87270000;
#10;x=-87260000;
#10;x=-87250000;
#10;x=-87240000;
#10;x=-87230000;
#10;x=-87220000;
#10;x=-87210000;
#10;x=-87200000;
#10;x=-87190000;
#10;x=-87180000;
#10;x=-87170000;
#10;x=-87160000;
#10;x=-87150000;
#10;x=-87140000;
#10;x=-87130000;
#10;x=-87120000;
#10;x=-87110000;
#10;x=-87100000;
#10;x=-87090000;
#10;x=-87080000;
#10;x=-87070000;
#10;x=-87060000;
#10;x=-87050000;
#10;x=-87040000;
#10;x=-87030000;
#10;x=-87020000;
#10;x=-87010000;
#10;x=-87000000;
#10;x=-86990000;
#10;x=-86980000;
#10;x=-86970000;
#10;x=-86960000;
#10;x=-86950000;
#10;x=-86940000;
#10;x=-86930000;
#10;x=-86920000;
#10;x=-86910000;
#10;x=-86900000;
#10;x=-86890000;
#10;x=-86880000;
#10;x=-86870000;
#10;x=-86860000;
#10;x=-86850000;
#10;x=-86840000;
#10;x=-86830000;
#10;x=-86820000;
#10;x=-86810000;
#10;x=-86800000;
#10;x=-86790000;
#10;x=-86780000;
#10;x=-86770000;
#10;x=-86760000;
#10;x=-86750000;
#10;x=-86740000;
#10;x=-86730000;
#10;x=-86720000;
#10;x=-86710000;
#10;x=-86700000;
#10;x=-86690000;
#10;x=-86680000;
#10;x=-86670000;
#10;x=-86660000;
#10;x=-86650000;
#10;x=-86640000;
#10;x=-86630000;
#10;x=-86620000;
#10;x=-86610000;
#10;x=-86600000;
#10;x=-86590000;
#10;x=-86580000;
#10;x=-86570000;
#10;x=-86560000;
#10;x=-86550000;
#10;x=-86540000;
#10;x=-86530000;
#10;x=-86520000;
#10;x=-86510000;
#10;x=-86500000;
#10;x=-86490000;
#10;x=-86480000;
#10;x=-86470000;
#10;x=-86460000;
#10;x=-86450000;
#10;x=-86440000;
#10;x=-86430000;
#10;x=-86420000;
#10;x=-86410000;
#10;x=-86400000;
#10;x=-86390000;
#10;x=-86380000;
#10;x=-86370000;
#10;x=-86360000;
#10;x=-86350000;
#10;x=-86340000;
#10;x=-86330000;
#10;x=-86320000;
#10;x=-86310000;
#10;x=-86300000;
#10;x=-86290000;
#10;x=-86280000;
#10;x=-86270000;
#10;x=-86260000;
#10;x=-86250000;
#10;x=-86240000;
#10;x=-86230000;
#10;x=-86220000;
#10;x=-86210000;
#10;x=-86200000;
#10;x=-86190000;
#10;x=-86180000;
#10;x=-86170000;
#10;x=-86160000;
#10;x=-86150000;
#10;x=-86140000;
#10;x=-86130000;
#10;x=-86120000;
#10;x=-86110000;
#10;x=-86100000;
#10;x=-86090000;
#10;x=-86080000;
#10;x=-86070000;
#10;x=-86060000;
#10;x=-86050000;
#10;x=-86040000;
#10;x=-86030000;
#10;x=-86020000;
#10;x=-86010000;
#10;x=-86000000;
#10;x=-85990000;
#10;x=-85980000;
#10;x=-85970000;
#10;x=-85960000;
#10;x=-85950000;
#10;x=-85940000;
#10;x=-85930000;
#10;x=-85920000;
#10;x=-85910000;
#10;x=-85900000;
#10;x=-85890000;
#10;x=-85880000;
#10;x=-85870000;
#10;x=-85860000;
#10;x=-85850000;
#10;x=-85840000;
#10;x=-85830000;
#10;x=-85820000;
#10;x=-85810000;
#10;x=-85800000;
#10;x=-85790000;
#10;x=-85780000;
#10;x=-85770000;
#10;x=-85760000;
#10;x=-85750000;
#10;x=-85740000;
#10;x=-85730000;
#10;x=-85720000;
#10;x=-85710000;
#10;x=-85700000;
#10;x=-85690000;
#10;x=-85680000;
#10;x=-85670000;
#10;x=-85660000;
#10;x=-85650000;
#10;x=-85640000;
#10;x=-85630000;
#10;x=-85620000;
#10;x=-85610000;
#10;x=-85600000;
#10;x=-85590000;
#10;x=-85580000;
#10;x=-85570000;
#10;x=-85560000;
#10;x=-85550000;
#10;x=-85540000;
#10;x=-85530000;
#10;x=-85520000;
#10;x=-85510000;
#10;x=-85500000;
#10;x=-85490000;
#10;x=-85480000;
#10;x=-85470000;
#10;x=-85460000;
#10;x=-85450000;
#10;x=-85440000;
#10;x=-85430000;
#10;x=-85420000;
#10;x=-85410000;
#10;x=-85400000;
#10;x=-85390000;
#10;x=-85380000;
#10;x=-85370000;
#10;x=-85360000;
#10;x=-85350000;
#10;x=-85340000;
#10;x=-85330000;
#10;x=-85320000;
#10;x=-85310000;
#10;x=-85300000;
#10;x=-85290000;
#10;x=-85280000;
#10;x=-85270000;
#10;x=-85260000;
#10;x=-85250000;
#10;x=-85240000;
#10;x=-85230000;
#10;x=-85220000;
#10;x=-85210000;
#10;x=-85200000;
#10;x=-85190000;
#10;x=-85180000;
#10;x=-85170000;
#10;x=-85160000;
#10;x=-85150000;
#10;x=-85140000;
#10;x=-85130000;
#10;x=-85120000;
#10;x=-85110000;
#10;x=-85100000;
#10;x=-85090000;
#10;x=-85080000;
#10;x=-85070000;
#10;x=-85060000;
#10;x=-85050000;
#10;x=-85040000;
#10;x=-85030000;
#10;x=-85020000;
#10;x=-85010000;
#10;x=-85000000;
#10;x=-84990000;
#10;x=-84980000;
#10;x=-84970000;
#10;x=-84960000;
#10;x=-84950000;
#10;x=-84940000;
#10;x=-84930000;
#10;x=-84920000;
#10;x=-84910000;
#10;x=-84900000;
#10;x=-84890000;
#10;x=-84880000;
#10;x=-84870000;
#10;x=-84860000;
#10;x=-84850000;
#10;x=-84840000;
#10;x=-84830000;
#10;x=-84820000;
#10;x=-84810000;
#10;x=-84800000;
#10;x=-84790000;
#10;x=-84780000;
#10;x=-84770000;
#10;x=-84760000;
#10;x=-84750000;
#10;x=-84740000;
#10;x=-84730000;
#10;x=-84720000;
#10;x=-84710000;
#10;x=-84700000;
#10;x=-84690000;
#10;x=-84680000;
#10;x=-84670000;
#10;x=-84660000;
#10;x=-84650000;
#10;x=-84640000;
#10;x=-84630000;
#10;x=-84620000;
#10;x=-84610000;
#10;x=-84600000;
#10;x=-84590000;
#10;x=-84580000;
#10;x=-84570000;
#10;x=-84560000;
#10;x=-84550000;
#10;x=-84540000;
#10;x=-84530000;
#10;x=-84520000;
#10;x=-84510000;
#10;x=-84500000;
#10;x=-84490000;
#10;x=-84480000;
#10;x=-84470000;
#10;x=-84460000;
#10;x=-84450000;
#10;x=-84440000;
#10;x=-84430000;
#10;x=-84420000;
#10;x=-84410000;
#10;x=-84400000;
#10;x=-84390000;
#10;x=-84380000;
#10;x=-84370000;
#10;x=-84360000;
#10;x=-84350000;
#10;x=-84340000;
#10;x=-84330000;
#10;x=-84320000;
#10;x=-84310000;
#10;x=-84300000;
#10;x=-84290000;
#10;x=-84280000;
#10;x=-84270000;
#10;x=-84260000;
#10;x=-84250000;
#10;x=-84240000;
#10;x=-84230000;
#10;x=-84220000;
#10;x=-84210000;
#10;x=-84200000;
#10;x=-84190000;
#10;x=-84180000;
#10;x=-84170000;
#10;x=-84160000;
#10;x=-84150000;
#10;x=-84140000;
#10;x=-84130000;
#10;x=-84120000;
#10;x=-84110000;
#10;x=-84100000;
#10;x=-84090000;
#10;x=-84080000;
#10;x=-84070000;
#10;x=-84060000;
#10;x=-84050000;
#10;x=-84040000;
#10;x=-84030000;
#10;x=-84020000;
#10;x=-84010000;
#10;x=-84000000;
#10;x=-83990000;
#10;x=-83980000;
#10;x=-83970000;
#10;x=-83960000;
#10;x=-83950000;
#10;x=-83940000;
#10;x=-83930000;
#10;x=-83920000;
#10;x=-83910000;
#10;x=-83900000;
#10;x=-83890000;
#10;x=-83880000;
#10;x=-83870000;
#10;x=-83860000;
#10;x=-83850000;
#10;x=-83840000;
#10;x=-83830000;
#10;x=-83820000;
#10;x=-83810000;
#10;x=-83800000;
#10;x=-83790000;
#10;x=-83780000;
#10;x=-83770000;
#10;x=-83760000;
#10;x=-83750000;
#10;x=-83740000;
#10;x=-83730000;
#10;x=-83720000;
#10;x=-83710000;
#10;x=-83700000;
#10;x=-83690000;
#10;x=-83680000;
#10;x=-83670000;
#10;x=-83660000;
#10;x=-83650000;
#10;x=-83640000;
#10;x=-83630000;
#10;x=-83620000;
#10;x=-83610000;
#10;x=-83600000;
#10;x=-83590000;
#10;x=-83580000;
#10;x=-83570000;
#10;x=-83560000;
#10;x=-83550000;
#10;x=-83540000;
#10;x=-83530000;
#10;x=-83520000;
#10;x=-83510000;
#10;x=-83500000;
#10;x=-83490000;
#10;x=-83480000;
#10;x=-83470000;
#10;x=-83460000;
#10;x=-83450000;
#10;x=-83440000;
#10;x=-83430000;
#10;x=-83420000;
#10;x=-83410000;
#10;x=-83400000;
#10;x=-83390000;
#10;x=-83380000;
#10;x=-83370000;
#10;x=-83360000;
#10;x=-83350000;
#10;x=-83340000;
#10;x=-83330000;
#10;x=-83320000;
#10;x=-83310000;
#10;x=-83300000;
#10;x=-83290000;
#10;x=-83280000;
#10;x=-83270000;
#10;x=-83260000;
#10;x=-83250000;
#10;x=-83240000;
#10;x=-83230000;
#10;x=-83220000;
#10;x=-83210000;
#10;x=-83200000;
#10;x=-83190000;
#10;x=-83180000;
#10;x=-83170000;
#10;x=-83160000;
#10;x=-83150000;
#10;x=-83140000;
#10;x=-83130000;
#10;x=-83120000;
#10;x=-83110000;
#10;x=-83100000;
#10;x=-83090000;
#10;x=-83080000;
#10;x=-83070000;
#10;x=-83060000;
#10;x=-83050000;
#10;x=-83040000;
#10;x=-83030000;
#10;x=-83020000;
#10;x=-83010000;
#10;x=-83000000;
#10;x=-82990000;
#10;x=-82980000;
#10;x=-82970000;
#10;x=-82960000;
#10;x=-82950000;
#10;x=-82940000;
#10;x=-82930000;
#10;x=-82920000;
#10;x=-82910000;
#10;x=-82900000;
#10;x=-82890000;
#10;x=-82880000;
#10;x=-82870000;
#10;x=-82860000;
#10;x=-82850000;
#10;x=-82840000;
#10;x=-82830000;
#10;x=-82820000;
#10;x=-82810000;
#10;x=-82800000;
#10;x=-82790000;
#10;x=-82780000;
#10;x=-82770000;
#10;x=-82760000;
#10;x=-82750000;
#10;x=-82740000;
#10;x=-82730000;
#10;x=-82720000;
#10;x=-82710000;
#10;x=-82700000;
#10;x=-82690000;
#10;x=-82680000;
#10;x=-82670000;
#10;x=-82660000;
#10;x=-82650000;
#10;x=-82640000;
#10;x=-82630000;
#10;x=-82620000;
#10;x=-82610000;
#10;x=-82600000;
#10;x=-82590000;
#10;x=-82580000;
#10;x=-82570000;
#10;x=-82560000;
#10;x=-82550000;
#10;x=-82540000;
#10;x=-82530000;
#10;x=-82520000;
#10;x=-82510000;
#10;x=-82500000;
#10;x=-82490000;
#10;x=-82480000;
#10;x=-82470000;
#10;x=-82460000;
#10;x=-82450000;
#10;x=-82440000;
#10;x=-82430000;
#10;x=-82420000;
#10;x=-82410000;
#10;x=-82400000;
#10;x=-82390000;
#10;x=-82380000;
#10;x=-82370000;
#10;x=-82360000;
#10;x=-82350000;
#10;x=-82340000;
#10;x=-82330000;
#10;x=-82320000;
#10;x=-82310000;
#10;x=-82300000;
#10;x=-82290000;
#10;x=-82280000;
#10;x=-82270000;
#10;x=-82260000;
#10;x=-82250000;
#10;x=-82240000;
#10;x=-82230000;
#10;x=-82220000;
#10;x=-82210000;
#10;x=-82200000;
#10;x=-82190000;
#10;x=-82180000;
#10;x=-82170000;
#10;x=-82160000;
#10;x=-82150000;
#10;x=-82140000;
#10;x=-82130000;
#10;x=-82120000;
#10;x=-82110000;
#10;x=-82100000;
#10;x=-82090000;
#10;x=-82080000;
#10;x=-82070000;
#10;x=-82060000;
#10;x=-82050000;
#10;x=-82040000;
#10;x=-82030000;
#10;x=-82020000;
#10;x=-82010000;
#10;x=-82000000;
#10;x=-81990000;
#10;x=-81980000;
#10;x=-81970000;
#10;x=-81960000;
#10;x=-81950000;
#10;x=-81940000;
#10;x=-81930000;
#10;x=-81920000;
#10;x=-81910000;
#10;x=-81900000;
#10;x=-81890000;
#10;x=-81880000;
#10;x=-81870000;
#10;x=-81860000;
#10;x=-81850000;
#10;x=-81840000;
#10;x=-81830000;
#10;x=-81820000;
#10;x=-81810000;
#10;x=-81800000;
#10;x=-81790000;
#10;x=-81780000;
#10;x=-81770000;
#10;x=-81760000;
#10;x=-81750000;
#10;x=-81740000;
#10;x=-81730000;
#10;x=-81720000;
#10;x=-81710000;
#10;x=-81700000;
#10;x=-81690000;
#10;x=-81680000;
#10;x=-81670000;
#10;x=-81660000;
#10;x=-81650000;
#10;x=-81640000;
#10;x=-81630000;
#10;x=-81620000;
#10;x=-81610000;
#10;x=-81600000;
#10;x=-81590000;
#10;x=-81580000;
#10;x=-81570000;
#10;x=-81560000;
#10;x=-81550000;
#10;x=-81540000;
#10;x=-81530000;
#10;x=-81520000;
#10;x=-81510000;
#10;x=-81500000;
#10;x=-81490000;
#10;x=-81480000;
#10;x=-81470000;
#10;x=-81460000;
#10;x=-81450000;
#10;x=-81440000;
#10;x=-81430000;
#10;x=-81420000;
#10;x=-81410000;
#10;x=-81400000;
#10;x=-81390000;
#10;x=-81380000;
#10;x=-81370000;
#10;x=-81360000;
#10;x=-81350000;
#10;x=-81340000;
#10;x=-81330000;
#10;x=-81320000;
#10;x=-81310000;
#10;x=-81300000;
#10;x=-81290000;
#10;x=-81280000;
#10;x=-81270000;
#10;x=-81260000;
#10;x=-81250000;
#10;x=-81240000;
#10;x=-81230000;
#10;x=-81220000;
#10;x=-81210000;
#10;x=-81200000;
#10;x=-81190000;
#10;x=-81180000;
#10;x=-81170000;
#10;x=-81160000;
#10;x=-81150000;
#10;x=-81140000;
#10;x=-81130000;
#10;x=-81120000;
#10;x=-81110000;
#10;x=-81100000;
#10;x=-81090000;
#10;x=-81080000;
#10;x=-81070000;
#10;x=-81060000;
#10;x=-81050000;
#10;x=-81040000;
#10;x=-81030000;
#10;x=-81020000;
#10;x=-81010000;
#10;x=-81000000;
#10;x=-80990000;
#10;x=-80980000;
#10;x=-80970000;
#10;x=-80960000;
#10;x=-80950000;
#10;x=-80940000;
#10;x=-80930000;
#10;x=-80920000;
#10;x=-80910000;
#10;x=-80900000;
#10;x=-80890000;
#10;x=-80880000;
#10;x=-80870000;
#10;x=-80860000;
#10;x=-80850000;
#10;x=-80840000;
#10;x=-80830000;
#10;x=-80820000;
#10;x=-80810000;
#10;x=-80800000;
#10;x=-80790000;
#10;x=-80780000;
#10;x=-80770000;
#10;x=-80760000;
#10;x=-80750000;
#10;x=-80740000;
#10;x=-80730000;
#10;x=-80720000;
#10;x=-80710000;
#10;x=-80700000;
#10;x=-80690000;
#10;x=-80680000;
#10;x=-80670000;
#10;x=-80660000;
#10;x=-80650000;
#10;x=-80640000;
#10;x=-80630000;
#10;x=-80620000;
#10;x=-80610000;
#10;x=-80600000;
#10;x=-80590000;
#10;x=-80580000;
#10;x=-80570000;
#10;x=-80560000;
#10;x=-80550000;
#10;x=-80540000;
#10;x=-80530000;
#10;x=-80520000;
#10;x=-80510000;
#10;x=-80500000;
#10;x=-80490000;
#10;x=-80480000;
#10;x=-80470000;
#10;x=-80460000;
#10;x=-80450000;
#10;x=-80440000;
#10;x=-80430000;
#10;x=-80420000;
#10;x=-80410000;
#10;x=-80400000;
#10;x=-80390000;
#10;x=-80380000;
#10;x=-80370000;
#10;x=-80360000;
#10;x=-80350000;
#10;x=-80340000;
#10;x=-80330000;
#10;x=-80320000;
#10;x=-80310000;
#10;x=-80300000;
#10;x=-80290000;
#10;x=-80280000;
#10;x=-80270000;
#10;x=-80260000;
#10;x=-80250000;
#10;x=-80240000;
#10;x=-80230000;
#10;x=-80220000;
#10;x=-80210000;
#10;x=-80200000;
#10;x=-80190000;
#10;x=-80180000;
#10;x=-80170000;
#10;x=-80160000;
#10;x=-80150000;
#10;x=-80140000;
#10;x=-80130000;
#10;x=-80120000;
#10;x=-80110000;
#10;x=-80100000;
#10;x=-80090000;
#10;x=-80080000;
#10;x=-80070000;
#10;x=-80060000;
#10;x=-80050000;
#10;x=-80040000;
#10;x=-80030000;
#10;x=-80020000;
#10;x=-80010000;
#10;x=-80000000;
#10;x=-79990000;
#10;x=-79980000;
#10;x=-79970000;
#10;x=-79960000;
#10;x=-79950000;
#10;x=-79940000;
#10;x=-79930000;
#10;x=-79920000;
#10;x=-79910000;
#10;x=-79900000;
#10;x=-79890000;
#10;x=-79880000;
#10;x=-79870000;
#10;x=-79860000;
#10;x=-79850000;
#10;x=-79840000;
#10;x=-79830000;
#10;x=-79820000;
#10;x=-79810000;
#10;x=-79800000;
#10;x=-79790000;
#10;x=-79780000;
#10;x=-79770000;
#10;x=-79760000;
#10;x=-79750000;
#10;x=-79740000;
#10;x=-79730000;
#10;x=-79720000;
#10;x=-79710000;
#10;x=-79700000;
#10;x=-79690000;
#10;x=-79680000;
#10;x=-79670000;
#10;x=-79660000;
#10;x=-79650000;
#10;x=-79640000;
#10;x=-79630000;
#10;x=-79620000;
#10;x=-79610000;
#10;x=-79600000;
#10;x=-79590000;
#10;x=-79580000;
#10;x=-79570000;
#10;x=-79560000;
#10;x=-79550000;
#10;x=-79540000;
#10;x=-79530000;
#10;x=-79520000;
#10;x=-79510000;
#10;x=-79500000;
#10;x=-79490000;
#10;x=-79480000;
#10;x=-79470000;
#10;x=-79460000;
#10;x=-79450000;
#10;x=-79440000;
#10;x=-79430000;
#10;x=-79420000;
#10;x=-79410000;
#10;x=-79400000;
#10;x=-79390000;
#10;x=-79380000;
#10;x=-79370000;
#10;x=-79360000;
#10;x=-79350000;
#10;x=-79340000;
#10;x=-79330000;
#10;x=-79320000;
#10;x=-79310000;
#10;x=-79300000;
#10;x=-79290000;
#10;x=-79280000;
#10;x=-79270000;
#10;x=-79260000;
#10;x=-79250000;
#10;x=-79240000;
#10;x=-79230000;
#10;x=-79220000;
#10;x=-79210000;
#10;x=-79200000;
#10;x=-79190000;
#10;x=-79180000;
#10;x=-79170000;
#10;x=-79160000;
#10;x=-79150000;
#10;x=-79140000;
#10;x=-79130000;
#10;x=-79120000;
#10;x=-79110000;
#10;x=-79100000;
#10;x=-79090000;
#10;x=-79080000;
#10;x=-79070000;
#10;x=-79060000;
#10;x=-79050000;
#10;x=-79040000;
#10;x=-79030000;
#10;x=-79020000;
#10;x=-79010000;
#10;x=-79000000;
#10;x=-78990000;
#10;x=-78980000;
#10;x=-78970000;
#10;x=-78960000;
#10;x=-78950000;
#10;x=-78940000;
#10;x=-78930000;
#10;x=-78920000;
#10;x=-78910000;
#10;x=-78900000;
#10;x=-78890000;
#10;x=-78880000;
#10;x=-78870000;
#10;x=-78860000;
#10;x=-78850000;
#10;x=-78840000;
#10;x=-78830000;
#10;x=-78820000;
#10;x=-78810000;
#10;x=-78800000;
#10;x=-78790000;
#10;x=-78780000;
#10;x=-78770000;
#10;x=-78760000;
#10;x=-78750000;
#10;x=-78740000;
#10;x=-78730000;
#10;x=-78720000;
#10;x=-78710000;
#10;x=-78700000;
#10;x=-78690000;
#10;x=-78680000;
#10;x=-78670000;
#10;x=-78660000;
#10;x=-78650000;
#10;x=-78640000;
#10;x=-78630000;
#10;x=-78620000;
#10;x=-78610000;
#10;x=-78600000;
#10;x=-78590000;
#10;x=-78580000;
#10;x=-78570000;
#10;x=-78560000;
#10;x=-78550000;
#10;x=-78540000;
#10;x=-78530000;
#10;x=-78520000;
#10;x=-78510000;
#10;x=-78500000;
#10;x=-78490000;
#10;x=-78480000;
#10;x=-78470000;
#10;x=-78460000;
#10;x=-78450000;
#10;x=-78440000;
#10;x=-78430000;
#10;x=-78420000;
#10;x=-78410000;
#10;x=-78400000;
#10;x=-78390000;
#10;x=-78380000;
#10;x=-78370000;
#10;x=-78360000;
#10;x=-78350000;
#10;x=-78340000;
#10;x=-78330000;
#10;x=-78320000;
#10;x=-78310000;
#10;x=-78300000;
#10;x=-78290000;
#10;x=-78280000;
#10;x=-78270000;
#10;x=-78260000;
#10;x=-78250000;
#10;x=-78240000;
#10;x=-78230000;
#10;x=-78220000;
#10;x=-78210000;
#10;x=-78200000;
#10;x=-78190000;
#10;x=-78180000;
#10;x=-78170000;
#10;x=-78160000;
#10;x=-78150000;
#10;x=-78140000;
#10;x=-78130000;
#10;x=-78120000;
#10;x=-78110000;
#10;x=-78100000;
#10;x=-78090000;
#10;x=-78080000;
#10;x=-78070000;
#10;x=-78060000;
#10;x=-78050000;
#10;x=-78040000;
#10;x=-78030000;
#10;x=-78020000;
#10;x=-78010000;
#10;x=-78000000;
#10;x=-77990000;
#10;x=-77980000;
#10;x=-77970000;
#10;x=-77960000;
#10;x=-77950000;
#10;x=-77940000;
#10;x=-77930000;
#10;x=-77920000;
#10;x=-77910000;
#10;x=-77900000;
#10;x=-77890000;
#10;x=-77880000;
#10;x=-77870000;
#10;x=-77860000;
#10;x=-77850000;
#10;x=-77840000;
#10;x=-77830000;
#10;x=-77820000;
#10;x=-77810000;
#10;x=-77800000;
#10;x=-77790000;
#10;x=-77780000;
#10;x=-77770000;
#10;x=-77760000;
#10;x=-77750000;
#10;x=-77740000;
#10;x=-77730000;
#10;x=-77720000;
#10;x=-77710000;
#10;x=-77700000;
#10;x=-77690000;
#10;x=-77680000;
#10;x=-77670000;
#10;x=-77660000;
#10;x=-77650000;
#10;x=-77640000;
#10;x=-77630000;
#10;x=-77620000;
#10;x=-77610000;
#10;x=-77600000;
#10;x=-77590000;
#10;x=-77580000;
#10;x=-77570000;
#10;x=-77560000;
#10;x=-77550000;
#10;x=-77540000;
#10;x=-77530000;
#10;x=-77520000;
#10;x=-77510000;
#10;x=-77500000;
#10;x=-77490000;
#10;x=-77480000;
#10;x=-77470000;
#10;x=-77460000;
#10;x=-77450000;
#10;x=-77440000;
#10;x=-77430000;
#10;x=-77420000;
#10;x=-77410000;
#10;x=-77400000;
#10;x=-77390000;
#10;x=-77380000;
#10;x=-77370000;
#10;x=-77360000;
#10;x=-77350000;
#10;x=-77340000;
#10;x=-77330000;
#10;x=-77320000;
#10;x=-77310000;
#10;x=-77300000;
#10;x=-77290000;
#10;x=-77280000;
#10;x=-77270000;
#10;x=-77260000;
#10;x=-77250000;
#10;x=-77240000;
#10;x=-77230000;
#10;x=-77220000;
#10;x=-77210000;
#10;x=-77200000;
#10;x=-77190000;
#10;x=-77180000;
#10;x=-77170000;
#10;x=-77160000;
#10;x=-77150000;
#10;x=-77140000;
#10;x=-77130000;
#10;x=-77120000;
#10;x=-77110000;
#10;x=-77100000;
#10;x=-77090000;
#10;x=-77080000;
#10;x=-77070000;
#10;x=-77060000;
#10;x=-77050000;
#10;x=-77040000;
#10;x=-77030000;
#10;x=-77020000;
#10;x=-77010000;
#10;x=-77000000;
#10;x=-76990000;
#10;x=-76980000;
#10;x=-76970000;
#10;x=-76960000;
#10;x=-76950000;
#10;x=-76940000;
#10;x=-76930000;
#10;x=-76920000;
#10;x=-76910000;
#10;x=-76900000;
#10;x=-76890000;
#10;x=-76880000;
#10;x=-76870000;
#10;x=-76860000;
#10;x=-76850000;
#10;x=-76840000;
#10;x=-76830000;
#10;x=-76820000;
#10;x=-76810000;
#10;x=-76800000;
#10;x=-76790000;
#10;x=-76780000;
#10;x=-76770000;
#10;x=-76760000;
#10;x=-76750000;
#10;x=-76740000;
#10;x=-76730000;
#10;x=-76720000;
#10;x=-76710000;
#10;x=-76700000;
#10;x=-76690000;
#10;x=-76680000;
#10;x=-76670000;
#10;x=-76660000;
#10;x=-76650000;
#10;x=-76640000;
#10;x=-76630000;
#10;x=-76620000;
#10;x=-76610000;
#10;x=-76600000;
#10;x=-76590000;
#10;x=-76580000;
#10;x=-76570000;
#10;x=-76560000;
#10;x=-76550000;
#10;x=-76540000;
#10;x=-76530000;
#10;x=-76520000;
#10;x=-76510000;
#10;x=-76500000;
#10;x=-76490000;
#10;x=-76480000;
#10;x=-76470000;
#10;x=-76460000;
#10;x=-76450000;
#10;x=-76440000;
#10;x=-76430000;
#10;x=-76420000;
#10;x=-76410000;
#10;x=-76400000;
#10;x=-76390000;
#10;x=-76380000;
#10;x=-76370000;
#10;x=-76360000;
#10;x=-76350000;
#10;x=-76340000;
#10;x=-76330000;
#10;x=-76320000;
#10;x=-76310000;
#10;x=-76300000;
#10;x=-76290000;
#10;x=-76280000;
#10;x=-76270000;
#10;x=-76260000;
#10;x=-76250000;
#10;x=-76240000;
#10;x=-76230000;
#10;x=-76220000;
#10;x=-76210000;
#10;x=-76200000;
#10;x=-76190000;
#10;x=-76180000;
#10;x=-76170000;
#10;x=-76160000;
#10;x=-76150000;
#10;x=-76140000;
#10;x=-76130000;
#10;x=-76120000;
#10;x=-76110000;
#10;x=-76100000;
#10;x=-76090000;
#10;x=-76080000;
#10;x=-76070000;
#10;x=-76060000;
#10;x=-76050000;
#10;x=-76040000;
#10;x=-76030000;
#10;x=-76020000;
#10;x=-76010000;
#10;x=-76000000;
#10;x=-75990000;
#10;x=-75980000;
#10;x=-75970000;
#10;x=-75960000;
#10;x=-75950000;
#10;x=-75940000;
#10;x=-75930000;
#10;x=-75920000;
#10;x=-75910000;
#10;x=-75900000;
#10;x=-75890000;
#10;x=-75880000;
#10;x=-75870000;
#10;x=-75860000;
#10;x=-75850000;
#10;x=-75840000;
#10;x=-75830000;
#10;x=-75820000;
#10;x=-75810000;
#10;x=-75800000;
#10;x=-75790000;
#10;x=-75780000;
#10;x=-75770000;
#10;x=-75760000;
#10;x=-75750000;
#10;x=-75740000;
#10;x=-75730000;
#10;x=-75720000;
#10;x=-75710000;
#10;x=-75700000;
#10;x=-75690000;
#10;x=-75680000;
#10;x=-75670000;
#10;x=-75660000;
#10;x=-75650000;
#10;x=-75640000;
#10;x=-75630000;
#10;x=-75620000;
#10;x=-75610000;
#10;x=-75600000;
#10;x=-75590000;
#10;x=-75580000;
#10;x=-75570000;
#10;x=-75560000;
#10;x=-75550000;
#10;x=-75540000;
#10;x=-75530000;
#10;x=-75520000;
#10;x=-75510000;
#10;x=-75500000;
#10;x=-75490000;
#10;x=-75480000;
#10;x=-75470000;
#10;x=-75460000;
#10;x=-75450000;
#10;x=-75440000;
#10;x=-75430000;
#10;x=-75420000;
#10;x=-75410000;
#10;x=-75400000;
#10;x=-75390000;
#10;x=-75380000;
#10;x=-75370000;
#10;x=-75360000;
#10;x=-75350000;
#10;x=-75340000;
#10;x=-75330000;
#10;x=-75320000;
#10;x=-75310000;
#10;x=-75300000;
#10;x=-75290000;
#10;x=-75280000;
#10;x=-75270000;
#10;x=-75260000;
#10;x=-75250000;
#10;x=-75240000;
#10;x=-75230000;
#10;x=-75220000;
#10;x=-75210000;
#10;x=-75200000;
#10;x=-75190000;
#10;x=-75180000;
#10;x=-75170000;
#10;x=-75160000;
#10;x=-75150000;
#10;x=-75140000;
#10;x=-75130000;
#10;x=-75120000;
#10;x=-75110000;
#10;x=-75100000;
#10;x=-75090000;
#10;x=-75080000;
#10;x=-75070000;
#10;x=-75060000;
#10;x=-75050000;
#10;x=-75040000;
#10;x=-75030000;
#10;x=-75020000;
#10;x=-75010000;
#10;x=-75000000;
#10;x=-74990000;
#10;x=-74980000;
#10;x=-74970000;
#10;x=-74960000;
#10;x=-74950000;
#10;x=-74940000;
#10;x=-74930000;
#10;x=-74920000;
#10;x=-74910000;
#10;x=-74900000;
#10;x=-74890000;
#10;x=-74880000;
#10;x=-74870000;
#10;x=-74860000;
#10;x=-74850000;
#10;x=-74840000;
#10;x=-74830000;
#10;x=-74820000;
#10;x=-74810000;
#10;x=-74800000;
#10;x=-74790000;
#10;x=-74780000;
#10;x=-74770000;
#10;x=-74760000;
#10;x=-74750000;
#10;x=-74740000;
#10;x=-74730000;
#10;x=-74720000;
#10;x=-74710000;
#10;x=-74700000;
#10;x=-74690000;
#10;x=-74680000;
#10;x=-74670000;
#10;x=-74660000;
#10;x=-74650000;
#10;x=-74640000;
#10;x=-74630000;
#10;x=-74620000;
#10;x=-74610000;
#10;x=-74600000;
#10;x=-74590000;
#10;x=-74580000;
#10;x=-74570000;
#10;x=-74560000;
#10;x=-74550000;
#10;x=-74540000;
#10;x=-74530000;
#10;x=-74520000;
#10;x=-74510000;
#10;x=-74500000;
#10;x=-74490000;
#10;x=-74480000;
#10;x=-74470000;
#10;x=-74460000;
#10;x=-74450000;
#10;x=-74440000;
#10;x=-74430000;
#10;x=-74420000;
#10;x=-74410000;
#10;x=-74400000;
#10;x=-74390000;
#10;x=-74380000;
#10;x=-74370000;
#10;x=-74360000;
#10;x=-74350000;
#10;x=-74340000;
#10;x=-74330000;
#10;x=-74320000;
#10;x=-74310000;
#10;x=-74300000;
#10;x=-74290000;
#10;x=-74280000;
#10;x=-74270000;
#10;x=-74260000;
#10;x=-74250000;
#10;x=-74240000;
#10;x=-74230000;
#10;x=-74220000;
#10;x=-74210000;
#10;x=-74200000;
#10;x=-74190000;
#10;x=-74180000;
#10;x=-74170000;
#10;x=-74160000;
#10;x=-74150000;
#10;x=-74140000;
#10;x=-74130000;
#10;x=-74120000;
#10;x=-74110000;
#10;x=-74100000;
#10;x=-74090000;
#10;x=-74080000;
#10;x=-74070000;
#10;x=-74060000;
#10;x=-74050000;
#10;x=-74040000;
#10;x=-74030000;
#10;x=-74020000;
#10;x=-74010000;
#10;x=-74000000;
#10;x=-73990000;
#10;x=-73980000;
#10;x=-73970000;
#10;x=-73960000;
#10;x=-73950000;
#10;x=-73940000;
#10;x=-73930000;
#10;x=-73920000;
#10;x=-73910000;
#10;x=-73900000;
#10;x=-73890000;
#10;x=-73880000;
#10;x=-73870000;
#10;x=-73860000;
#10;x=-73850000;
#10;x=-73840000;
#10;x=-73830000;
#10;x=-73820000;
#10;x=-73810000;
#10;x=-73800000;
#10;x=-73790000;
#10;x=-73780000;
#10;x=-73770000;
#10;x=-73760000;
#10;x=-73750000;
#10;x=-73740000;
#10;x=-73730000;
#10;x=-73720000;
#10;x=-73710000;
#10;x=-73700000;
#10;x=-73690000;
#10;x=-73680000;
#10;x=-73670000;
#10;x=-73660000;
#10;x=-73650000;
#10;x=-73640000;
#10;x=-73630000;
#10;x=-73620000;
#10;x=-73610000;
#10;x=-73600000;
#10;x=-73590000;
#10;x=-73580000;
#10;x=-73570000;
#10;x=-73560000;
#10;x=-73550000;
#10;x=-73540000;
#10;x=-73530000;
#10;x=-73520000;
#10;x=-73510000;
#10;x=-73500000;
#10;x=-73490000;
#10;x=-73480000;
#10;x=-73470000;
#10;x=-73460000;
#10;x=-73450000;
#10;x=-73440000;
#10;x=-73430000;
#10;x=-73420000;
#10;x=-73410000;
#10;x=-73400000;
#10;x=-73390000;
#10;x=-73380000;
#10;x=-73370000;
#10;x=-73360000;
#10;x=-73350000;
#10;x=-73340000;
#10;x=-73330000;
#10;x=-73320000;
#10;x=-73310000;
#10;x=-73300000;
#10;x=-73290000;
#10;x=-73280000;
#10;x=-73270000;
#10;x=-73260000;
#10;x=-73250000;
#10;x=-73240000;
#10;x=-73230000;
#10;x=-73220000;
#10;x=-73210000;
#10;x=-73200000;
#10;x=-73190000;
#10;x=-73180000;
#10;x=-73170000;
#10;x=-73160000;
#10;x=-73150000;
#10;x=-73140000;
#10;x=-73130000;
#10;x=-73120000;
#10;x=-73110000;
#10;x=-73100000;
#10;x=-73090000;
#10;x=-73080000;
#10;x=-73070000;
#10;x=-73060000;
#10;x=-73050000;
#10;x=-73040000;
#10;x=-73030000;
#10;x=-73020000;
#10;x=-73010000;
#10;x=-73000000;
#10;x=-72990000;
#10;x=-72980000;
#10;x=-72970000;
#10;x=-72960000;
#10;x=-72950000;
#10;x=-72940000;
#10;x=-72930000;
#10;x=-72920000;
#10;x=-72910000;
#10;x=-72900000;
#10;x=-72890000;
#10;x=-72880000;
#10;x=-72870000;
#10;x=-72860000;
#10;x=-72850000;
#10;x=-72840000;
#10;x=-72830000;
#10;x=-72820000;
#10;x=-72810000;
#10;x=-72800000;
#10;x=-72790000;
#10;x=-72780000;
#10;x=-72770000;
#10;x=-72760000;
#10;x=-72750000;
#10;x=-72740000;
#10;x=-72730000;
#10;x=-72720000;
#10;x=-72710000;
#10;x=-72700000;
#10;x=-72690000;
#10;x=-72680000;
#10;x=-72670000;
#10;x=-72660000;
#10;x=-72650000;
#10;x=-72640000;
#10;x=-72630000;
#10;x=-72620000;
#10;x=-72610000;
#10;x=-72600000;
#10;x=-72590000;
#10;x=-72580000;
#10;x=-72570000;
#10;x=-72560000;
#10;x=-72550000;
#10;x=-72540000;
#10;x=-72530000;
#10;x=-72520000;
#10;x=-72510000;
#10;x=-72500000;
#10;x=-72490000;
#10;x=-72480000;
#10;x=-72470000;
#10;x=-72460000;
#10;x=-72450000;
#10;x=-72440000;
#10;x=-72430000;
#10;x=-72420000;
#10;x=-72410000;
#10;x=-72400000;
#10;x=-72390000;
#10;x=-72380000;
#10;x=-72370000;
#10;x=-72360000;
#10;x=-72350000;
#10;x=-72340000;
#10;x=-72330000;
#10;x=-72320000;
#10;x=-72310000;
#10;x=-72300000;
#10;x=-72290000;
#10;x=-72280000;
#10;x=-72270000;
#10;x=-72260000;
#10;x=-72250000;
#10;x=-72240000;
#10;x=-72230000;
#10;x=-72220000;
#10;x=-72210000;
#10;x=-72200000;
#10;x=-72190000;
#10;x=-72180000;
#10;x=-72170000;
#10;x=-72160000;
#10;x=-72150000;
#10;x=-72140000;
#10;x=-72130000;
#10;x=-72120000;
#10;x=-72110000;
#10;x=-72100000;
#10;x=-72090000;
#10;x=-72080000;
#10;x=-72070000;
#10;x=-72060000;
#10;x=-72050000;
#10;x=-72040000;
#10;x=-72030000;
#10;x=-72020000;
#10;x=-72010000;
#10;x=-72000000;
#10;x=-71990000;
#10;x=-71980000;
#10;x=-71970000;
#10;x=-71960000;
#10;x=-71950000;
#10;x=-71940000;
#10;x=-71930000;
#10;x=-71920000;
#10;x=-71910000;
#10;x=-71900000;
#10;x=-71890000;
#10;x=-71880000;
#10;x=-71870000;
#10;x=-71860000;
#10;x=-71850000;
#10;x=-71840000;
#10;x=-71830000;
#10;x=-71820000;
#10;x=-71810000;
#10;x=-71800000;
#10;x=-71790000;
#10;x=-71780000;
#10;x=-71770000;
#10;x=-71760000;
#10;x=-71750000;
#10;x=-71740000;
#10;x=-71730000;
#10;x=-71720000;
#10;x=-71710000;
#10;x=-71700000;
#10;x=-71690000;
#10;x=-71680000;
#10;x=-71670000;
#10;x=-71660000;
#10;x=-71650000;
#10;x=-71640000;
#10;x=-71630000;
#10;x=-71620000;
#10;x=-71610000;
#10;x=-71600000;
#10;x=-71590000;
#10;x=-71580000;
#10;x=-71570000;
#10;x=-71560000;
#10;x=-71550000;
#10;x=-71540000;
#10;x=-71530000;
#10;x=-71520000;
#10;x=-71510000;
#10;x=-71500000;
#10;x=-71490000;
#10;x=-71480000;
#10;x=-71470000;
#10;x=-71460000;
#10;x=-71450000;
#10;x=-71440000;
#10;x=-71430000;
#10;x=-71420000;
#10;x=-71410000;
#10;x=-71400000;
#10;x=-71390000;
#10;x=-71380000;
#10;x=-71370000;
#10;x=-71360000;
#10;x=-71350000;
#10;x=-71340000;
#10;x=-71330000;
#10;x=-71320000;
#10;x=-71310000;
#10;x=-71300000;
#10;x=-71290000;
#10;x=-71280000;
#10;x=-71270000;
#10;x=-71260000;
#10;x=-71250000;
#10;x=-71240000;
#10;x=-71230000;
#10;x=-71220000;
#10;x=-71210000;
#10;x=-71200000;
#10;x=-71190000;
#10;x=-71180000;
#10;x=-71170000;
#10;x=-71160000;
#10;x=-71150000;
#10;x=-71140000;
#10;x=-71130000;
#10;x=-71120000;
#10;x=-71110000;
#10;x=-71100000;
#10;x=-71090000;
#10;x=-71080000;
#10;x=-71070000;
#10;x=-71060000;
#10;x=-71050000;
#10;x=-71040000;
#10;x=-71030000;
#10;x=-71020000;
#10;x=-71010000;
#10;x=-71000000;
#10;x=-70990000;
#10;x=-70980000;
#10;x=-70970000;
#10;x=-70960000;
#10;x=-70950000;
#10;x=-70940000;
#10;x=-70930000;
#10;x=-70920000;
#10;x=-70910000;
#10;x=-70900000;
#10;x=-70890000;
#10;x=-70880000;
#10;x=-70870000;
#10;x=-70860000;
#10;x=-70850000;
#10;x=-70840000;
#10;x=-70830000;
#10;x=-70820000;
#10;x=-70810000;
#10;x=-70800000;
#10;x=-70790000;
#10;x=-70780000;
#10;x=-70770000;
#10;x=-70760000;
#10;x=-70750000;
#10;x=-70740000;
#10;x=-70730000;
#10;x=-70720000;
#10;x=-70710000;
#10;x=-70700000;
#10;x=-70690000;
#10;x=-70680000;
#10;x=-70670000;
#10;x=-70660000;
#10;x=-70650000;
#10;x=-70640000;
#10;x=-70630000;
#10;x=-70620000;
#10;x=-70610000;
#10;x=-70600000;
#10;x=-70590000;
#10;x=-70580000;
#10;x=-70570000;
#10;x=-70560000;
#10;x=-70550000;
#10;x=-70540000;
#10;x=-70530000;
#10;x=-70520000;
#10;x=-70510000;
#10;x=-70500000;
#10;x=-70490000;
#10;x=-70480000;
#10;x=-70470000;
#10;x=-70460000;
#10;x=-70450000;
#10;x=-70440000;
#10;x=-70430000;
#10;x=-70420000;
#10;x=-70410000;
#10;x=-70400000;
#10;x=-70390000;
#10;x=-70380000;
#10;x=-70370000;
#10;x=-70360000;
#10;x=-70350000;
#10;x=-70340000;
#10;x=-70330000;
#10;x=-70320000;
#10;x=-70310000;
#10;x=-70300000;
#10;x=-70290000;
#10;x=-70280000;
#10;x=-70270000;
#10;x=-70260000;
#10;x=-70250000;
#10;x=-70240000;
#10;x=-70230000;
#10;x=-70220000;
#10;x=-70210000;
#10;x=-70200000;
#10;x=-70190000;
#10;x=-70180000;
#10;x=-70170000;
#10;x=-70160000;
#10;x=-70150000;
#10;x=-70140000;
#10;x=-70130000;
#10;x=-70120000;
#10;x=-70110000;
#10;x=-70100000;
#10;x=-70090000;
#10;x=-70080000;
#10;x=-70070000;
#10;x=-70060000;
#10;x=-70050000;
#10;x=-70040000;
#10;x=-70030000;
#10;x=-70020000;
#10;x=-70010000;
#10;x=-70000000;
#10;x=-69990000;
#10;x=-69980000;
#10;x=-69970000;
#10;x=-69960000;
#10;x=-69950000;
#10;x=-69940000;
#10;x=-69930000;
#10;x=-69920000;
#10;x=-69910000;
#10;x=-69900000;
#10;x=-69890000;
#10;x=-69880000;
#10;x=-69870000;
#10;x=-69860000;
#10;x=-69850000;
#10;x=-69840000;
#10;x=-69830000;
#10;x=-69820000;
#10;x=-69810000;
#10;x=-69800000;
#10;x=-69790000;
#10;x=-69780000;
#10;x=-69770000;
#10;x=-69760000;
#10;x=-69750000;
#10;x=-69740000;
#10;x=-69730000;
#10;x=-69720000;
#10;x=-69710000;
#10;x=-69700000;
#10;x=-69690000;
#10;x=-69680000;
#10;x=-69670000;
#10;x=-69660000;
#10;x=-69650000;
#10;x=-69640000;
#10;x=-69630000;
#10;x=-69620000;
#10;x=-69610000;
#10;x=-69600000;
#10;x=-69590000;
#10;x=-69580000;
#10;x=-69570000;
#10;x=-69560000;
#10;x=-69550000;
#10;x=-69540000;
#10;x=-69530000;
#10;x=-69520000;
#10;x=-69510000;
#10;x=-69500000;
#10;x=-69490000;
#10;x=-69480000;
#10;x=-69470000;
#10;x=-69460000;
#10;x=-69450000;
#10;x=-69440000;
#10;x=-69430000;
#10;x=-69420000;
#10;x=-69410000;
#10;x=-69400000;
#10;x=-69390000;
#10;x=-69380000;
#10;x=-69370000;
#10;x=-69360000;
#10;x=-69350000;
#10;x=-69340000;
#10;x=-69330000;
#10;x=-69320000;
#10;x=-69310000;
#10;x=-69300000;
#10;x=-69290000;
#10;x=-69280000;
#10;x=-69270000;
#10;x=-69260000;
#10;x=-69250000;
#10;x=-69240000;
#10;x=-69230000;
#10;x=-69220000;
#10;x=-69210000;
#10;x=-69200000;
#10;x=-69190000;
#10;x=-69180000;
#10;x=-69170000;
#10;x=-69160000;
#10;x=-69150000;
#10;x=-69140000;
#10;x=-69130000;
#10;x=-69120000;
#10;x=-69110000;
#10;x=-69100000;
#10;x=-69090000;
#10;x=-69080000;
#10;x=-69070000;
#10;x=-69060000;
#10;x=-69050000;
#10;x=-69040000;
#10;x=-69030000;
#10;x=-69020000;
#10;x=-69010000;
#10;x=-69000000;
#10;x=-68990000;
#10;x=-68980000;
#10;x=-68970000;
#10;x=-68960000;
#10;x=-68950000;
#10;x=-68940000;
#10;x=-68930000;
#10;x=-68920000;
#10;x=-68910000;
#10;x=-68900000;
#10;x=-68890000;
#10;x=-68880000;
#10;x=-68870000;
#10;x=-68860000;
#10;x=-68850000;
#10;x=-68840000;
#10;x=-68830000;
#10;x=-68820000;
#10;x=-68810000;
#10;x=-68800000;
#10;x=-68790000;
#10;x=-68780000;
#10;x=-68770000;
#10;x=-68760000;
#10;x=-68750000;
#10;x=-68740000;
#10;x=-68730000;
#10;x=-68720000;
#10;x=-68710000;
#10;x=-68700000;
#10;x=-68690000;
#10;x=-68680000;
#10;x=-68670000;
#10;x=-68660000;
#10;x=-68650000;
#10;x=-68640000;
#10;x=-68630000;
#10;x=-68620000;
#10;x=-68610000;
#10;x=-68600000;
#10;x=-68590000;
#10;x=-68580000;
#10;x=-68570000;
#10;x=-68560000;
#10;x=-68550000;
#10;x=-68540000;
#10;x=-68530000;
#10;x=-68520000;
#10;x=-68510000;
#10;x=-68500000;
#10;x=-68490000;
#10;x=-68480000;
#10;x=-68470000;
#10;x=-68460000;
#10;x=-68450000;
#10;x=-68440000;
#10;x=-68430000;
#10;x=-68420000;
#10;x=-68410000;
#10;x=-68400000;
#10;x=-68390000;
#10;x=-68380000;
#10;x=-68370000;
#10;x=-68360000;
#10;x=-68350000;
#10;x=-68340000;
#10;x=-68330000;
#10;x=-68320000;
#10;x=-68310000;
#10;x=-68300000;
#10;x=-68290000;
#10;x=-68280000;
#10;x=-68270000;
#10;x=-68260000;
#10;x=-68250000;
#10;x=-68240000;
#10;x=-68230000;
#10;x=-68220000;
#10;x=-68210000;
#10;x=-68200000;
#10;x=-68190000;
#10;x=-68180000;
#10;x=-68170000;
#10;x=-68160000;
#10;x=-68150000;
#10;x=-68140000;
#10;x=-68130000;
#10;x=-68120000;
#10;x=-68110000;
#10;x=-68100000;
#10;x=-68090000;
#10;x=-68080000;
#10;x=-68070000;
#10;x=-68060000;
#10;x=-68050000;
#10;x=-68040000;
#10;x=-68030000;
#10;x=-68020000;
#10;x=-68010000;
#10;x=-68000000;
#10;x=-67990000;
#10;x=-67980000;
#10;x=-67970000;
#10;x=-67960000;
#10;x=-67950000;
#10;x=-67940000;
#10;x=-67930000;
#10;x=-67920000;
#10;x=-67910000;
#10;x=-67900000;
#10;x=-67890000;
#10;x=-67880000;
#10;x=-67870000;
#10;x=-67860000;
#10;x=-67850000;
#10;x=-67840000;
#10;x=-67830000;
#10;x=-67820000;
#10;x=-67810000;
#10;x=-67800000;
#10;x=-67790000;
#10;x=-67780000;
#10;x=-67770000;
#10;x=-67760000;
#10;x=-67750000;
#10;x=-67740000;
#10;x=-67730000;
#10;x=-67720000;
#10;x=-67710000;
#10;x=-67700000;
#10;x=-67690000;
#10;x=-67680000;
#10;x=-67670000;
#10;x=-67660000;
#10;x=-67650000;
#10;x=-67640000;
#10;x=-67630000;
#10;x=-67620000;
#10;x=-67610000;
#10;x=-67600000;
#10;x=-67590000;
#10;x=-67580000;
#10;x=-67570000;
#10;x=-67560000;
#10;x=-67550000;
#10;x=-67540000;
#10;x=-67530000;
#10;x=-67520000;
#10;x=-67510000;
#10;x=-67500000;
#10;x=-67490000;
#10;x=-67480000;
#10;x=-67470000;
#10;x=-67460000;
#10;x=-67450000;
#10;x=-67440000;
#10;x=-67430000;
#10;x=-67420000;
#10;x=-67410000;
#10;x=-67400000;
#10;x=-67390000;
#10;x=-67380000;
#10;x=-67370000;
#10;x=-67360000;
#10;x=-67350000;
#10;x=-67340000;
#10;x=-67330000;
#10;x=-67320000;
#10;x=-67310000;
#10;x=-67300000;
#10;x=-67290000;
#10;x=-67280000;
#10;x=-67270000;
#10;x=-67260000;
#10;x=-67250000;
#10;x=-67240000;
#10;x=-67230000;
#10;x=-67220000;
#10;x=-67210000;
#10;x=-67200000;
#10;x=-67190000;
#10;x=-67180000;
#10;x=-67170000;
#10;x=-67160000;
#10;x=-67150000;
#10;x=-67140000;
#10;x=-67130000;
#10;x=-67120000;
#10;x=-67110000;
#10;x=-67100000;
#10;x=-67090000;
#10;x=-67080000;
#10;x=-67070000;
#10;x=-67060000;
#10;x=-67050000;
#10;x=-67040000;
#10;x=-67030000;
#10;x=-67020000;
#10;x=-67010000;
#10;x=-67000000;
#10;x=-66990000;
#10;x=-66980000;
#10;x=-66970000;
#10;x=-66960000;
#10;x=-66950000;
#10;x=-66940000;
#10;x=-66930000;
#10;x=-66920000;
#10;x=-66910000;
#10;x=-66900000;
#10;x=-66890000;
#10;x=-66880000;
#10;x=-66870000;
#10;x=-66860000;
#10;x=-66850000;
#10;x=-66840000;
#10;x=-66830000;
#10;x=-66820000;
#10;x=-66810000;
#10;x=-66800000;
#10;x=-66790000;
#10;x=-66780000;
#10;x=-66770000;
#10;x=-66760000;
#10;x=-66750000;
#10;x=-66740000;
#10;x=-66730000;
#10;x=-66720000;
#10;x=-66710000;
#10;x=-66700000;
#10;x=-66690000;
#10;x=-66680000;
#10;x=-66670000;
#10;x=-66660000;
#10;x=-66650000;
#10;x=-66640000;
#10;x=-66630000;
#10;x=-66620000;
#10;x=-66610000;
#10;x=-66600000;
#10;x=-66590000;
#10;x=-66580000;
#10;x=-66570000;
#10;x=-66560000;
#10;x=-66550000;
#10;x=-66540000;
#10;x=-66530000;
#10;x=-66520000;
#10;x=-66510000;
#10;x=-66500000;
#10;x=-66490000;
#10;x=-66480000;
#10;x=-66470000;
#10;x=-66460000;
#10;x=-66450000;
#10;x=-66440000;
#10;x=-66430000;
#10;x=-66420000;
#10;x=-66410000;
#10;x=-66400000;
#10;x=-66390000;
#10;x=-66380000;
#10;x=-66370000;
#10;x=-66360000;
#10;x=-66350000;
#10;x=-66340000;
#10;x=-66330000;
#10;x=-66320000;
#10;x=-66310000;
#10;x=-66300000;
#10;x=-66290000;
#10;x=-66280000;
#10;x=-66270000;
#10;x=-66260000;
#10;x=-66250000;
#10;x=-66240000;
#10;x=-66230000;
#10;x=-66220000;
#10;x=-66210000;
#10;x=-66200000;
#10;x=-66190000;
#10;x=-66180000;
#10;x=-66170000;
#10;x=-66160000;
#10;x=-66150000;
#10;x=-66140000;
#10;x=-66130000;
#10;x=-66120000;
#10;x=-66110000;
#10;x=-66100000;
#10;x=-66090000;
#10;x=-66080000;
#10;x=-66070000;
#10;x=-66060000;
#10;x=-66050000;
#10;x=-66040000;
#10;x=-66030000;
#10;x=-66020000;
#10;x=-66010000;
#10;x=-66000000;
#10;x=-65990000;
#10;x=-65980000;
#10;x=-65970000;
#10;x=-65960000;
#10;x=-65950000;
#10;x=-65940000;
#10;x=-65930000;
#10;x=-65920000;
#10;x=-65910000;
#10;x=-65900000;
#10;x=-65890000;
#10;x=-65880000;
#10;x=-65870000;
#10;x=-65860000;
#10;x=-65850000;
#10;x=-65840000;
#10;x=-65830000;
#10;x=-65820000;
#10;x=-65810000;
#10;x=-65800000;
#10;x=-65790000;
#10;x=-65780000;
#10;x=-65770000;
#10;x=-65760000;
#10;x=-65750000;
#10;x=-65740000;
#10;x=-65730000;
#10;x=-65720000;
#10;x=-65710000;
#10;x=-65700000;
#10;x=-65690000;
#10;x=-65680000;
#10;x=-65670000;
#10;x=-65660000;
#10;x=-65650000;
#10;x=-65640000;
#10;x=-65630000;
#10;x=-65620000;
#10;x=-65610000;
#10;x=-65600000;
#10;x=-65590000;
#10;x=-65580000;
#10;x=-65570000;
#10;x=-65560000;
#10;x=-65550000;
#10;x=-65540000;
#10;x=-65530000;
#10;x=-65520000;
#10;x=-65510000;
#10;x=-65500000;
#10;x=-65490000;
#10;x=-65480000;
#10;x=-65470000;
#10;x=-65460000;
#10;x=-65450000;
#10;x=-65440000;
#10;x=-65430000;
#10;x=-65420000;
#10;x=-65410000;
#10;x=-65400000;
#10;x=-65390000;
#10;x=-65380000;
#10;x=-65370000;
#10;x=-65360000;
#10;x=-65350000;
#10;x=-65340000;
#10;x=-65330000;
#10;x=-65320000;
#10;x=-65310000;
#10;x=-65300000;
#10;x=-65290000;
#10;x=-65280000;
#10;x=-65270000;
#10;x=-65260000;
#10;x=-65250000;
#10;x=-65240000;
#10;x=-65230000;
#10;x=-65220000;
#10;x=-65210000;
#10;x=-65200000;
#10;x=-65190000;
#10;x=-65180000;
#10;x=-65170000;
#10;x=-65160000;
#10;x=-65150000;
#10;x=-65140000;
#10;x=-65130000;
#10;x=-65120000;
#10;x=-65110000;
#10;x=-65100000;
#10;x=-65090000;
#10;x=-65080000;
#10;x=-65070000;
#10;x=-65060000;
#10;x=-65050000;
#10;x=-65040000;
#10;x=-65030000;
#10;x=-65020000;
#10;x=-65010000;
#10;x=-65000000;
#10;x=-64990000;
#10;x=-64980000;
#10;x=-64970000;
#10;x=-64960000;
#10;x=-64950000;
#10;x=-64940000;
#10;x=-64930000;
#10;x=-64920000;
#10;x=-64910000;
#10;x=-64900000;
#10;x=-64890000;
#10;x=-64880000;
#10;x=-64870000;
#10;x=-64860000;
#10;x=-64850000;
#10;x=-64840000;
#10;x=-64830000;
#10;x=-64820000;
#10;x=-64810000;
#10;x=-64800000;
#10;x=-64790000;
#10;x=-64780000;
#10;x=-64770000;
#10;x=-64760000;
#10;x=-64750000;
#10;x=-64740000;
#10;x=-64730000;
#10;x=-64720000;
#10;x=-64710000;
#10;x=-64700000;
#10;x=-64690000;
#10;x=-64680000;
#10;x=-64670000;
#10;x=-64660000;
#10;x=-64650000;
#10;x=-64640000;
#10;x=-64630000;
#10;x=-64620000;
#10;x=-64610000;
#10;x=-64600000;
#10;x=-64590000;
#10;x=-64580000;
#10;x=-64570000;
#10;x=-64560000;
#10;x=-64550000;
#10;x=-64540000;
#10;x=-64530000;
#10;x=-64520000;
#10;x=-64510000;
#10;x=-64500000;
#10;x=-64490000;
#10;x=-64480000;
#10;x=-64470000;
#10;x=-64460000;
#10;x=-64450000;
#10;x=-64440000;
#10;x=-64430000;
#10;x=-64420000;
#10;x=-64410000;
#10;x=-64400000;
#10;x=-64390000;
#10;x=-64380000;
#10;x=-64370000;
#10;x=-64360000;
#10;x=-64350000;
#10;x=-64340000;
#10;x=-64330000;
#10;x=-64320000;
#10;x=-64310000;
#10;x=-64300000;
#10;x=-64290000;
#10;x=-64280000;
#10;x=-64270000;
#10;x=-64260000;
#10;x=-64250000;
#10;x=-64240000;
#10;x=-64230000;
#10;x=-64220000;
#10;x=-64210000;
#10;x=-64200000;
#10;x=-64190000;
#10;x=-64180000;
#10;x=-64170000;
#10;x=-64160000;
#10;x=-64150000;
#10;x=-64140000;
#10;x=-64130000;
#10;x=-64120000;
#10;x=-64110000;
#10;x=-64100000;
#10;x=-64090000;
#10;x=-64080000;
#10;x=-64070000;
#10;x=-64060000;
#10;x=-64050000;
#10;x=-64040000;
#10;x=-64030000;
#10;x=-64020000;
#10;x=-64010000;
#10;x=-64000000;
#10;x=-63990000;
#10;x=-63980000;
#10;x=-63970000;
#10;x=-63960000;
#10;x=-63950000;
#10;x=-63940000;
#10;x=-63930000;
#10;x=-63920000;
#10;x=-63910000;
#10;x=-63900000;
#10;x=-63890000;
#10;x=-63880000;
#10;x=-63870000;
#10;x=-63860000;
#10;x=-63850000;
#10;x=-63840000;
#10;x=-63830000;
#10;x=-63820000;
#10;x=-63810000;
#10;x=-63800000;
#10;x=-63790000;
#10;x=-63780000;
#10;x=-63770000;
#10;x=-63760000;
#10;x=-63750000;
#10;x=-63740000;
#10;x=-63730000;
#10;x=-63720000;
#10;x=-63710000;
#10;x=-63700000;
#10;x=-63690000;
#10;x=-63680000;
#10;x=-63670000;
#10;x=-63660000;
#10;x=-63650000;
#10;x=-63640000;
#10;x=-63630000;
#10;x=-63620000;
#10;x=-63610000;
#10;x=-63600000;
#10;x=-63590000;
#10;x=-63580000;
#10;x=-63570000;
#10;x=-63560000;
#10;x=-63550000;
#10;x=-63540000;
#10;x=-63530000;
#10;x=-63520000;
#10;x=-63510000;
#10;x=-63500000;
#10;x=-63490000;
#10;x=-63480000;
#10;x=-63470000;
#10;x=-63460000;
#10;x=-63450000;
#10;x=-63440000;
#10;x=-63430000;
#10;x=-63420000;
#10;x=-63410000;
#10;x=-63400000;
#10;x=-63390000;
#10;x=-63380000;
#10;x=-63370000;
#10;x=-63360000;
#10;x=-63350000;
#10;x=-63340000;
#10;x=-63330000;
#10;x=-63320000;
#10;x=-63310000;
#10;x=-63300000;
#10;x=-63290000;
#10;x=-63280000;
#10;x=-63270000;
#10;x=-63260000;
#10;x=-63250000;
#10;x=-63240000;
#10;x=-63230000;
#10;x=-63220000;
#10;x=-63210000;
#10;x=-63200000;
#10;x=-63190000;
#10;x=-63180000;
#10;x=-63170000;
#10;x=-63160000;
#10;x=-63150000;
#10;x=-63140000;
#10;x=-63130000;
#10;x=-63120000;
#10;x=-63110000;
#10;x=-63100000;
#10;x=-63090000;
#10;x=-63080000;
#10;x=-63070000;
#10;x=-63060000;
#10;x=-63050000;
#10;x=-63040000;
#10;x=-63030000;
#10;x=-63020000;
#10;x=-63010000;
#10;x=-63000000;
#10;x=-62990000;
#10;x=-62980000;
#10;x=-62970000;
#10;x=-62960000;
#10;x=-62950000;
#10;x=-62940000;
#10;x=-62930000;
#10;x=-62920000;
#10;x=-62910000;
#10;x=-62900000;
#10;x=-62890000;
#10;x=-62880000;
#10;x=-62870000;
#10;x=-62860000;
#10;x=-62850000;
#10;x=-62840000;
#10;x=-62830000;
#10;x=-62820000;
#10;x=-62810000;
#10;x=-62800000;
#10;x=-62790000;
#10;x=-62780000;
#10;x=-62770000;
#10;x=-62760000;
#10;x=-62750000;
#10;x=-62740000;
#10;x=-62730000;
#10;x=-62720000;
#10;x=-62710000;
#10;x=-62700000;
#10;x=-62690000;
#10;x=-62680000;
#10;x=-62670000;
#10;x=-62660000;
#10;x=-62650000;
#10;x=-62640000;
#10;x=-62630000;
#10;x=-62620000;
#10;x=-62610000;
#10;x=-62600000;
#10;x=-62590000;
#10;x=-62580000;
#10;x=-62570000;
#10;x=-62560000;
#10;x=-62550000;
#10;x=-62540000;
#10;x=-62530000;
#10;x=-62520000;
#10;x=-62510000;
#10;x=-62500000;
#10;x=-62490000;
#10;x=-62480000;
#10;x=-62470000;
#10;x=-62460000;
#10;x=-62450000;
#10;x=-62440000;
#10;x=-62430000;
#10;x=-62420000;
#10;x=-62410000;
#10;x=-62400000;
#10;x=-62390000;
#10;x=-62380000;
#10;x=-62370000;
#10;x=-62360000;
#10;x=-62350000;
#10;x=-62340000;
#10;x=-62330000;
#10;x=-62320000;
#10;x=-62310000;
#10;x=-62300000;
#10;x=-62290000;
#10;x=-62280000;
#10;x=-62270000;
#10;x=-62260000;
#10;x=-62250000;
#10;x=-62240000;
#10;x=-62230000;
#10;x=-62220000;
#10;x=-62210000;
#10;x=-62200000;
#10;x=-62190000;
#10;x=-62180000;
#10;x=-62170000;
#10;x=-62160000;
#10;x=-62150000;
#10;x=-62140000;
#10;x=-62130000;
#10;x=-62120000;
#10;x=-62110000;
#10;x=-62100000;
#10;x=-62090000;
#10;x=-62080000;
#10;x=-62070000;
#10;x=-62060000;
#10;x=-62050000;
#10;x=-62040000;
#10;x=-62030000;
#10;x=-62020000;
#10;x=-62010000;
#10;x=-62000000;
#10;x=-61990000;
#10;x=-61980000;
#10;x=-61970000;
#10;x=-61960000;
#10;x=-61950000;
#10;x=-61940000;
#10;x=-61930000;
#10;x=-61920000;
#10;x=-61910000;
#10;x=-61900000;
#10;x=-61890000;
#10;x=-61880000;
#10;x=-61870000;
#10;x=-61860000;
#10;x=-61850000;
#10;x=-61840000;
#10;x=-61830000;
#10;x=-61820000;
#10;x=-61810000;
#10;x=-61800000;
#10;x=-61790000;
#10;x=-61780000;
#10;x=-61770000;
#10;x=-61760000;
#10;x=-61750000;
#10;x=-61740000;
#10;x=-61730000;
#10;x=-61720000;
#10;x=-61710000;
#10;x=-61700000;
#10;x=-61690000;
#10;x=-61680000;
#10;x=-61670000;
#10;x=-61660000;
#10;x=-61650000;
#10;x=-61640000;
#10;x=-61630000;
#10;x=-61620000;
#10;x=-61610000;
#10;x=-61600000;
#10;x=-61590000;
#10;x=-61580000;
#10;x=-61570000;
#10;x=-61560000;
#10;x=-61550000;
#10;x=-61540000;
#10;x=-61530000;
#10;x=-61520000;
#10;x=-61510000;
#10;x=-61500000;
#10;x=-61490000;
#10;x=-61480000;
#10;x=-61470000;
#10;x=-61460000;
#10;x=-61450000;
#10;x=-61440000;
#10;x=-61430000;
#10;x=-61420000;
#10;x=-61410000;
#10;x=-61400000;
#10;x=-61390000;
#10;x=-61380000;
#10;x=-61370000;
#10;x=-61360000;
#10;x=-61350000;
#10;x=-61340000;
#10;x=-61330000;
#10;x=-61320000;
#10;x=-61310000;
#10;x=-61300000;
#10;x=-61290000;
#10;x=-61280000;
#10;x=-61270000;
#10;x=-61260000;
#10;x=-61250000;
#10;x=-61240000;
#10;x=-61230000;
#10;x=-61220000;
#10;x=-61210000;
#10;x=-61200000;
#10;x=-61190000;
#10;x=-61180000;
#10;x=-61170000;
#10;x=-61160000;
#10;x=-61150000;
#10;x=-61140000;
#10;x=-61130000;
#10;x=-61120000;
#10;x=-61110000;
#10;x=-61100000;
#10;x=-61090000;
#10;x=-61080000;
#10;x=-61070000;
#10;x=-61060000;
#10;x=-61050000;
#10;x=-61040000;
#10;x=-61030000;
#10;x=-61020000;
#10;x=-61010000;
#10;x=-61000000;
#10;x=-60990000;
#10;x=-60980000;
#10;x=-60970000;
#10;x=-60960000;
#10;x=-60950000;
#10;x=-60940000;
#10;x=-60930000;
#10;x=-60920000;
#10;x=-60910000;
#10;x=-60900000;
#10;x=-60890000;
#10;x=-60880000;
#10;x=-60870000;
#10;x=-60860000;
#10;x=-60850000;
#10;x=-60840000;
#10;x=-60830000;
#10;x=-60820000;
#10;x=-60810000;
#10;x=-60800000;
#10;x=-60790000;
#10;x=-60780000;
#10;x=-60770000;
#10;x=-60760000;
#10;x=-60750000;
#10;x=-60740000;
#10;x=-60730000;
#10;x=-60720000;
#10;x=-60710000;
#10;x=-60700000;
#10;x=-60690000;
#10;x=-60680000;
#10;x=-60670000;
#10;x=-60660000;
#10;x=-60650000;
#10;x=-60640000;
#10;x=-60630000;
#10;x=-60620000;
#10;x=-60610000;
#10;x=-60600000;
#10;x=-60590000;
#10;x=-60580000;
#10;x=-60570000;
#10;x=-60560000;
#10;x=-60550000;
#10;x=-60540000;
#10;x=-60530000;
#10;x=-60520000;
#10;x=-60510000;
#10;x=-60500000;
#10;x=-60490000;
#10;x=-60480000;
#10;x=-60470000;
#10;x=-60460000;
#10;x=-60450000;
#10;x=-60440000;
#10;x=-60430000;
#10;x=-60420000;
#10;x=-60410000;
#10;x=-60400000;
#10;x=-60390000;
#10;x=-60380000;
#10;x=-60370000;
#10;x=-60360000;
#10;x=-60350000;
#10;x=-60340000;
#10;x=-60330000;
#10;x=-60320000;
#10;x=-60310000;
#10;x=-60300000;
#10;x=-60290000;
#10;x=-60280000;
#10;x=-60270000;
#10;x=-60260000;
#10;x=-60250000;
#10;x=-60240000;
#10;x=-60230000;
#10;x=-60220000;
#10;x=-60210000;
#10;x=-60200000;
#10;x=-60190000;
#10;x=-60180000;
#10;x=-60170000;
#10;x=-60160000;
#10;x=-60150000;
#10;x=-60140000;
#10;x=-60130000;
#10;x=-60120000;
#10;x=-60110000;
#10;x=-60100000;
#10;x=-60090000;
#10;x=-60080000;
#10;x=-60070000;
#10;x=-60060000;
#10;x=-60050000;
#10;x=-60040000;
#10;x=-60030000;
#10;x=-60020000;
#10;x=-60010000;
#10;x=-60000000;
#10;x=-59990000;
#10;x=-59980000;
#10;x=-59970000;
#10;x=-59960000;
#10;x=-59950000;
#10;x=-59940000;
#10;x=-59930000;
#10;x=-59920000;
#10;x=-59910000;
#10;x=-59900000;
#10;x=-59890000;
#10;x=-59880000;
#10;x=-59870000;
#10;x=-59860000;
#10;x=-59850000;
#10;x=-59840000;
#10;x=-59830000;
#10;x=-59820000;
#10;x=-59810000;
#10;x=-59800000;
#10;x=-59790000;
#10;x=-59780000;
#10;x=-59770000;
#10;x=-59760000;
#10;x=-59750000;
#10;x=-59740000;
#10;x=-59730000;
#10;x=-59720000;
#10;x=-59710000;
#10;x=-59700000;
#10;x=-59690000;
#10;x=-59680000;
#10;x=-59670000;
#10;x=-59660000;
#10;x=-59650000;
#10;x=-59640000;
#10;x=-59630000;
#10;x=-59620000;
#10;x=-59610000;
#10;x=-59600000;
#10;x=-59590000;
#10;x=-59580000;
#10;x=-59570000;
#10;x=-59560000;
#10;x=-59550000;
#10;x=-59540000;
#10;x=-59530000;
#10;x=-59520000;
#10;x=-59510000;
#10;x=-59500000;
#10;x=-59490000;
#10;x=-59480000;
#10;x=-59470000;
#10;x=-59460000;
#10;x=-59450000;
#10;x=-59440000;
#10;x=-59430000;
#10;x=-59420000;
#10;x=-59410000;
#10;x=-59400000;
#10;x=-59390000;
#10;x=-59380000;
#10;x=-59370000;
#10;x=-59360000;
#10;x=-59350000;
#10;x=-59340000;
#10;x=-59330000;
#10;x=-59320000;
#10;x=-59310000;
#10;x=-59300000;
#10;x=-59290000;
#10;x=-59280000;
#10;x=-59270000;
#10;x=-59260000;
#10;x=-59250000;
#10;x=-59240000;
#10;x=-59230000;
#10;x=-59220000;
#10;x=-59210000;
#10;x=-59200000;
#10;x=-59190000;
#10;x=-59180000;
#10;x=-59170000;
#10;x=-59160000;
#10;x=-59150000;
#10;x=-59140000;
#10;x=-59130000;
#10;x=-59120000;
#10;x=-59110000;
#10;x=-59100000;
#10;x=-59090000;
#10;x=-59080000;
#10;x=-59070000;
#10;x=-59060000;
#10;x=-59050000;
#10;x=-59040000;
#10;x=-59030000;
#10;x=-59020000;
#10;x=-59010000;
#10;x=-59000000;
#10;x=-58990000;
#10;x=-58980000;
#10;x=-58970000;
#10;x=-58960000;
#10;x=-58950000;
#10;x=-58940000;
#10;x=-58930000;
#10;x=-58920000;
#10;x=-58910000;
#10;x=-58900000;
#10;x=-58890000;
#10;x=-58880000;
#10;x=-58870000;
#10;x=-58860000;
#10;x=-58850000;
#10;x=-58840000;
#10;x=-58830000;
#10;x=-58820000;
#10;x=-58810000;
#10;x=-58800000;
#10;x=-58790000;
#10;x=-58780000;
#10;x=-58770000;
#10;x=-58760000;
#10;x=-58750000;
#10;x=-58740000;
#10;x=-58730000;
#10;x=-58720000;
#10;x=-58710000;
#10;x=-58700000;
#10;x=-58690000;
#10;x=-58680000;
#10;x=-58670000;
#10;x=-58660000;
#10;x=-58650000;
#10;x=-58640000;
#10;x=-58630000;
#10;x=-58620000;
#10;x=-58610000;
#10;x=-58600000;
#10;x=-58590000;
#10;x=-58580000;
#10;x=-58570000;
#10;x=-58560000;
#10;x=-58550000;
#10;x=-58540000;
#10;x=-58530000;
#10;x=-58520000;
#10;x=-58510000;
#10;x=-58500000;
#10;x=-58490000;
#10;x=-58480000;
#10;x=-58470000;
#10;x=-58460000;
#10;x=-58450000;
#10;x=-58440000;
#10;x=-58430000;
#10;x=-58420000;
#10;x=-58410000;
#10;x=-58400000;
#10;x=-58390000;
#10;x=-58380000;
#10;x=-58370000;
#10;x=-58360000;
#10;x=-58350000;
#10;x=-58340000;
#10;x=-58330000;
#10;x=-58320000;
#10;x=-58310000;
#10;x=-58300000;
#10;x=-58290000;
#10;x=-58280000;
#10;x=-58270000;
#10;x=-58260000;
#10;x=-58250000;
#10;x=-58240000;
#10;x=-58230000;
#10;x=-58220000;
#10;x=-58210000;
#10;x=-58200000;
#10;x=-58190000;
#10;x=-58180000;
#10;x=-58170000;
#10;x=-58160000;
#10;x=-58150000;
#10;x=-58140000;
#10;x=-58130000;
#10;x=-58120000;
#10;x=-58110000;
#10;x=-58100000;
#10;x=-58090000;
#10;x=-58080000;
#10;x=-58070000;
#10;x=-58060000;
#10;x=-58050000;
#10;x=-58040000;
#10;x=-58030000;
#10;x=-58020000;
#10;x=-58010000;
#10;x=-58000000;
#10;x=-57990000;
#10;x=-57980000;
#10;x=-57970000;
#10;x=-57960000;
#10;x=-57950000;
#10;x=-57940000;
#10;x=-57930000;
#10;x=-57920000;
#10;x=-57910000;
#10;x=-57900000;
#10;x=-57890000;
#10;x=-57880000;
#10;x=-57870000;
#10;x=-57860000;
#10;x=-57850000;
#10;x=-57840000;
#10;x=-57830000;
#10;x=-57820000;
#10;x=-57810000;
#10;x=-57800000;
#10;x=-57790000;
#10;x=-57780000;
#10;x=-57770000;
#10;x=-57760000;
#10;x=-57750000;
#10;x=-57740000;
#10;x=-57730000;
#10;x=-57720000;
#10;x=-57710000;
#10;x=-57700000;
#10;x=-57690000;
#10;x=-57680000;
#10;x=-57670000;
#10;x=-57660000;
#10;x=-57650000;
#10;x=-57640000;
#10;x=-57630000;
#10;x=-57620000;
#10;x=-57610000;
#10;x=-57600000;
#10;x=-57590000;
#10;x=-57580000;
#10;x=-57570000;
#10;x=-57560000;
#10;x=-57550000;
#10;x=-57540000;
#10;x=-57530000;
#10;x=-57520000;
#10;x=-57510000;
#10;x=-57500000;
#10;x=-57490000;
#10;x=-57480000;
#10;x=-57470000;
#10;x=-57460000;
#10;x=-57450000;
#10;x=-57440000;
#10;x=-57430000;
#10;x=-57420000;
#10;x=-57410000;
#10;x=-57400000;
#10;x=-57390000;
#10;x=-57380000;
#10;x=-57370000;
#10;x=-57360000;
#10;x=-57350000;
#10;x=-57340000;
#10;x=-57330000;
#10;x=-57320000;
#10;x=-57310000;
#10;x=-57300000;
#10;x=-57290000;
#10;x=-57280000;
#10;x=-57270000;
#10;x=-57260000;
#10;x=-57250000;
#10;x=-57240000;
#10;x=-57230000;
#10;x=-57220000;
#10;x=-57210000;
#10;x=-57200000;
#10;x=-57190000;
#10;x=-57180000;
#10;x=-57170000;
#10;x=-57160000;
#10;x=-57150000;
#10;x=-57140000;
#10;x=-57130000;
#10;x=-57120000;
#10;x=-57110000;
#10;x=-57100000;
#10;x=-57090000;
#10;x=-57080000;
#10;x=-57070000;
#10;x=-57060000;
#10;x=-57050000;
#10;x=-57040000;
#10;x=-57030000;
#10;x=-57020000;
#10;x=-57010000;
#10;x=-57000000;
#10;x=-56990000;
#10;x=-56980000;
#10;x=-56970000;
#10;x=-56960000;
#10;x=-56950000;
#10;x=-56940000;
#10;x=-56930000;
#10;x=-56920000;
#10;x=-56910000;
#10;x=-56900000;
#10;x=-56890000;
#10;x=-56880000;
#10;x=-56870000;
#10;x=-56860000;
#10;x=-56850000;
#10;x=-56840000;
#10;x=-56830000;
#10;x=-56820000;
#10;x=-56810000;
#10;x=-56800000;
#10;x=-56790000;
#10;x=-56780000;
#10;x=-56770000;
#10;x=-56760000;
#10;x=-56750000;
#10;x=-56740000;
#10;x=-56730000;
#10;x=-56720000;
#10;x=-56710000;
#10;x=-56700000;
#10;x=-56690000;
#10;x=-56680000;
#10;x=-56670000;
#10;x=-56660000;
#10;x=-56650000;
#10;x=-56640000;
#10;x=-56630000;
#10;x=-56620000;
#10;x=-56610000;
#10;x=-56600000;
#10;x=-56590000;
#10;x=-56580000;
#10;x=-56570000;
#10;x=-56560000;
#10;x=-56550000;
#10;x=-56540000;
#10;x=-56530000;
#10;x=-56520000;
#10;x=-56510000;
#10;x=-56500000;
#10;x=-56490000;
#10;x=-56480000;
#10;x=-56470000;
#10;x=-56460000;
#10;x=-56450000;
#10;x=-56440000;
#10;x=-56430000;
#10;x=-56420000;
#10;x=-56410000;
#10;x=-56400000;
#10;x=-56390000;
#10;x=-56380000;
#10;x=-56370000;
#10;x=-56360000;
#10;x=-56350000;
#10;x=-56340000;
#10;x=-56330000;
#10;x=-56320000;
#10;x=-56310000;
#10;x=-56300000;
#10;x=-56290000;
#10;x=-56280000;
#10;x=-56270000;
#10;x=-56260000;
#10;x=-56250000;
#10;x=-56240000;
#10;x=-56230000;
#10;x=-56220000;
#10;x=-56210000;
#10;x=-56200000;
#10;x=-56190000;
#10;x=-56180000;
#10;x=-56170000;
#10;x=-56160000;
#10;x=-56150000;
#10;x=-56140000;
#10;x=-56130000;
#10;x=-56120000;
#10;x=-56110000;
#10;x=-56100000;
#10;x=-56090000;
#10;x=-56080000;
#10;x=-56070000;
#10;x=-56060000;
#10;x=-56050000;
#10;x=-56040000;
#10;x=-56030000;
#10;x=-56020000;
#10;x=-56010000;
#10;x=-56000000;
#10;x=-55990000;
#10;x=-55980000;
#10;x=-55970000;
#10;x=-55960000;
#10;x=-55950000;
#10;x=-55940000;
#10;x=-55930000;
#10;x=-55920000;
#10;x=-55910000;
#10;x=-55900000;
#10;x=-55890000;
#10;x=-55880000;
#10;x=-55870000;
#10;x=-55860000;
#10;x=-55850000;
#10;x=-55840000;
#10;x=-55830000;
#10;x=-55820000;
#10;x=-55810000;
#10;x=-55800000;
#10;x=-55790000;
#10;x=-55780000;
#10;x=-55770000;
#10;x=-55760000;
#10;x=-55750000;
#10;x=-55740000;
#10;x=-55730000;
#10;x=-55720000;
#10;x=-55710000;
#10;x=-55700000;
#10;x=-55690000;
#10;x=-55680000;
#10;x=-55670000;
#10;x=-55660000;
#10;x=-55650000;
#10;x=-55640000;
#10;x=-55630000;
#10;x=-55620000;
#10;x=-55610000;
#10;x=-55600000;
#10;x=-55590000;
#10;x=-55580000;
#10;x=-55570000;
#10;x=-55560000;
#10;x=-55550000;
#10;x=-55540000;
#10;x=-55530000;
#10;x=-55520000;
#10;x=-55510000;
#10;x=-55500000;
#10;x=-55490000;
#10;x=-55480000;
#10;x=-55470000;
#10;x=-55460000;
#10;x=-55450000;
#10;x=-55440000;
#10;x=-55430000;
#10;x=-55420000;
#10;x=-55410000;
#10;x=-55400000;
#10;x=-55390000;
#10;x=-55380000;
#10;x=-55370000;
#10;x=-55360000;
#10;x=-55350000;
#10;x=-55340000;
#10;x=-55330000;
#10;x=-55320000;
#10;x=-55310000;
#10;x=-55300000;
#10;x=-55290000;
#10;x=-55280000;
#10;x=-55270000;
#10;x=-55260000;
#10;x=-55250000;
#10;x=-55240000;
#10;x=-55230000;
#10;x=-55220000;
#10;x=-55210000;
#10;x=-55200000;
#10;x=-55190000;
#10;x=-55180000;
#10;x=-55170000;
#10;x=-55160000;
#10;x=-55150000;
#10;x=-55140000;
#10;x=-55130000;
#10;x=-55120000;
#10;x=-55110000;
#10;x=-55100000;
#10;x=-55090000;
#10;x=-55080000;
#10;x=-55070000;
#10;x=-55060000;
#10;x=-55050000;
#10;x=-55040000;
#10;x=-55030000;
#10;x=-55020000;
#10;x=-55010000;
#10;x=-55000000;
#10;x=-54990000;
#10;x=-54980000;
#10;x=-54970000;
#10;x=-54960000;
#10;x=-54950000;
#10;x=-54940000;
#10;x=-54930000;
#10;x=-54920000;
#10;x=-54910000;
#10;x=-54900000;
#10;x=-54890000;
#10;x=-54880000;
#10;x=-54870000;
#10;x=-54860000;
#10;x=-54850000;
#10;x=-54840000;
#10;x=-54830000;
#10;x=-54820000;
#10;x=-54810000;
#10;x=-54800000;
#10;x=-54790000;
#10;x=-54780000;
#10;x=-54770000;
#10;x=-54760000;
#10;x=-54750000;
#10;x=-54740000;
#10;x=-54730000;
#10;x=-54720000;
#10;x=-54710000;
#10;x=-54700000;
#10;x=-54690000;
#10;x=-54680000;
#10;x=-54670000;
#10;x=-54660000;
#10;x=-54650000;
#10;x=-54640000;
#10;x=-54630000;
#10;x=-54620000;
#10;x=-54610000;
#10;x=-54600000;
#10;x=-54590000;
#10;x=-54580000;
#10;x=-54570000;
#10;x=-54560000;
#10;x=-54550000;
#10;x=-54540000;
#10;x=-54530000;
#10;x=-54520000;
#10;x=-54510000;
#10;x=-54500000;
#10;x=-54490000;
#10;x=-54480000;
#10;x=-54470000;
#10;x=-54460000;
#10;x=-54450000;
#10;x=-54440000;
#10;x=-54430000;
#10;x=-54420000;
#10;x=-54410000;
#10;x=-54400000;
#10;x=-54390000;
#10;x=-54380000;
#10;x=-54370000;
#10;x=-54360000;
#10;x=-54350000;
#10;x=-54340000;
#10;x=-54330000;
#10;x=-54320000;
#10;x=-54310000;
#10;x=-54300000;
#10;x=-54290000;
#10;x=-54280000;
#10;x=-54270000;
#10;x=-54260000;
#10;x=-54250000;
#10;x=-54240000;
#10;x=-54230000;
#10;x=-54220000;
#10;x=-54210000;
#10;x=-54200000;
#10;x=-54190000;
#10;x=-54180000;
#10;x=-54170000;
#10;x=-54160000;
#10;x=-54150000;
#10;x=-54140000;
#10;x=-54130000;
#10;x=-54120000;
#10;x=-54110000;
#10;x=-54100000;
#10;x=-54090000;
#10;x=-54080000;
#10;x=-54070000;
#10;x=-54060000;
#10;x=-54050000;
#10;x=-54040000;
#10;x=-54030000;
#10;x=-54020000;
#10;x=-54010000;
#10;x=-54000000;
#10;x=-53990000;
#10;x=-53980000;
#10;x=-53970000;
#10;x=-53960000;
#10;x=-53950000;
#10;x=-53940000;
#10;x=-53930000;
#10;x=-53920000;
#10;x=-53910000;
#10;x=-53900000;
#10;x=-53890000;
#10;x=-53880000;
#10;x=-53870000;
#10;x=-53860000;
#10;x=-53850000;
#10;x=-53840000;
#10;x=-53830000;
#10;x=-53820000;
#10;x=-53810000;
#10;x=-53800000;
#10;x=-53790000;
#10;x=-53780000;
#10;x=-53770000;
#10;x=-53760000;
#10;x=-53750000;
#10;x=-53740000;
#10;x=-53730000;
#10;x=-53720000;
#10;x=-53710000;
#10;x=-53700000;
#10;x=-53690000;
#10;x=-53680000;
#10;x=-53670000;
#10;x=-53660000;
#10;x=-53650000;
#10;x=-53640000;
#10;x=-53630000;
#10;x=-53620000;
#10;x=-53610000;
#10;x=-53600000;
#10;x=-53590000;
#10;x=-53580000;
#10;x=-53570000;
#10;x=-53560000;
#10;x=-53550000;
#10;x=-53540000;
#10;x=-53530000;
#10;x=-53520000;
#10;x=-53510000;
#10;x=-53500000;
#10;x=-53490000;
#10;x=-53480000;
#10;x=-53470000;
#10;x=-53460000;
#10;x=-53450000;
#10;x=-53440000;
#10;x=-53430000;
#10;x=-53420000;
#10;x=-53410000;
#10;x=-53400000;
#10;x=-53390000;
#10;x=-53380000;
#10;x=-53370000;
#10;x=-53360000;
#10;x=-53350000;
#10;x=-53340000;
#10;x=-53330000;
#10;x=-53320000;
#10;x=-53310000;
#10;x=-53300000;
#10;x=-53290000;
#10;x=-53280000;
#10;x=-53270000;
#10;x=-53260000;
#10;x=-53250000;
#10;x=-53240000;
#10;x=-53230000;
#10;x=-53220000;
#10;x=-53210000;
#10;x=-53200000;
#10;x=-53190000;
#10;x=-53180000;
#10;x=-53170000;
#10;x=-53160000;
#10;x=-53150000;
#10;x=-53140000;
#10;x=-53130000;
#10;x=-53120000;
#10;x=-53110000;
#10;x=-53100000;
#10;x=-53090000;
#10;x=-53080000;
#10;x=-53070000;
#10;x=-53060000;
#10;x=-53050000;
#10;x=-53040000;
#10;x=-53030000;
#10;x=-53020000;
#10;x=-53010000;
#10;x=-53000000;
#10;x=-52990000;
#10;x=-52980000;
#10;x=-52970000;
#10;x=-52960000;
#10;x=-52950000;
#10;x=-52940000;
#10;x=-52930000;
#10;x=-52920000;
#10;x=-52910000;
#10;x=-52900000;
#10;x=-52890000;
#10;x=-52880000;
#10;x=-52870000;
#10;x=-52860000;
#10;x=-52850000;
#10;x=-52840000;
#10;x=-52830000;
#10;x=-52820000;
#10;x=-52810000;
#10;x=-52800000;
#10;x=-52790000;
#10;x=-52780000;
#10;x=-52770000;
#10;x=-52760000;
#10;x=-52750000;
#10;x=-52740000;
#10;x=-52730000;
#10;x=-52720000;
#10;x=-52710000;
#10;x=-52700000;
#10;x=-52690000;
#10;x=-52680000;
#10;x=-52670000;
#10;x=-52660000;
#10;x=-52650000;
#10;x=-52640000;
#10;x=-52630000;
#10;x=-52620000;
#10;x=-52610000;
#10;x=-52600000;
#10;x=-52590000;
#10;x=-52580000;
#10;x=-52570000;
#10;x=-52560000;
#10;x=-52550000;
#10;x=-52540000;
#10;x=-52530000;
#10;x=-52520000;
#10;x=-52510000;
#10;x=-52500000;
#10;x=-52490000;
#10;x=-52480000;
#10;x=-52470000;
#10;x=-52460000;
#10;x=-52450000;
#10;x=-52440000;
#10;x=-52430000;
#10;x=-52420000;
#10;x=-52410000;
#10;x=-52400000;
#10;x=-52390000;
#10;x=-52380000;
#10;x=-52370000;
#10;x=-52360000;
#10;x=-52350000;
#10;x=-52340000;
#10;x=-52330000;
#10;x=-52320000;
#10;x=-52310000;
#10;x=-52300000;
#10;x=-52290000;
#10;x=-52280000;
#10;x=-52270000;
#10;x=-52260000;
#10;x=-52250000;
#10;x=-52240000;
#10;x=-52230000;
#10;x=-52220000;
#10;x=-52210000;
#10;x=-52200000;
#10;x=-52190000;
#10;x=-52180000;
#10;x=-52170000;
#10;x=-52160000;
#10;x=-52150000;
#10;x=-52140000;
#10;x=-52130000;
#10;x=-52120000;
#10;x=-52110000;
#10;x=-52100000;
#10;x=-52090000;
#10;x=-52080000;
#10;x=-52070000;
#10;x=-52060000;
#10;x=-52050000;
#10;x=-52040000;
#10;x=-52030000;
#10;x=-52020000;
#10;x=-52010000;
#10;x=-52000000;
#10;x=-51990000;
#10;x=-51980000;
#10;x=-51970000;
#10;x=-51960000;
#10;x=-51950000;
#10;x=-51940000;
#10;x=-51930000;
#10;x=-51920000;
#10;x=-51910000;
#10;x=-51900000;
#10;x=-51890000;
#10;x=-51880000;
#10;x=-51870000;
#10;x=-51860000;
#10;x=-51850000;
#10;x=-51840000;
#10;x=-51830000;
#10;x=-51820000;
#10;x=-51810000;
#10;x=-51800000;
#10;x=-51790000;
#10;x=-51780000;
#10;x=-51770000;
#10;x=-51760000;
#10;x=-51750000;
#10;x=-51740000;
#10;x=-51730000;
#10;x=-51720000;
#10;x=-51710000;
#10;x=-51700000;
#10;x=-51690000;
#10;x=-51680000;
#10;x=-51670000;
#10;x=-51660000;
#10;x=-51650000;
#10;x=-51640000;
#10;x=-51630000;
#10;x=-51620000;
#10;x=-51610000;
#10;x=-51600000;
#10;x=-51590000;
#10;x=-51580000;
#10;x=-51570000;
#10;x=-51560000;
#10;x=-51550000;
#10;x=-51540000;
#10;x=-51530000;
#10;x=-51520000;
#10;x=-51510000;
#10;x=-51500000;
#10;x=-51490000;
#10;x=-51480000;
#10;x=-51470000;
#10;x=-51460000;
#10;x=-51450000;
#10;x=-51440000;
#10;x=-51430000;
#10;x=-51420000;
#10;x=-51410000;
#10;x=-51400000;
#10;x=-51390000;
#10;x=-51380000;
#10;x=-51370000;
#10;x=-51360000;
#10;x=-51350000;
#10;x=-51340000;
#10;x=-51330000;
#10;x=-51320000;
#10;x=-51310000;
#10;x=-51300000;
#10;x=-51290000;
#10;x=-51280000;
#10;x=-51270000;
#10;x=-51260000;
#10;x=-51250000;
#10;x=-51240000;
#10;x=-51230000;
#10;x=-51220000;
#10;x=-51210000;
#10;x=-51200000;
#10;x=-51190000;
#10;x=-51180000;
#10;x=-51170000;
#10;x=-51160000;
#10;x=-51150000;
#10;x=-51140000;
#10;x=-51130000;
#10;x=-51120000;
#10;x=-51110000;
#10;x=-51100000;
#10;x=-51090000;
#10;x=-51080000;
#10;x=-51070000;
#10;x=-51060000;
#10;x=-51050000;
#10;x=-51040000;
#10;x=-51030000;
#10;x=-51020000;
#10;x=-51010000;
#10;x=-51000000;
#10;x=-50990000;
#10;x=-50980000;
#10;x=-50970000;
#10;x=-50960000;
#10;x=-50950000;
#10;x=-50940000;
#10;x=-50930000;
#10;x=-50920000;
#10;x=-50910000;
#10;x=-50900000;
#10;x=-50890000;
#10;x=-50880000;
#10;x=-50870000;
#10;x=-50860000;
#10;x=-50850000;
#10;x=-50840000;
#10;x=-50830000;
#10;x=-50820000;
#10;x=-50810000;
#10;x=-50800000;
#10;x=-50790000;
#10;x=-50780000;
#10;x=-50770000;
#10;x=-50760000;
#10;x=-50750000;
#10;x=-50740000;
#10;x=-50730000;
#10;x=-50720000;
#10;x=-50710000;
#10;x=-50700000;
#10;x=-50690000;
#10;x=-50680000;
#10;x=-50670000;
#10;x=-50660000;
#10;x=-50650000;
#10;x=-50640000;
#10;x=-50630000;
#10;x=-50620000;
#10;x=-50610000;
#10;x=-50600000;
#10;x=-50590000;
#10;x=-50580000;
#10;x=-50570000;
#10;x=-50560000;
#10;x=-50550000;
#10;x=-50540000;
#10;x=-50530000;
#10;x=-50520000;
#10;x=-50510000;
#10;x=-50500000;
#10;x=-50490000;
#10;x=-50480000;
#10;x=-50470000;
#10;x=-50460000;
#10;x=-50450000;
#10;x=-50440000;
#10;x=-50430000;
#10;x=-50420000;
#10;x=-50410000;
#10;x=-50400000;
#10;x=-50390000;
#10;x=-50380000;
#10;x=-50370000;
#10;x=-50360000;
#10;x=-50350000;
#10;x=-50340000;
#10;x=-50330000;
#10;x=-50320000;
#10;x=-50310000;
#10;x=-50300000;
#10;x=-50290000;
#10;x=-50280000;
#10;x=-50270000;
#10;x=-50260000;
#10;x=-50250000;
#10;x=-50240000;
#10;x=-50230000;
#10;x=-50220000;
#10;x=-50210000;
#10;x=-50200000;
#10;x=-50190000;
#10;x=-50180000;
#10;x=-50170000;
#10;x=-50160000;
#10;x=-50150000;
#10;x=-50140000;
#10;x=-50130000;
#10;x=-50120000;
#10;x=-50110000;
#10;x=-50100000;
#10;x=-50090000;
#10;x=-50080000;
#10;x=-50070000;
#10;x=-50060000;
#10;x=-50050000;
#10;x=-50040000;
#10;x=-50030000;
#10;x=-50020000;
#10;x=-50010000;
#10;x=-50000000;
#10;x=-49990000;
#10;x=-49980000;
#10;x=-49970000;
#10;x=-49960000;
#10;x=-49950000;
#10;x=-49940000;
#10;x=-49930000;
#10;x=-49920000;
#10;x=-49910000;
#10;x=-49900000;
#10;x=-49890000;
#10;x=-49880000;
#10;x=-49870000;
#10;x=-49860000;
#10;x=-49850000;
#10;x=-49840000;
#10;x=-49830000;
#10;x=-49820000;
#10;x=-49810000;
#10;x=-49800000;
#10;x=-49790000;
#10;x=-49780000;
#10;x=-49770000;
#10;x=-49760000;
#10;x=-49750000;
#10;x=-49740000;
#10;x=-49730000;
#10;x=-49720000;
#10;x=-49710000;
#10;x=-49700000;
#10;x=-49690000;
#10;x=-49680000;
#10;x=-49670000;
#10;x=-49660000;
#10;x=-49650000;
#10;x=-49640000;
#10;x=-49630000;
#10;x=-49620000;
#10;x=-49610000;
#10;x=-49600000;
#10;x=-49590000;
#10;x=-49580000;
#10;x=-49570000;
#10;x=-49560000;
#10;x=-49550000;
#10;x=-49540000;
#10;x=-49530000;
#10;x=-49520000;
#10;x=-49510000;
#10;x=-49500000;
#10;x=-49490000;
#10;x=-49480000;
#10;x=-49470000;
#10;x=-49460000;
#10;x=-49450000;
#10;x=-49440000;
#10;x=-49430000;
#10;x=-49420000;
#10;x=-49410000;
#10;x=-49400000;
#10;x=-49390000;
#10;x=-49380000;
#10;x=-49370000;
#10;x=-49360000;
#10;x=-49350000;
#10;x=-49340000;
#10;x=-49330000;
#10;x=-49320000;
#10;x=-49310000;
#10;x=-49300000;
#10;x=-49290000;
#10;x=-49280000;
#10;x=-49270000;
#10;x=-49260000;
#10;x=-49250000;
#10;x=-49240000;
#10;x=-49230000;
#10;x=-49220000;
#10;x=-49210000;
#10;x=-49200000;
#10;x=-49190000;
#10;x=-49180000;
#10;x=-49170000;
#10;x=-49160000;
#10;x=-49150000;
#10;x=-49140000;
#10;x=-49130000;
#10;x=-49120000;
#10;x=-49110000;
#10;x=-49100000;
#10;x=-49090000;
#10;x=-49080000;
#10;x=-49070000;
#10;x=-49060000;
#10;x=-49050000;
#10;x=-49040000;
#10;x=-49030000;
#10;x=-49020000;
#10;x=-49010000;
#10;x=-49000000;
#10;x=-48990000;
#10;x=-48980000;
#10;x=-48970000;
#10;x=-48960000;
#10;x=-48950000;
#10;x=-48940000;
#10;x=-48930000;
#10;x=-48920000;
#10;x=-48910000;
#10;x=-48900000;
#10;x=-48890000;
#10;x=-48880000;
#10;x=-48870000;
#10;x=-48860000;
#10;x=-48850000;
#10;x=-48840000;
#10;x=-48830000;
#10;x=-48820000;
#10;x=-48810000;
#10;x=-48800000;
#10;x=-48790000;
#10;x=-48780000;
#10;x=-48770000;
#10;x=-48760000;
#10;x=-48750000;
#10;x=-48740000;
#10;x=-48730000;
#10;x=-48720000;
#10;x=-48710000;
#10;x=-48700000;
#10;x=-48690000;
#10;x=-48680000;
#10;x=-48670000;
#10;x=-48660000;
#10;x=-48650000;
#10;x=-48640000;
#10;x=-48630000;
#10;x=-48620000;
#10;x=-48610000;
#10;x=-48600000;
#10;x=-48590000;
#10;x=-48580000;
#10;x=-48570000;
#10;x=-48560000;
#10;x=-48550000;
#10;x=-48540000;
#10;x=-48530000;
#10;x=-48520000;
#10;x=-48510000;
#10;x=-48500000;
#10;x=-48490000;
#10;x=-48480000;
#10;x=-48470000;
#10;x=-48460000;
#10;x=-48450000;
#10;x=-48440000;
#10;x=-48430000;
#10;x=-48420000;
#10;x=-48410000;
#10;x=-48400000;
#10;x=-48390000;
#10;x=-48380000;
#10;x=-48370000;
#10;x=-48360000;
#10;x=-48350000;
#10;x=-48340000;
#10;x=-48330000;
#10;x=-48320000;
#10;x=-48310000;
#10;x=-48300000;
#10;x=-48290000;
#10;x=-48280000;
#10;x=-48270000;
#10;x=-48260000;
#10;x=-48250000;
#10;x=-48240000;
#10;x=-48230000;
#10;x=-48220000;
#10;x=-48210000;
#10;x=-48200000;
#10;x=-48190000;
#10;x=-48180000;
#10;x=-48170000;
#10;x=-48160000;
#10;x=-48150000;
#10;x=-48140000;
#10;x=-48130000;
#10;x=-48120000;
#10;x=-48110000;
#10;x=-48100000;
#10;x=-48090000;
#10;x=-48080000;
#10;x=-48070000;
#10;x=-48060000;
#10;x=-48050000;
#10;x=-48040000;
#10;x=-48030000;
#10;x=-48020000;
#10;x=-48010000;
#10;x=-48000000;
#10;x=-47990000;
#10;x=-47980000;
#10;x=-47970000;
#10;x=-47960000;
#10;x=-47950000;
#10;x=-47940000;
#10;x=-47930000;
#10;x=-47920000;
#10;x=-47910000;
#10;x=-47900000;
#10;x=-47890000;
#10;x=-47880000;
#10;x=-47870000;
#10;x=-47860000;
#10;x=-47850000;
#10;x=-47840000;
#10;x=-47830000;
#10;x=-47820000;
#10;x=-47810000;
#10;x=-47800000;
#10;x=-47790000;
#10;x=-47780000;
#10;x=-47770000;
#10;x=-47760000;
#10;x=-47750000;
#10;x=-47740000;
#10;x=-47730000;
#10;x=-47720000;
#10;x=-47710000;
#10;x=-47700000;
#10;x=-47690000;
#10;x=-47680000;
#10;x=-47670000;
#10;x=-47660000;
#10;x=-47650000;
#10;x=-47640000;
#10;x=-47630000;
#10;x=-47620000;
#10;x=-47610000;
#10;x=-47600000;
#10;x=-47590000;
#10;x=-47580000;
#10;x=-47570000;
#10;x=-47560000;
#10;x=-47550000;
#10;x=-47540000;
#10;x=-47530000;
#10;x=-47520000;
#10;x=-47510000;
#10;x=-47500000;
#10;x=-47490000;
#10;x=-47480000;
#10;x=-47470000;
#10;x=-47460000;
#10;x=-47450000;
#10;x=-47440000;
#10;x=-47430000;
#10;x=-47420000;
#10;x=-47410000;
#10;x=-47400000;
#10;x=-47390000;
#10;x=-47380000;
#10;x=-47370000;
#10;x=-47360000;
#10;x=-47350000;
#10;x=-47340000;
#10;x=-47330000;
#10;x=-47320000;
#10;x=-47310000;
#10;x=-47300000;
#10;x=-47290000;
#10;x=-47280000;
#10;x=-47270000;
#10;x=-47260000;
#10;x=-47250000;
#10;x=-47240000;
#10;x=-47230000;
#10;x=-47220000;
#10;x=-47210000;
#10;x=-47200000;
#10;x=-47190000;
#10;x=-47180000;
#10;x=-47170000;
#10;x=-47160000;
#10;x=-47150000;
#10;x=-47140000;
#10;x=-47130000;
#10;x=-47120000;
#10;x=-47110000;
#10;x=-47100000;
#10;x=-47090000;
#10;x=-47080000;
#10;x=-47070000;
#10;x=-47060000;
#10;x=-47050000;
#10;x=-47040000;
#10;x=-47030000;
#10;x=-47020000;
#10;x=-47010000;
#10;x=-47000000;
#10;x=-46990000;
#10;x=-46980000;
#10;x=-46970000;
#10;x=-46960000;
#10;x=-46950000;
#10;x=-46940000;
#10;x=-46930000;
#10;x=-46920000;
#10;x=-46910000;
#10;x=-46900000;
#10;x=-46890000;
#10;x=-46880000;
#10;x=-46870000;
#10;x=-46860000;
#10;x=-46850000;
#10;x=-46840000;
#10;x=-46830000;
#10;x=-46820000;
#10;x=-46810000;
#10;x=-46800000;
#10;x=-46790000;
#10;x=-46780000;
#10;x=-46770000;
#10;x=-46760000;
#10;x=-46750000;
#10;x=-46740000;
#10;x=-46730000;
#10;x=-46720000;
#10;x=-46710000;
#10;x=-46700000;
#10;x=-46690000;
#10;x=-46680000;
#10;x=-46670000;
#10;x=-46660000;
#10;x=-46650000;
#10;x=-46640000;
#10;x=-46630000;
#10;x=-46620000;
#10;x=-46610000;
#10;x=-46600000;
#10;x=-46590000;
#10;x=-46580000;
#10;x=-46570000;
#10;x=-46560000;
#10;x=-46550000;
#10;x=-46540000;
#10;x=-46530000;
#10;x=-46520000;
#10;x=-46510000;
#10;x=-46500000;
#10;x=-46490000;
#10;x=-46480000;
#10;x=-46470000;
#10;x=-46460000;
#10;x=-46450000;
#10;x=-46440000;
#10;x=-46430000;
#10;x=-46420000;
#10;x=-46410000;
#10;x=-46400000;
#10;x=-46390000;
#10;x=-46380000;
#10;x=-46370000;
#10;x=-46360000;
#10;x=-46350000;
#10;x=-46340000;
#10;x=-46330000;
#10;x=-46320000;
#10;x=-46310000;
#10;x=-46300000;
#10;x=-46290000;
#10;x=-46280000;
#10;x=-46270000;
#10;x=-46260000;
#10;x=-46250000;
#10;x=-46240000;
#10;x=-46230000;
#10;x=-46220000;
#10;x=-46210000;
#10;x=-46200000;
#10;x=-46190000;
#10;x=-46180000;
#10;x=-46170000;
#10;x=-46160000;
#10;x=-46150000;
#10;x=-46140000;
#10;x=-46130000;
#10;x=-46120000;
#10;x=-46110000;
#10;x=-46100000;
#10;x=-46090000;
#10;x=-46080000;
#10;x=-46070000;
#10;x=-46060000;
#10;x=-46050000;
#10;x=-46040000;
#10;x=-46030000;
#10;x=-46020000;
#10;x=-46010000;
#10;x=-46000000;
#10;x=-45990000;
#10;x=-45980000;
#10;x=-45970000;
#10;x=-45960000;
#10;x=-45950000;
#10;x=-45940000;
#10;x=-45930000;
#10;x=-45920000;
#10;x=-45910000;
#10;x=-45900000;
#10;x=-45890000;
#10;x=-45880000;
#10;x=-45870000;
#10;x=-45860000;
#10;x=-45850000;
#10;x=-45840000;
#10;x=-45830000;
#10;x=-45820000;
#10;x=-45810000;
#10;x=-45800000;
#10;x=-45790000;
#10;x=-45780000;
#10;x=-45770000;
#10;x=-45760000;
#10;x=-45750000;
#10;x=-45740000;
#10;x=-45730000;
#10;x=-45720000;
#10;x=-45710000;
#10;x=-45700000;
#10;x=-45690000;
#10;x=-45680000;
#10;x=-45670000;
#10;x=-45660000;
#10;x=-45650000;
#10;x=-45640000;
#10;x=-45630000;
#10;x=-45620000;
#10;x=-45610000;
#10;x=-45600000;
#10;x=-45590000;
#10;x=-45580000;
#10;x=-45570000;
#10;x=-45560000;
#10;x=-45550000;
#10;x=-45540000;
#10;x=-45530000;
#10;x=-45520000;
#10;x=-45510000;
#10;x=-45500000;
#10;x=-45490000;
#10;x=-45480000;
#10;x=-45470000;
#10;x=-45460000;
#10;x=-45450000;
#10;x=-45440000;
#10;x=-45430000;
#10;x=-45420000;
#10;x=-45410000;
#10;x=-45400000;
#10;x=-45390000;
#10;x=-45380000;
#10;x=-45370000;
#10;x=-45360000;
#10;x=-45350000;
#10;x=-45340000;
#10;x=-45330000;
#10;x=-45320000;
#10;x=-45310000;
#10;x=-45300000;
#10;x=-45290000;
#10;x=-45280000;
#10;x=-45270000;
#10;x=-45260000;
#10;x=-45250000;
#10;x=-45240000;
#10;x=-45230000;
#10;x=-45220000;
#10;x=-45210000;
#10;x=-45200000;
#10;x=-45190000;
#10;x=-45180000;
#10;x=-45170000;
#10;x=-45160000;
#10;x=-45150000;
#10;x=-45140000;
#10;x=-45130000;
#10;x=-45120000;
#10;x=-45110000;
#10;x=-45100000;
#10;x=-45090000;
#10;x=-45080000;
#10;x=-45070000;
#10;x=-45060000;
#10;x=-45050000;
#10;x=-45040000;
#10;x=-45030000;
#10;x=-45020000;
#10;x=-45010000;
#10;x=-45000000;
#10;x=-44990000;
#10;x=-44980000;
#10;x=-44970000;
#10;x=-44960000;
#10;x=-44950000;
#10;x=-44940000;
#10;x=-44930000;
#10;x=-44920000;
#10;x=-44910000;
#10;x=-44900000;
#10;x=-44890000;
#10;x=-44880000;
#10;x=-44870000;
#10;x=-44860000;
#10;x=-44850000;
#10;x=-44840000;
#10;x=-44830000;
#10;x=-44820000;
#10;x=-44810000;
#10;x=-44800000;
#10;x=-44790000;
#10;x=-44780000;
#10;x=-44770000;
#10;x=-44760000;
#10;x=-44750000;
#10;x=-44740000;
#10;x=-44730000;
#10;x=-44720000;
#10;x=-44710000;
#10;x=-44700000;
#10;x=-44690000;
#10;x=-44680000;
#10;x=-44670000;
#10;x=-44660000;
#10;x=-44650000;
#10;x=-44640000;
#10;x=-44630000;
#10;x=-44620000;
#10;x=-44610000;
#10;x=-44600000;
#10;x=-44590000;
#10;x=-44580000;
#10;x=-44570000;
#10;x=-44560000;
#10;x=-44550000;
#10;x=-44540000;
#10;x=-44530000;
#10;x=-44520000;
#10;x=-44510000;
#10;x=-44500000;
#10;x=-44490000;
#10;x=-44480000;
#10;x=-44470000;
#10;x=-44460000;
#10;x=-44450000;
#10;x=-44440000;
#10;x=-44430000;
#10;x=-44420000;
#10;x=-44410000;
#10;x=-44400000;
#10;x=-44390000;
#10;x=-44380000;
#10;x=-44370000;
#10;x=-44360000;
#10;x=-44350000;
#10;x=-44340000;
#10;x=-44330000;
#10;x=-44320000;
#10;x=-44310000;
#10;x=-44300000;
#10;x=-44290000;
#10;x=-44280000;
#10;x=-44270000;
#10;x=-44260000;
#10;x=-44250000;
#10;x=-44240000;
#10;x=-44230000;
#10;x=-44220000;
#10;x=-44210000;
#10;x=-44200000;
#10;x=-44190000;
#10;x=-44180000;
#10;x=-44170000;
#10;x=-44160000;
#10;x=-44150000;
#10;x=-44140000;
#10;x=-44130000;
#10;x=-44120000;
#10;x=-44110000;
#10;x=-44100000;
#10;x=-44090000;
#10;x=-44080000;
#10;x=-44070000;
#10;x=-44060000;
#10;x=-44050000;
#10;x=-44040000;
#10;x=-44030000;
#10;x=-44020000;
#10;x=-44010000;
#10;x=-44000000;
#10;x=-43990000;
#10;x=-43980000;
#10;x=-43970000;
#10;x=-43960000;
#10;x=-43950000;
#10;x=-43940000;
#10;x=-43930000;
#10;x=-43920000;
#10;x=-43910000;
#10;x=-43900000;
#10;x=-43890000;
#10;x=-43880000;
#10;x=-43870000;
#10;x=-43860000;
#10;x=-43850000;
#10;x=-43840000;
#10;x=-43830000;
#10;x=-43820000;
#10;x=-43810000;
#10;x=-43800000;
#10;x=-43790000;
#10;x=-43780000;
#10;x=-43770000;
#10;x=-43760000;
#10;x=-43750000;
#10;x=-43740000;
#10;x=-43730000;
#10;x=-43720000;
#10;x=-43710000;
#10;x=-43700000;
#10;x=-43690000;
#10;x=-43680000;
#10;x=-43670000;
#10;x=-43660000;
#10;x=-43650000;
#10;x=-43640000;
#10;x=-43630000;
#10;x=-43620000;
#10;x=-43610000;
#10;x=-43600000;
#10;x=-43590000;
#10;x=-43580000;
#10;x=-43570000;
#10;x=-43560000;
#10;x=-43550000;
#10;x=-43540000;
#10;x=-43530000;
#10;x=-43520000;
#10;x=-43510000;
#10;x=-43500000;
#10;x=-43490000;
#10;x=-43480000;
#10;x=-43470000;
#10;x=-43460000;
#10;x=-43450000;
#10;x=-43440000;
#10;x=-43430000;
#10;x=-43420000;
#10;x=-43410000;
#10;x=-43400000;
#10;x=-43390000;
#10;x=-43380000;
#10;x=-43370000;
#10;x=-43360000;
#10;x=-43350000;
#10;x=-43340000;
#10;x=-43330000;
#10;x=-43320000;
#10;x=-43310000;
#10;x=-43300000;
#10;x=-43290000;
#10;x=-43280000;
#10;x=-43270000;
#10;x=-43260000;
#10;x=-43250000;
#10;x=-43240000;
#10;x=-43230000;
#10;x=-43220000;
#10;x=-43210000;
#10;x=-43200000;
#10;x=-43190000;
#10;x=-43180000;
#10;x=-43170000;
#10;x=-43160000;
#10;x=-43150000;
#10;x=-43140000;
#10;x=-43130000;
#10;x=-43120000;
#10;x=-43110000;
#10;x=-43100000;
#10;x=-43090000;
#10;x=-43080000;
#10;x=-43070000;
#10;x=-43060000;
#10;x=-43050000;
#10;x=-43040000;
#10;x=-43030000;
#10;x=-43020000;
#10;x=-43010000;
#10;x=-43000000;
#10;x=-42990000;
#10;x=-42980000;
#10;x=-42970000;
#10;x=-42960000;
#10;x=-42950000;
#10;x=-42940000;
#10;x=-42930000;
#10;x=-42920000;
#10;x=-42910000;
#10;x=-42900000;
#10;x=-42890000;
#10;x=-42880000;
#10;x=-42870000;
#10;x=-42860000;
#10;x=-42850000;
#10;x=-42840000;
#10;x=-42830000;
#10;x=-42820000;
#10;x=-42810000;
#10;x=-42800000;
#10;x=-42790000;
#10;x=-42780000;
#10;x=-42770000;
#10;x=-42760000;
#10;x=-42750000;
#10;x=-42740000;
#10;x=-42730000;
#10;x=-42720000;
#10;x=-42710000;
#10;x=-42700000;
#10;x=-42690000;
#10;x=-42680000;
#10;x=-42670000;
#10;x=-42660000;
#10;x=-42650000;
#10;x=-42640000;
#10;x=-42630000;
#10;x=-42620000;
#10;x=-42610000;
#10;x=-42600000;
#10;x=-42590000;
#10;x=-42580000;
#10;x=-42570000;
#10;x=-42560000;
#10;x=-42550000;
#10;x=-42540000;
#10;x=-42530000;
#10;x=-42520000;
#10;x=-42510000;
#10;x=-42500000;
#10;x=-42490000;
#10;x=-42480000;
#10;x=-42470000;
#10;x=-42460000;
#10;x=-42450000;
#10;x=-42440000;
#10;x=-42430000;
#10;x=-42420000;
#10;x=-42410000;
#10;x=-42400000;
#10;x=-42390000;
#10;x=-42380000;
#10;x=-42370000;
#10;x=-42360000;
#10;x=-42350000;
#10;x=-42340000;
#10;x=-42330000;
#10;x=-42320000;
#10;x=-42310000;
#10;x=-42300000;
#10;x=-42290000;
#10;x=-42280000;
#10;x=-42270000;
#10;x=-42260000;
#10;x=-42250000;
#10;x=-42240000;
#10;x=-42230000;
#10;x=-42220000;
#10;x=-42210000;
#10;x=-42200000;
#10;x=-42190000;
#10;x=-42180000;
#10;x=-42170000;
#10;x=-42160000;
#10;x=-42150000;
#10;x=-42140000;
#10;x=-42130000;
#10;x=-42120000;
#10;x=-42110000;
#10;x=-42100000;
#10;x=-42090000;
#10;x=-42080000;
#10;x=-42070000;
#10;x=-42060000;
#10;x=-42050000;
#10;x=-42040000;
#10;x=-42030000;
#10;x=-42020000;
#10;x=-42010000;
#10;x=-42000000;
#10;x=-41990000;
#10;x=-41980000;
#10;x=-41970000;
#10;x=-41960000;
#10;x=-41950000;
#10;x=-41940000;
#10;x=-41930000;
#10;x=-41920000;
#10;x=-41910000;
#10;x=-41900000;
#10;x=-41890000;
#10;x=-41880000;
#10;x=-41870000;
#10;x=-41860000;
#10;x=-41850000;
#10;x=-41840000;
#10;x=-41830000;
#10;x=-41820000;
#10;x=-41810000;
#10;x=-41800000;
#10;x=-41790000;
#10;x=-41780000;
#10;x=-41770000;
#10;x=-41760000;
#10;x=-41750000;
#10;x=-41740000;
#10;x=-41730000;
#10;x=-41720000;
#10;x=-41710000;
#10;x=-41700000;
#10;x=-41690000;
#10;x=-41680000;
#10;x=-41670000;
#10;x=-41660000;
#10;x=-41650000;
#10;x=-41640000;
#10;x=-41630000;
#10;x=-41620000;
#10;x=-41610000;
#10;x=-41600000;
#10;x=-41590000;
#10;x=-41580000;
#10;x=-41570000;
#10;x=-41560000;
#10;x=-41550000;
#10;x=-41540000;
#10;x=-41530000;
#10;x=-41520000;
#10;x=-41510000;
#10;x=-41500000;
#10;x=-41490000;
#10;x=-41480000;
#10;x=-41470000;
#10;x=-41460000;
#10;x=-41450000;
#10;x=-41440000;
#10;x=-41430000;
#10;x=-41420000;
#10;x=-41410000;
#10;x=-41400000;
#10;x=-41390000;
#10;x=-41380000;
#10;x=-41370000;
#10;x=-41360000;
#10;x=-41350000;
#10;x=-41340000;
#10;x=-41330000;
#10;x=-41320000;
#10;x=-41310000;
#10;x=-41300000;
#10;x=-41290000;
#10;x=-41280000;
#10;x=-41270000;
#10;x=-41260000;
#10;x=-41250000;
#10;x=-41240000;
#10;x=-41230000;
#10;x=-41220000;
#10;x=-41210000;
#10;x=-41200000;
#10;x=-41190000;
#10;x=-41180000;
#10;x=-41170000;
#10;x=-41160000;
#10;x=-41150000;
#10;x=-41140000;
#10;x=-41130000;
#10;x=-41120000;
#10;x=-41110000;
#10;x=-41100000;
#10;x=-41090000;
#10;x=-41080000;
#10;x=-41070000;
#10;x=-41060000;
#10;x=-41050000;
#10;x=-41040000;
#10;x=-41030000;
#10;x=-41020000;
#10;x=-41010000;
#10;x=-41000000;
#10;x=-40990000;
#10;x=-40980000;
#10;x=-40970000;
#10;x=-40960000;
#10;x=-40950000;
#10;x=-40940000;
#10;x=-40930000;
#10;x=-40920000;
#10;x=-40910000;
#10;x=-40900000;
#10;x=-40890000;
#10;x=-40880000;
#10;x=-40870000;
#10;x=-40860000;
#10;x=-40850000;
#10;x=-40840000;
#10;x=-40830000;
#10;x=-40820000;
#10;x=-40810000;
#10;x=-40800000;
#10;x=-40790000;
#10;x=-40780000;
#10;x=-40770000;
#10;x=-40760000;
#10;x=-40750000;
#10;x=-40740000;
#10;x=-40730000;
#10;x=-40720000;
#10;x=-40710000;
#10;x=-40700000;
#10;x=-40690000;
#10;x=-40680000;
#10;x=-40670000;
#10;x=-40660000;
#10;x=-40650000;
#10;x=-40640000;
#10;x=-40630000;
#10;x=-40620000;
#10;x=-40610000;
#10;x=-40600000;
#10;x=-40590000;
#10;x=-40580000;
#10;x=-40570000;
#10;x=-40560000;
#10;x=-40550000;
#10;x=-40540000;
#10;x=-40530000;
#10;x=-40520000;
#10;x=-40510000;
#10;x=-40500000;
#10;x=-40490000;
#10;x=-40480000;
#10;x=-40470000;
#10;x=-40460000;
#10;x=-40450000;
#10;x=-40440000;
#10;x=-40430000;
#10;x=-40420000;
#10;x=-40410000;
#10;x=-40400000;
#10;x=-40390000;
#10;x=-40380000;
#10;x=-40370000;
#10;x=-40360000;
#10;x=-40350000;
#10;x=-40340000;
#10;x=-40330000;
#10;x=-40320000;
#10;x=-40310000;
#10;x=-40300000;
#10;x=-40290000;
#10;x=-40280000;
#10;x=-40270000;
#10;x=-40260000;
#10;x=-40250000;
#10;x=-40240000;
#10;x=-40230000;
#10;x=-40220000;
#10;x=-40210000;
#10;x=-40200000;
#10;x=-40190000;
#10;x=-40180000;
#10;x=-40170000;
#10;x=-40160000;
#10;x=-40150000;
#10;x=-40140000;
#10;x=-40130000;
#10;x=-40120000;
#10;x=-40110000;
#10;x=-40100000;
#10;x=-40090000;
#10;x=-40080000;
#10;x=-40070000;
#10;x=-40060000;
#10;x=-40050000;
#10;x=-40040000;
#10;x=-40030000;
#10;x=-40020000;
#10;x=-40010000;
#10;x=-40000000;
#10;x=-39990000;
#10;x=-39980000;
#10;x=-39970000;
#10;x=-39960000;
#10;x=-39950000;
#10;x=-39940000;
#10;x=-39930000;
#10;x=-39920000;
#10;x=-39910000;
#10;x=-39900000;
#10;x=-39890000;
#10;x=-39880000;
#10;x=-39870000;
#10;x=-39860000;
#10;x=-39850000;
#10;x=-39840000;
#10;x=-39830000;
#10;x=-39820000;
#10;x=-39810000;
#10;x=-39800000;
#10;x=-39790000;
#10;x=-39780000;
#10;x=-39770000;
#10;x=-39760000;
#10;x=-39750000;
#10;x=-39740000;
#10;x=-39730000;
#10;x=-39720000;
#10;x=-39710000;
#10;x=-39700000;
#10;x=-39690000;
#10;x=-39680000;
#10;x=-39670000;
#10;x=-39660000;
#10;x=-39650000;
#10;x=-39640000;
#10;x=-39630000;
#10;x=-39620000;
#10;x=-39610000;
#10;x=-39600000;
#10;x=-39590000;
#10;x=-39580000;
#10;x=-39570000;
#10;x=-39560000;
#10;x=-39550000;
#10;x=-39540000;
#10;x=-39530000;
#10;x=-39520000;
#10;x=-39510000;
#10;x=-39500000;
#10;x=-39490000;
#10;x=-39480000;
#10;x=-39470000;
#10;x=-39460000;
#10;x=-39450000;
#10;x=-39440000;
#10;x=-39430000;
#10;x=-39420000;
#10;x=-39410000;
#10;x=-39400000;
#10;x=-39390000;
#10;x=-39380000;
#10;x=-39370000;
#10;x=-39360000;
#10;x=-39350000;
#10;x=-39340000;
#10;x=-39330000;
#10;x=-39320000;
#10;x=-39310000;
#10;x=-39300000;
#10;x=-39290000;
#10;x=-39280000;
#10;x=-39270000;
#10;x=-39260000;
#10;x=-39250000;
#10;x=-39240000;
#10;x=-39230000;
#10;x=-39220000;
#10;x=-39210000;
#10;x=-39200000;
#10;x=-39190000;
#10;x=-39180000;
#10;x=-39170000;
#10;x=-39160000;
#10;x=-39150000;
#10;x=-39140000;
#10;x=-39130000;
#10;x=-39120000;
#10;x=-39110000;
#10;x=-39100000;
#10;x=-39090000;
#10;x=-39080000;
#10;x=-39070000;
#10;x=-39060000;
#10;x=-39050000;
#10;x=-39040000;
#10;x=-39030000;
#10;x=-39020000;
#10;x=-39010000;
#10;x=-39000000;
#10;x=-38990000;
#10;x=-38980000;
#10;x=-38970000;
#10;x=-38960000;
#10;x=-38950000;
#10;x=-38940000;
#10;x=-38930000;
#10;x=-38920000;
#10;x=-38910000;
#10;x=-38900000;
#10;x=-38890000;
#10;x=-38880000;
#10;x=-38870000;
#10;x=-38860000;
#10;x=-38850000;
#10;x=-38840000;
#10;x=-38830000;
#10;x=-38820000;
#10;x=-38810000;
#10;x=-38800000;
#10;x=-38790000;
#10;x=-38780000;
#10;x=-38770000;
#10;x=-38760000;
#10;x=-38750000;
#10;x=-38740000;
#10;x=-38730000;
#10;x=-38720000;
#10;x=-38710000;
#10;x=-38700000;
#10;x=-38690000;
#10;x=-38680000;
#10;x=-38670000;
#10;x=-38660000;
#10;x=-38650000;
#10;x=-38640000;
#10;x=-38630000;
#10;x=-38620000;
#10;x=-38610000;
#10;x=-38600000;
#10;x=-38590000;
#10;x=-38580000;
#10;x=-38570000;
#10;x=-38560000;
#10;x=-38550000;
#10;x=-38540000;
#10;x=-38530000;
#10;x=-38520000;
#10;x=-38510000;
#10;x=-38500000;
#10;x=-38490000;
#10;x=-38480000;
#10;x=-38470000;
#10;x=-38460000;
#10;x=-38450000;
#10;x=-38440000;
#10;x=-38430000;
#10;x=-38420000;
#10;x=-38410000;
#10;x=-38400000;
#10;x=-38390000;
#10;x=-38380000;
#10;x=-38370000;
#10;x=-38360000;
#10;x=-38350000;
#10;x=-38340000;
#10;x=-38330000;
#10;x=-38320000;
#10;x=-38310000;
#10;x=-38300000;
#10;x=-38290000;
#10;x=-38280000;
#10;x=-38270000;
#10;x=-38260000;
#10;x=-38250000;
#10;x=-38240000;
#10;x=-38230000;
#10;x=-38220000;
#10;x=-38210000;
#10;x=-38200000;
#10;x=-38190000;
#10;x=-38180000;
#10;x=-38170000;
#10;x=-38160000;
#10;x=-38150000;
#10;x=-38140000;
#10;x=-38130000;
#10;x=-38120000;
#10;x=-38110000;
#10;x=-38100000;
#10;x=-38090000;
#10;x=-38080000;
#10;x=-38070000;
#10;x=-38060000;
#10;x=-38050000;
#10;x=-38040000;
#10;x=-38030000;
#10;x=-38020000;
#10;x=-38010000;
#10;x=-38000000;
#10;x=-37990000;
#10;x=-37980000;
#10;x=-37970000;
#10;x=-37960000;
#10;x=-37950000;
#10;x=-37940000;
#10;x=-37930000;
#10;x=-37920000;
#10;x=-37910000;
#10;x=-37900000;
#10;x=-37890000;
#10;x=-37880000;
#10;x=-37870000;
#10;x=-37860000;
#10;x=-37850000;
#10;x=-37840000;
#10;x=-37830000;
#10;x=-37820000;
#10;x=-37810000;
#10;x=-37800000;
#10;x=-37790000;
#10;x=-37780000;
#10;x=-37770000;
#10;x=-37760000;
#10;x=-37750000;
#10;x=-37740000;
#10;x=-37730000;
#10;x=-37720000;
#10;x=-37710000;
#10;x=-37700000;
#10;x=-37690000;
#10;x=-37680000;
#10;x=-37670000;
#10;x=-37660000;
#10;x=-37650000;
#10;x=-37640000;
#10;x=-37630000;
#10;x=-37620000;
#10;x=-37610000;
#10;x=-37600000;
#10;x=-37590000;
#10;x=-37580000;
#10;x=-37570000;
#10;x=-37560000;
#10;x=-37550000;
#10;x=-37540000;
#10;x=-37530000;
#10;x=-37520000;
#10;x=-37510000;
#10;x=-37500000;
#10;x=-37490000;
#10;x=-37480000;
#10;x=-37470000;
#10;x=-37460000;
#10;x=-37450000;
#10;x=-37440000;
#10;x=-37430000;
#10;x=-37420000;
#10;x=-37410000;
#10;x=-37400000;
#10;x=-37390000;
#10;x=-37380000;
#10;x=-37370000;
#10;x=-37360000;
#10;x=-37350000;
#10;x=-37340000;
#10;x=-37330000;
#10;x=-37320000;
#10;x=-37310000;
#10;x=-37300000;
#10;x=-37290000;
#10;x=-37280000;
#10;x=-37270000;
#10;x=-37260000;
#10;x=-37250000;
#10;x=-37240000;
#10;x=-37230000;
#10;x=-37220000;
#10;x=-37210000;
#10;x=-37200000;
#10;x=-37190000;
#10;x=-37180000;
#10;x=-37170000;
#10;x=-37160000;
#10;x=-37150000;
#10;x=-37140000;
#10;x=-37130000;
#10;x=-37120000;
#10;x=-37110000;
#10;x=-37100000;
#10;x=-37090000;
#10;x=-37080000;
#10;x=-37070000;
#10;x=-37060000;
#10;x=-37050000;
#10;x=-37040000;
#10;x=-37030000;
#10;x=-37020000;
#10;x=-37010000;
#10;x=-37000000;
#10;x=-36990000;
#10;x=-36980000;
#10;x=-36970000;
#10;x=-36960000;
#10;x=-36950000;
#10;x=-36940000;
#10;x=-36930000;
#10;x=-36920000;
#10;x=-36910000;
#10;x=-36900000;
#10;x=-36890000;
#10;x=-36880000;
#10;x=-36870000;
#10;x=-36860000;
#10;x=-36850000;
#10;x=-36840000;
#10;x=-36830000;
#10;x=-36820000;
#10;x=-36810000;
#10;x=-36800000;
#10;x=-36790000;
#10;x=-36780000;
#10;x=-36770000;
#10;x=-36760000;
#10;x=-36750000;
#10;x=-36740000;
#10;x=-36730000;
#10;x=-36720000;
#10;x=-36710000;
#10;x=-36700000;
#10;x=-36690000;
#10;x=-36680000;
#10;x=-36670000;
#10;x=-36660000;
#10;x=-36650000;
#10;x=-36640000;
#10;x=-36630000;
#10;x=-36620000;
#10;x=-36610000;
#10;x=-36600000;
#10;x=-36590000;
#10;x=-36580000;
#10;x=-36570000;
#10;x=-36560000;
#10;x=-36550000;
#10;x=-36540000;
#10;x=-36530000;
#10;x=-36520000;
#10;x=-36510000;
#10;x=-36500000;
#10;x=-36490000;
#10;x=-36480000;
#10;x=-36470000;
#10;x=-36460000;
#10;x=-36450000;
#10;x=-36440000;
#10;x=-36430000;
#10;x=-36420000;
#10;x=-36410000;
#10;x=-36400000;
#10;x=-36390000;
#10;x=-36380000;
#10;x=-36370000;
#10;x=-36360000;
#10;x=-36350000;
#10;x=-36340000;
#10;x=-36330000;
#10;x=-36320000;
#10;x=-36310000;
#10;x=-36300000;
#10;x=-36290000;
#10;x=-36280000;
#10;x=-36270000;
#10;x=-36260000;
#10;x=-36250000;
#10;x=-36240000;
#10;x=-36230000;
#10;x=-36220000;
#10;x=-36210000;
#10;x=-36200000;
#10;x=-36190000;
#10;x=-36180000;
#10;x=-36170000;
#10;x=-36160000;
#10;x=-36150000;
#10;x=-36140000;
#10;x=-36130000;
#10;x=-36120000;
#10;x=-36110000;
#10;x=-36100000;
#10;x=-36090000;
#10;x=-36080000;
#10;x=-36070000;
#10;x=-36060000;
#10;x=-36050000;
#10;x=-36040000;
#10;x=-36030000;
#10;x=-36020000;
#10;x=-36010000;
#10;x=-36000000;
#10;x=-35990000;
#10;x=-35980000;
#10;x=-35970000;
#10;x=-35960000;
#10;x=-35950000;
#10;x=-35940000;
#10;x=-35930000;
#10;x=-35920000;
#10;x=-35910000;
#10;x=-35900000;
#10;x=-35890000;
#10;x=-35880000;
#10;x=-35870000;
#10;x=-35860000;
#10;x=-35850000;
#10;x=-35840000;
#10;x=-35830000;
#10;x=-35820000;
#10;x=-35810000;
#10;x=-35800000;
#10;x=-35790000;
#10;x=-35780000;
#10;x=-35770000;
#10;x=-35760000;
#10;x=-35750000;
#10;x=-35740000;
#10;x=-35730000;
#10;x=-35720000;
#10;x=-35710000;
#10;x=-35700000;
#10;x=-35690000;
#10;x=-35680000;
#10;x=-35670000;
#10;x=-35660000;
#10;x=-35650000;
#10;x=-35640000;
#10;x=-35630000;
#10;x=-35620000;
#10;x=-35610000;
#10;x=-35600000;
#10;x=-35590000;
#10;x=-35580000;
#10;x=-35570000;
#10;x=-35560000;
#10;x=-35550000;
#10;x=-35540000;
#10;x=-35530000;
#10;x=-35520000;
#10;x=-35510000;
#10;x=-35500000;
#10;x=-35490000;
#10;x=-35480000;
#10;x=-35470000;
#10;x=-35460000;
#10;x=-35450000;
#10;x=-35440000;
#10;x=-35430000;
#10;x=-35420000;
#10;x=-35410000;
#10;x=-35400000;
#10;x=-35390000;
#10;x=-35380000;
#10;x=-35370000;
#10;x=-35360000;
#10;x=-35350000;
#10;x=-35340000;
#10;x=-35330000;
#10;x=-35320000;
#10;x=-35310000;
#10;x=-35300000;
#10;x=-35290000;
#10;x=-35280000;
#10;x=-35270000;
#10;x=-35260000;
#10;x=-35250000;
#10;x=-35240000;
#10;x=-35230000;
#10;x=-35220000;
#10;x=-35210000;
#10;x=-35200000;
#10;x=-35190000;
#10;x=-35180000;
#10;x=-35170000;
#10;x=-35160000;
#10;x=-35150000;
#10;x=-35140000;
#10;x=-35130000;
#10;x=-35120000;
#10;x=-35110000;
#10;x=-35100000;
#10;x=-35090000;
#10;x=-35080000;
#10;x=-35070000;
#10;x=-35060000;
#10;x=-35050000;
#10;x=-35040000;
#10;x=-35030000;
#10;x=-35020000;
#10;x=-35010000;
#10;x=-35000000;
#10;x=-34990000;
#10;x=-34980000;
#10;x=-34970000;
#10;x=-34960000;
#10;x=-34950000;
#10;x=-34940000;
#10;x=-34930000;
#10;x=-34920000;
#10;x=-34910000;
#10;x=-34900000;
#10;x=-34890000;
#10;x=-34880000;
#10;x=-34870000;
#10;x=-34860000;
#10;x=-34850000;
#10;x=-34840000;
#10;x=-34830000;
#10;x=-34820000;
#10;x=-34810000;
#10;x=-34800000;
#10;x=-34790000;
#10;x=-34780000;
#10;x=-34770000;
#10;x=-34760000;
#10;x=-34750000;
#10;x=-34740000;
#10;x=-34730000;
#10;x=-34720000;
#10;x=-34710000;
#10;x=-34700000;
#10;x=-34690000;
#10;x=-34680000;
#10;x=-34670000;
#10;x=-34660000;
#10;x=-34650000;
#10;x=-34640000;
#10;x=-34630000;
#10;x=-34620000;
#10;x=-34610000;
#10;x=-34600000;
#10;x=-34590000;
#10;x=-34580000;
#10;x=-34570000;
#10;x=-34560000;
#10;x=-34550000;
#10;x=-34540000;
#10;x=-34530000;
#10;x=-34520000;
#10;x=-34510000;
#10;x=-34500000;
#10;x=-34490000;
#10;x=-34480000;
#10;x=-34470000;
#10;x=-34460000;
#10;x=-34450000;
#10;x=-34440000;
#10;x=-34430000;
#10;x=-34420000;
#10;x=-34410000;
#10;x=-34400000;
#10;x=-34390000;
#10;x=-34380000;
#10;x=-34370000;
#10;x=-34360000;
#10;x=-34350000;
#10;x=-34340000;
#10;x=-34330000;
#10;x=-34320000;
#10;x=-34310000;
#10;x=-34300000;
#10;x=-34290000;
#10;x=-34280000;
#10;x=-34270000;
#10;x=-34260000;
#10;x=-34250000;
#10;x=-34240000;
#10;x=-34230000;
#10;x=-34220000;
#10;x=-34210000;
#10;x=-34200000;
#10;x=-34190000;
#10;x=-34180000;
#10;x=-34170000;
#10;x=-34160000;
#10;x=-34150000;
#10;x=-34140000;
#10;x=-34130000;
#10;x=-34120000;
#10;x=-34110000;
#10;x=-34100000;
#10;x=-34090000;
#10;x=-34080000;
#10;x=-34070000;
#10;x=-34060000;
#10;x=-34050000;
#10;x=-34040000;
#10;x=-34030000;
#10;x=-34020000;
#10;x=-34010000;
#10;x=-34000000;
#10;x=-33990000;
#10;x=-33980000;
#10;x=-33970000;
#10;x=-33960000;
#10;x=-33950000;
#10;x=-33940000;
#10;x=-33930000;
#10;x=-33920000;
#10;x=-33910000;
#10;x=-33900000;
#10;x=-33890000;
#10;x=-33880000;
#10;x=-33870000;
#10;x=-33860000;
#10;x=-33850000;
#10;x=-33840000;
#10;x=-33830000;
#10;x=-33820000;
#10;x=-33810000;
#10;x=-33800000;
#10;x=-33790000;
#10;x=-33780000;
#10;x=-33770000;
#10;x=-33760000;
#10;x=-33750000;
#10;x=-33740000;
#10;x=-33730000;
#10;x=-33720000;
#10;x=-33710000;
#10;x=-33700000;
#10;x=-33690000;
#10;x=-33680000;
#10;x=-33670000;
#10;x=-33660000;
#10;x=-33650000;
#10;x=-33640000;
#10;x=-33630000;
#10;x=-33620000;
#10;x=-33610000;
#10;x=-33600000;
#10;x=-33590000;
#10;x=-33580000;
#10;x=-33570000;
#10;x=-33560000;
#10;x=-33550000;
#10;x=-33540000;
#10;x=-33530000;
#10;x=-33520000;
#10;x=-33510000;
#10;x=-33500000;
#10;x=-33490000;
#10;x=-33480000;
#10;x=-33470000;
#10;x=-33460000;
#10;x=-33450000;
#10;x=-33440000;
#10;x=-33430000;
#10;x=-33420000;
#10;x=-33410000;
#10;x=-33400000;
#10;x=-33390000;
#10;x=-33380000;
#10;x=-33370000;
#10;x=-33360000;
#10;x=-33350000;
#10;x=-33340000;
#10;x=-33330000;
#10;x=-33320000;
#10;x=-33310000;
#10;x=-33300000;
#10;x=-33290000;
#10;x=-33280000;
#10;x=-33270000;
#10;x=-33260000;
#10;x=-33250000;
#10;x=-33240000;
#10;x=-33230000;
#10;x=-33220000;
#10;x=-33210000;
#10;x=-33200000;
#10;x=-33190000;
#10;x=-33180000;
#10;x=-33170000;
#10;x=-33160000;
#10;x=-33150000;
#10;x=-33140000;
#10;x=-33130000;
#10;x=-33120000;
#10;x=-33110000;
#10;x=-33100000;
#10;x=-33090000;
#10;x=-33080000;
#10;x=-33070000;
#10;x=-33060000;
#10;x=-33050000;
#10;x=-33040000;
#10;x=-33030000;
#10;x=-33020000;
#10;x=-33010000;
#10;x=-33000000;
#10;x=-32990000;
#10;x=-32980000;
#10;x=-32970000;
#10;x=-32960000;
#10;x=-32950000;
#10;x=-32940000;
#10;x=-32930000;
#10;x=-32920000;
#10;x=-32910000;
#10;x=-32900000;
#10;x=-32890000;
#10;x=-32880000;
#10;x=-32870000;
#10;x=-32860000;
#10;x=-32850000;
#10;x=-32840000;
#10;x=-32830000;
#10;x=-32820000;
#10;x=-32810000;
#10;x=-32800000;
#10;x=-32790000;
#10;x=-32780000;
#10;x=-32770000;
#10;x=-32760000;
#10;x=-32750000;
#10;x=-32740000;
#10;x=-32730000;
#10;x=-32720000;
#10;x=-32710000;
#10;x=-32700000;
#10;x=-32690000;
#10;x=-32680000;
#10;x=-32670000;
#10;x=-32660000;
#10;x=-32650000;
#10;x=-32640000;
#10;x=-32630000;
#10;x=-32620000;
#10;x=-32610000;
#10;x=-32600000;
#10;x=-32590000;
#10;x=-32580000;
#10;x=-32570000;
#10;x=-32560000;
#10;x=-32550000;
#10;x=-32540000;
#10;x=-32530000;
#10;x=-32520000;
#10;x=-32510000;
#10;x=-32500000;
#10;x=-32490000;
#10;x=-32480000;
#10;x=-32470000;
#10;x=-32460000;
#10;x=-32450000;
#10;x=-32440000;
#10;x=-32430000;
#10;x=-32420000;
#10;x=-32410000;
#10;x=-32400000;
#10;x=-32390000;
#10;x=-32380000;
#10;x=-32370000;
#10;x=-32360000;
#10;x=-32350000;
#10;x=-32340000;
#10;x=-32330000;
#10;x=-32320000;
#10;x=-32310000;
#10;x=-32300000;
#10;x=-32290000;
#10;x=-32280000;
#10;x=-32270000;
#10;x=-32260000;
#10;x=-32250000;
#10;x=-32240000;
#10;x=-32230000;
#10;x=-32220000;
#10;x=-32210000;
#10;x=-32200000;
#10;x=-32190000;
#10;x=-32180000;
#10;x=-32170000;
#10;x=-32160000;
#10;x=-32150000;
#10;x=-32140000;
#10;x=-32130000;
#10;x=-32120000;
#10;x=-32110000;
#10;x=-32100000;
#10;x=-32090000;
#10;x=-32080000;
#10;x=-32070000;
#10;x=-32060000;
#10;x=-32050000;
#10;x=-32040000;
#10;x=-32030000;
#10;x=-32020000;
#10;x=-32010000;
#10;x=-32000000;
#10;x=-31990000;
#10;x=-31980000;
#10;x=-31970000;
#10;x=-31960000;
#10;x=-31950000;
#10;x=-31940000;
#10;x=-31930000;
#10;x=-31920000;
#10;x=-31910000;
#10;x=-31900000;
#10;x=-31890000;
#10;x=-31880000;
#10;x=-31870000;
#10;x=-31860000;
#10;x=-31850000;
#10;x=-31840000;
#10;x=-31830000;
#10;x=-31820000;
#10;x=-31810000;
#10;x=-31800000;
#10;x=-31790000;
#10;x=-31780000;
#10;x=-31770000;
#10;x=-31760000;
#10;x=-31750000;
#10;x=-31740000;
#10;x=-31730000;
#10;x=-31720000;
#10;x=-31710000;
#10;x=-31700000;
#10;x=-31690000;
#10;x=-31680000;
#10;x=-31670000;
#10;x=-31660000;
#10;x=-31650000;
#10;x=-31640000;
#10;x=-31630000;
#10;x=-31620000;
#10;x=-31610000;
#10;x=-31600000;
#10;x=-31590000;
#10;x=-31580000;
#10;x=-31570000;
#10;x=-31560000;
#10;x=-31550000;
#10;x=-31540000;
#10;x=-31530000;
#10;x=-31520000;
#10;x=-31510000;
#10;x=-31500000;
#10;x=-31490000;
#10;x=-31480000;
#10;x=-31470000;
#10;x=-31460000;
#10;x=-31450000;
#10;x=-31440000;
#10;x=-31430000;
#10;x=-31420000;
#10;x=-31410000;
#10;x=-31400000;
#10;x=-31390000;
#10;x=-31380000;
#10;x=-31370000;
#10;x=-31360000;
#10;x=-31350000;
#10;x=-31340000;
#10;x=-31330000;
#10;x=-31320000;
#10;x=-31310000;
#10;x=-31300000;
#10;x=-31290000;
#10;x=-31280000;
#10;x=-31270000;
#10;x=-31260000;
#10;x=-31250000;
#10;x=-31240000;
#10;x=-31230000;
#10;x=-31220000;
#10;x=-31210000;
#10;x=-31200000;
#10;x=-31190000;
#10;x=-31180000;
#10;x=-31170000;
#10;x=-31160000;
#10;x=-31150000;
#10;x=-31140000;
#10;x=-31130000;
#10;x=-31120000;
#10;x=-31110000;
#10;x=-31100000;
#10;x=-31090000;
#10;x=-31080000;
#10;x=-31070000;
#10;x=-31060000;
#10;x=-31050000;
#10;x=-31040000;
#10;x=-31030000;
#10;x=-31020000;
#10;x=-31010000;
#10;x=-31000000;
#10;x=-30990000;
#10;x=-30980000;
#10;x=-30970000;
#10;x=-30960000;
#10;x=-30950000;
#10;x=-30940000;
#10;x=-30930000;
#10;x=-30920000;
#10;x=-30910000;
#10;x=-30900000;
#10;x=-30890000;
#10;x=-30880000;
#10;x=-30870000;
#10;x=-30860000;
#10;x=-30850000;
#10;x=-30840000;
#10;x=-30830000;
#10;x=-30820000;
#10;x=-30810000;
#10;x=-30800000;
#10;x=-30790000;
#10;x=-30780000;
#10;x=-30770000;
#10;x=-30760000;
#10;x=-30750000;
#10;x=-30740000;
#10;x=-30730000;
#10;x=-30720000;
#10;x=-30710000;
#10;x=-30700000;
#10;x=-30690000;
#10;x=-30680000;
#10;x=-30670000;
#10;x=-30660000;
#10;x=-30650000;
#10;x=-30640000;
#10;x=-30630000;
#10;x=-30620000;
#10;x=-30610000;
#10;x=-30600000;
#10;x=-30590000;
#10;x=-30580000;
#10;x=-30570000;
#10;x=-30560000;
#10;x=-30550000;
#10;x=-30540000;
#10;x=-30530000;
#10;x=-30520000;
#10;x=-30510000;
#10;x=-30500000;
#10;x=-30490000;
#10;x=-30480000;
#10;x=-30470000;
#10;x=-30460000;
#10;x=-30450000;
#10;x=-30440000;
#10;x=-30430000;
#10;x=-30420000;
#10;x=-30410000;
#10;x=-30400000;
#10;x=-30390000;
#10;x=-30380000;
#10;x=-30370000;
#10;x=-30360000;
#10;x=-30350000;
#10;x=-30340000;
#10;x=-30330000;
#10;x=-30320000;
#10;x=-30310000;
#10;x=-30300000;
#10;x=-30290000;
#10;x=-30280000;
#10;x=-30270000;
#10;x=-30260000;
#10;x=-30250000;
#10;x=-30240000;
#10;x=-30230000;
#10;x=-30220000;
#10;x=-30210000;
#10;x=-30200000;
#10;x=-30190000;
#10;x=-30180000;
#10;x=-30170000;
#10;x=-30160000;
#10;x=-30150000;
#10;x=-30140000;
#10;x=-30130000;
#10;x=-30120000;
#10;x=-30110000;
#10;x=-30100000;
#10;x=-30090000;
#10;x=-30080000;
#10;x=-30070000;
#10;x=-30060000;
#10;x=-30050000;
#10;x=-30040000;
#10;x=-30030000;
#10;x=-30020000;
#10;x=-30010000;
#10;x=-30000000;
#10;x=-29990000;
#10;x=-29980000;
#10;x=-29970000;
#10;x=-29960000;
#10;x=-29950000;
#10;x=-29940000;
#10;x=-29930000;
#10;x=-29920000;
#10;x=-29910000;
#10;x=-29900000;
#10;x=-29890000;
#10;x=-29880000;
#10;x=-29870000;
#10;x=-29860000;
#10;x=-29850000;
#10;x=-29840000;
#10;x=-29830000;
#10;x=-29820000;
#10;x=-29810000;
#10;x=-29800000;
#10;x=-29790000;
#10;x=-29780000;
#10;x=-29770000;
#10;x=-29760000;
#10;x=-29750000;
#10;x=-29740000;
#10;x=-29730000;
#10;x=-29720000;
#10;x=-29710000;
#10;x=-29700000;
#10;x=-29690000;
#10;x=-29680000;
#10;x=-29670000;
#10;x=-29660000;
#10;x=-29650000;
#10;x=-29640000;
#10;x=-29630000;
#10;x=-29620000;
#10;x=-29610000;
#10;x=-29600000;
#10;x=-29590000;
#10;x=-29580000;
#10;x=-29570000;
#10;x=-29560000;
#10;x=-29550000;
#10;x=-29540000;
#10;x=-29530000;
#10;x=-29520000;
#10;x=-29510000;
#10;x=-29500000;
#10;x=-29490000;
#10;x=-29480000;
#10;x=-29470000;
#10;x=-29460000;
#10;x=-29450000;
#10;x=-29440000;
#10;x=-29430000;
#10;x=-29420000;
#10;x=-29410000;
#10;x=-29400000;
#10;x=-29390000;
#10;x=-29380000;
#10;x=-29370000;
#10;x=-29360000;
#10;x=-29350000;
#10;x=-29340000;
#10;x=-29330000;
#10;x=-29320000;
#10;x=-29310000;
#10;x=-29300000;
#10;x=-29290000;
#10;x=-29280000;
#10;x=-29270000;
#10;x=-29260000;
#10;x=-29250000;
#10;x=-29240000;
#10;x=-29230000;
#10;x=-29220000;
#10;x=-29210000;
#10;x=-29200000;
#10;x=-29190000;
#10;x=-29180000;
#10;x=-29170000;
#10;x=-29160000;
#10;x=-29150000;
#10;x=-29140000;
#10;x=-29130000;
#10;x=-29120000;
#10;x=-29110000;
#10;x=-29100000;
#10;x=-29090000;
#10;x=-29080000;
#10;x=-29070000;
#10;x=-29060000;
#10;x=-29050000;
#10;x=-29040000;
#10;x=-29030000;
#10;x=-29020000;
#10;x=-29010000;
#10;x=-29000000;
#10;x=-28990000;
#10;x=-28980000;
#10;x=-28970000;
#10;x=-28960000;
#10;x=-28950000;
#10;x=-28940000;
#10;x=-28930000;
#10;x=-28920000;
#10;x=-28910000;
#10;x=-28900000;
#10;x=-28890000;
#10;x=-28880000;
#10;x=-28870000;
#10;x=-28860000;
#10;x=-28850000;
#10;x=-28840000;
#10;x=-28830000;
#10;x=-28820000;
#10;x=-28810000;
#10;x=-28800000;
#10;x=-28790000;
#10;x=-28780000;
#10;x=-28770000;
#10;x=-28760000;
#10;x=-28750000;
#10;x=-28740000;
#10;x=-28730000;
#10;x=-28720000;
#10;x=-28710000;
#10;x=-28700000;
#10;x=-28690000;
#10;x=-28680000;
#10;x=-28670000;
#10;x=-28660000;
#10;x=-28650000;
#10;x=-28640000;
#10;x=-28630000;
#10;x=-28620000;
#10;x=-28610000;
#10;x=-28600000;
#10;x=-28590000;
#10;x=-28580000;
#10;x=-28570000;
#10;x=-28560000;
#10;x=-28550000;
#10;x=-28540000;
#10;x=-28530000;
#10;x=-28520000;
#10;x=-28510000;
#10;x=-28500000;
#10;x=-28490000;
#10;x=-28480000;
#10;x=-28470000;
#10;x=-28460000;
#10;x=-28450000;
#10;x=-28440000;
#10;x=-28430000;
#10;x=-28420000;
#10;x=-28410000;
#10;x=-28400000;
#10;x=-28390000;
#10;x=-28380000;
#10;x=-28370000;
#10;x=-28360000;
#10;x=-28350000;
#10;x=-28340000;
#10;x=-28330000;
#10;x=-28320000;
#10;x=-28310000;
#10;x=-28300000;
#10;x=-28290000;
#10;x=-28280000;
#10;x=-28270000;
#10;x=-28260000;
#10;x=-28250000;
#10;x=-28240000;
#10;x=-28230000;
#10;x=-28220000;
#10;x=-28210000;
#10;x=-28200000;
#10;x=-28190000;
#10;x=-28180000;
#10;x=-28170000;
#10;x=-28160000;
#10;x=-28150000;
#10;x=-28140000;
#10;x=-28130000;
#10;x=-28120000;
#10;x=-28110000;
#10;x=-28100000;
#10;x=-28090000;
#10;x=-28080000;
#10;x=-28070000;
#10;x=-28060000;
#10;x=-28050000;
#10;x=-28040000;
#10;x=-28030000;
#10;x=-28020000;
#10;x=-28010000;
#10;x=-28000000;
#10;x=-27990000;
#10;x=-27980000;
#10;x=-27970000;
#10;x=-27960000;
#10;x=-27950000;
#10;x=-27940000;
#10;x=-27930000;
#10;x=-27920000;
#10;x=-27910000;
#10;x=-27900000;
#10;x=-27890000;
#10;x=-27880000;
#10;x=-27870000;
#10;x=-27860000;
#10;x=-27850000;
#10;x=-27840000;
#10;x=-27830000;
#10;x=-27820000;
#10;x=-27810000;
#10;x=-27800000;
#10;x=-27790000;
#10;x=-27780000;
#10;x=-27770000;
#10;x=-27760000;
#10;x=-27750000;
#10;x=-27740000;
#10;x=-27730000;
#10;x=-27720000;
#10;x=-27710000;
#10;x=-27700000;
#10;x=-27690000;
#10;x=-27680000;
#10;x=-27670000;
#10;x=-27660000;
#10;x=-27650000;
#10;x=-27640000;
#10;x=-27630000;
#10;x=-27620000;
#10;x=-27610000;
#10;x=-27600000;
#10;x=-27590000;
#10;x=-27580000;
#10;x=-27570000;
#10;x=-27560000;
#10;x=-27550000;
#10;x=-27540000;
#10;x=-27530000;
#10;x=-27520000;
#10;x=-27510000;
#10;x=-27500000;
#10;x=-27490000;
#10;x=-27480000;
#10;x=-27470000;
#10;x=-27460000;
#10;x=-27450000;
#10;x=-27440000;
#10;x=-27430000;
#10;x=-27420000;
#10;x=-27410000;
#10;x=-27400000;
#10;x=-27390000;
#10;x=-27380000;
#10;x=-27370000;
#10;x=-27360000;
#10;x=-27350000;
#10;x=-27340000;
#10;x=-27330000;
#10;x=-27320000;
#10;x=-27310000;
#10;x=-27300000;
#10;x=-27290000;
#10;x=-27280000;
#10;x=-27270000;
#10;x=-27260000;
#10;x=-27250000;
#10;x=-27240000;
#10;x=-27230000;
#10;x=-27220000;
#10;x=-27210000;
#10;x=-27200000;
#10;x=-27190000;
#10;x=-27180000;
#10;x=-27170000;
#10;x=-27160000;
#10;x=-27150000;
#10;x=-27140000;
#10;x=-27130000;
#10;x=-27120000;
#10;x=-27110000;
#10;x=-27100000;
#10;x=-27090000;
#10;x=-27080000;
#10;x=-27070000;
#10;x=-27060000;
#10;x=-27050000;
#10;x=-27040000;
#10;x=-27030000;
#10;x=-27020000;
#10;x=-27010000;
#10;x=-27000000;
#10;x=-26990000;
#10;x=-26980000;
#10;x=-26970000;
#10;x=-26960000;
#10;x=-26950000;
#10;x=-26940000;
#10;x=-26930000;
#10;x=-26920000;
#10;x=-26910000;
#10;x=-26900000;
#10;x=-26890000;
#10;x=-26880000;
#10;x=-26870000;
#10;x=-26860000;
#10;x=-26850000;
#10;x=-26840000;
#10;x=-26830000;
#10;x=-26820000;
#10;x=-26810000;
#10;x=-26800000;
#10;x=-26790000;
#10;x=-26780000;
#10;x=-26770000;
#10;x=-26760000;
#10;x=-26750000;
#10;x=-26740000;
#10;x=-26730000;
#10;x=-26720000;
#10;x=-26710000;
#10;x=-26700000;
#10;x=-26690000;
#10;x=-26680000;
#10;x=-26670000;
#10;x=-26660000;
#10;x=-26650000;
#10;x=-26640000;
#10;x=-26630000;
#10;x=-26620000;
#10;x=-26610000;
#10;x=-26600000;
#10;x=-26590000;
#10;x=-26580000;
#10;x=-26570000;
#10;x=-26560000;
#10;x=-26550000;
#10;x=-26540000;
#10;x=-26530000;
#10;x=-26520000;
#10;x=-26510000;
#10;x=-26500000;
#10;x=-26490000;
#10;x=-26480000;
#10;x=-26470000;
#10;x=-26460000;
#10;x=-26450000;
#10;x=-26440000;
#10;x=-26430000;
#10;x=-26420000;
#10;x=-26410000;
#10;x=-26400000;
#10;x=-26390000;
#10;x=-26380000;
#10;x=-26370000;
#10;x=-26360000;
#10;x=-26350000;
#10;x=-26340000;
#10;x=-26330000;
#10;x=-26320000;
#10;x=-26310000;
#10;x=-26300000;
#10;x=-26290000;
#10;x=-26280000;
#10;x=-26270000;
#10;x=-26260000;
#10;x=-26250000;
#10;x=-26240000;
#10;x=-26230000;
#10;x=-26220000;
#10;x=-26210000;
#10;x=-26200000;
#10;x=-26190000;
#10;x=-26180000;
#10;x=-26170000;
#10;x=-26160000;
#10;x=-26150000;
#10;x=-26140000;
#10;x=-26130000;
#10;x=-26120000;
#10;x=-26110000;
#10;x=-26100000;
#10;x=-26090000;
#10;x=-26080000;
#10;x=-26070000;
#10;x=-26060000;
#10;x=-26050000;
#10;x=-26040000;
#10;x=-26030000;
#10;x=-26020000;
#10;x=-26010000;
#10;x=-26000000;
#10;x=-25990000;
#10;x=-25980000;
#10;x=-25970000;
#10;x=-25960000;
#10;x=-25950000;
#10;x=-25940000;
#10;x=-25930000;
#10;x=-25920000;
#10;x=-25910000;
#10;x=-25900000;
#10;x=-25890000;
#10;x=-25880000;
#10;x=-25870000;
#10;x=-25860000;
#10;x=-25850000;
#10;x=-25840000;
#10;x=-25830000;
#10;x=-25820000;
#10;x=-25810000;
#10;x=-25800000;
#10;x=-25790000;
#10;x=-25780000;
#10;x=-25770000;
#10;x=-25760000;
#10;x=-25750000;
#10;x=-25740000;
#10;x=-25730000;
#10;x=-25720000;
#10;x=-25710000;
#10;x=-25700000;
#10;x=-25690000;
#10;x=-25680000;
#10;x=-25670000;
#10;x=-25660000;
#10;x=-25650000;
#10;x=-25640000;
#10;x=-25630000;
#10;x=-25620000;
#10;x=-25610000;
#10;x=-25600000;
#10;x=-25590000;
#10;x=-25580000;
#10;x=-25570000;
#10;x=-25560000;
#10;x=-25550000;
#10;x=-25540000;
#10;x=-25530000;
#10;x=-25520000;
#10;x=-25510000;
#10;x=-25500000;
#10;x=-25490000;
#10;x=-25480000;
#10;x=-25470000;
#10;x=-25460000;
#10;x=-25450000;
#10;x=-25440000;
#10;x=-25430000;
#10;x=-25420000;
#10;x=-25410000;
#10;x=-25400000;
#10;x=-25390000;
#10;x=-25380000;
#10;x=-25370000;
#10;x=-25360000;
#10;x=-25350000;
#10;x=-25340000;
#10;x=-25330000;
#10;x=-25320000;
#10;x=-25310000;
#10;x=-25300000;
#10;x=-25290000;
#10;x=-25280000;
#10;x=-25270000;
#10;x=-25260000;
#10;x=-25250000;
#10;x=-25240000;
#10;x=-25230000;
#10;x=-25220000;
#10;x=-25210000;
#10;x=-25200000;
#10;x=-25190000;
#10;x=-25180000;
#10;x=-25170000;
#10;x=-25160000;
#10;x=-25150000;
#10;x=-25140000;
#10;x=-25130000;
#10;x=-25120000;
#10;x=-25110000;
#10;x=-25100000;
#10;x=-25090000;
#10;x=-25080000;
#10;x=-25070000;
#10;x=-25060000;
#10;x=-25050000;
#10;x=-25040000;
#10;x=-25030000;
#10;x=-25020000;
#10;x=-25010000;
#10;x=-25000000;
#10;x=-24990000;
#10;x=-24980000;
#10;x=-24970000;
#10;x=-24960000;
#10;x=-24950000;
#10;x=-24940000;
#10;x=-24930000;
#10;x=-24920000;
#10;x=-24910000;
#10;x=-24900000;
#10;x=-24890000;
#10;x=-24880000;
#10;x=-24870000;
#10;x=-24860000;
#10;x=-24850000;
#10;x=-24840000;
#10;x=-24830000;
#10;x=-24820000;
#10;x=-24810000;
#10;x=-24800000;
#10;x=-24790000;
#10;x=-24780000;
#10;x=-24770000;
#10;x=-24760000;
#10;x=-24750000;
#10;x=-24740000;
#10;x=-24730000;
#10;x=-24720000;
#10;x=-24710000;
#10;x=-24700000;
#10;x=-24690000;
#10;x=-24680000;
#10;x=-24670000;
#10;x=-24660000;
#10;x=-24650000;
#10;x=-24640000;
#10;x=-24630000;
#10;x=-24620000;
#10;x=-24610000;
#10;x=-24600000;
#10;x=-24590000;
#10;x=-24580000;
#10;x=-24570000;
#10;x=-24560000;
#10;x=-24550000;
#10;x=-24540000;
#10;x=-24530000;
#10;x=-24520000;
#10;x=-24510000;
#10;x=-24500000;
#10;x=-24490000;
#10;x=-24480000;
#10;x=-24470000;
#10;x=-24460000;
#10;x=-24450000;
#10;x=-24440000;
#10;x=-24430000;
#10;x=-24420000;
#10;x=-24410000;
#10;x=-24400000;
#10;x=-24390000;
#10;x=-24380000;
#10;x=-24370000;
#10;x=-24360000;
#10;x=-24350000;
#10;x=-24340000;
#10;x=-24330000;
#10;x=-24320000;
#10;x=-24310000;
#10;x=-24300000;
#10;x=-24290000;
#10;x=-24280000;
#10;x=-24270000;
#10;x=-24260000;
#10;x=-24250000;
#10;x=-24240000;
#10;x=-24230000;
#10;x=-24220000;
#10;x=-24210000;
#10;x=-24200000;
#10;x=-24190000;
#10;x=-24180000;
#10;x=-24170000;
#10;x=-24160000;
#10;x=-24150000;
#10;x=-24140000;
#10;x=-24130000;
#10;x=-24120000;
#10;x=-24110000;
#10;x=-24100000;
#10;x=-24090000;
#10;x=-24080000;
#10;x=-24070000;
#10;x=-24060000;
#10;x=-24050000;
#10;x=-24040000;
#10;x=-24030000;
#10;x=-24020000;
#10;x=-24010000;
#10;x=-24000000;
#10;x=-23990000;
#10;x=-23980000;
#10;x=-23970000;
#10;x=-23960000;
#10;x=-23950000;
#10;x=-23940000;
#10;x=-23930000;
#10;x=-23920000;
#10;x=-23910000;
#10;x=-23900000;
#10;x=-23890000;
#10;x=-23880000;
#10;x=-23870000;
#10;x=-23860000;
#10;x=-23850000;
#10;x=-23840000;
#10;x=-23830000;
#10;x=-23820000;
#10;x=-23810000;
#10;x=-23800000;
#10;x=-23790000;
#10;x=-23780000;
#10;x=-23770000;
#10;x=-23760000;
#10;x=-23750000;
#10;x=-23740000;
#10;x=-23730000;
#10;x=-23720000;
#10;x=-23710000;
#10;x=-23700000;
#10;x=-23690000;
#10;x=-23680000;
#10;x=-23670000;
#10;x=-23660000;
#10;x=-23650000;
#10;x=-23640000;
#10;x=-23630000;
#10;x=-23620000;
#10;x=-23610000;
#10;x=-23600000;
#10;x=-23590000;
#10;x=-23580000;
#10;x=-23570000;
#10;x=-23560000;
#10;x=-23550000;
#10;x=-23540000;
#10;x=-23530000;
#10;x=-23520000;
#10;x=-23510000;
#10;x=-23500000;
#10;x=-23490000;
#10;x=-23480000;
#10;x=-23470000;
#10;x=-23460000;
#10;x=-23450000;
#10;x=-23440000;
#10;x=-23430000;
#10;x=-23420000;
#10;x=-23410000;
#10;x=-23400000;
#10;x=-23390000;
#10;x=-23380000;
#10;x=-23370000;
#10;x=-23360000;
#10;x=-23350000;
#10;x=-23340000;
#10;x=-23330000;
#10;x=-23320000;
#10;x=-23310000;
#10;x=-23300000;
#10;x=-23290000;
#10;x=-23280000;
#10;x=-23270000;
#10;x=-23260000;
#10;x=-23250000;
#10;x=-23240000;
#10;x=-23230000;
#10;x=-23220000;
#10;x=-23210000;
#10;x=-23200000;
#10;x=-23190000;
#10;x=-23180000;
#10;x=-23170000;
#10;x=-23160000;
#10;x=-23150000;
#10;x=-23140000;
#10;x=-23130000;
#10;x=-23120000;
#10;x=-23110000;
#10;x=-23100000;
#10;x=-23090000;
#10;x=-23080000;
#10;x=-23070000;
#10;x=-23060000;
#10;x=-23050000;
#10;x=-23040000;
#10;x=-23030000;
#10;x=-23020000;
#10;x=-23010000;
#10;x=-23000000;
#10;x=-22990000;
#10;x=-22980000;
#10;x=-22970000;
#10;x=-22960000;
#10;x=-22950000;
#10;x=-22940000;
#10;x=-22930000;
#10;x=-22920000;
#10;x=-22910000;
#10;x=-22900000;
#10;x=-22890000;
#10;x=-22880000;
#10;x=-22870000;
#10;x=-22860000;
#10;x=-22850000;
#10;x=-22840000;
#10;x=-22830000;
#10;x=-22820000;
#10;x=-22810000;
#10;x=-22800000;
#10;x=-22790000;
#10;x=-22780000;
#10;x=-22770000;
#10;x=-22760000;
#10;x=-22750000;
#10;x=-22740000;
#10;x=-22730000;
#10;x=-22720000;
#10;x=-22710000;
#10;x=-22700000;
#10;x=-22690000;
#10;x=-22680000;
#10;x=-22670000;
#10;x=-22660000;
#10;x=-22650000;
#10;x=-22640000;
#10;x=-22630000;
#10;x=-22620000;
#10;x=-22610000;
#10;x=-22600000;
#10;x=-22590000;
#10;x=-22580000;
#10;x=-22570000;
#10;x=-22560000;
#10;x=-22550000;
#10;x=-22540000;
#10;x=-22530000;
#10;x=-22520000;
#10;x=-22510000;
#10;x=-22500000;
#10;x=-22490000;
#10;x=-22480000;
#10;x=-22470000;
#10;x=-22460000;
#10;x=-22450000;
#10;x=-22440000;
#10;x=-22430000;
#10;x=-22420000;
#10;x=-22410000;
#10;x=-22400000;
#10;x=-22390000;
#10;x=-22380000;
#10;x=-22370000;
#10;x=-22360000;
#10;x=-22350000;
#10;x=-22340000;
#10;x=-22330000;
#10;x=-22320000;
#10;x=-22310000;
#10;x=-22300000;
#10;x=-22290000;
#10;x=-22280000;
#10;x=-22270000;
#10;x=-22260000;
#10;x=-22250000;
#10;x=-22240000;
#10;x=-22230000;
#10;x=-22220000;
#10;x=-22210000;
#10;x=-22200000;
#10;x=-22190000;
#10;x=-22180000;
#10;x=-22170000;
#10;x=-22160000;
#10;x=-22150000;
#10;x=-22140000;
#10;x=-22130000;
#10;x=-22120000;
#10;x=-22110000;
#10;x=-22100000;
#10;x=-22090000;
#10;x=-22080000;
#10;x=-22070000;
#10;x=-22060000;
#10;x=-22050000;
#10;x=-22040000;
#10;x=-22030000;
#10;x=-22020000;
#10;x=-22010000;
#10;x=-22000000;
#10;x=-21990000;
#10;x=-21980000;
#10;x=-21970000;
#10;x=-21960000;
#10;x=-21950000;
#10;x=-21940000;
#10;x=-21930000;
#10;x=-21920000;
#10;x=-21910000;
#10;x=-21900000;
#10;x=-21890000;
#10;x=-21880000;
#10;x=-21870000;
#10;x=-21860000;
#10;x=-21850000;
#10;x=-21840000;
#10;x=-21830000;
#10;x=-21820000;
#10;x=-21810000;
#10;x=-21800000;
#10;x=-21790000;
#10;x=-21780000;
#10;x=-21770000;
#10;x=-21760000;
#10;x=-21750000;
#10;x=-21740000;
#10;x=-21730000;
#10;x=-21720000;
#10;x=-21710000;
#10;x=-21700000;
#10;x=-21690000;
#10;x=-21680000;
#10;x=-21670000;
#10;x=-21660000;
#10;x=-21650000;
#10;x=-21640000;
#10;x=-21630000;
#10;x=-21620000;
#10;x=-21610000;
#10;x=-21600000;
#10;x=-21590000;
#10;x=-21580000;
#10;x=-21570000;
#10;x=-21560000;
#10;x=-21550000;
#10;x=-21540000;
#10;x=-21530000;
#10;x=-21520000;
#10;x=-21510000;
#10;x=-21500000;
#10;x=-21490000;
#10;x=-21480000;
#10;x=-21470000;
#10;x=-21460000;
#10;x=-21450000;
#10;x=-21440000;
#10;x=-21430000;
#10;x=-21420000;
#10;x=-21410000;
#10;x=-21400000;
#10;x=-21390000;
#10;x=-21380000;
#10;x=-21370000;
#10;x=-21360000;
#10;x=-21350000;
#10;x=-21340000;
#10;x=-21330000;
#10;x=-21320000;
#10;x=-21310000;
#10;x=-21300000;
#10;x=-21290000;
#10;x=-21280000;
#10;x=-21270000;
#10;x=-21260000;
#10;x=-21250000;
#10;x=-21240000;
#10;x=-21230000;
#10;x=-21220000;
#10;x=-21210000;
#10;x=-21200000;
#10;x=-21190000;
#10;x=-21180000;
#10;x=-21170000;
#10;x=-21160000;
#10;x=-21150000;
#10;x=-21140000;
#10;x=-21130000;
#10;x=-21120000;
#10;x=-21110000;
#10;x=-21100000;
#10;x=-21090000;
#10;x=-21080000;
#10;x=-21070000;
#10;x=-21060000;
#10;x=-21050000;
#10;x=-21040000;
#10;x=-21030000;
#10;x=-21020000;
#10;x=-21010000;
#10;x=-21000000;
#10;x=-20990000;
#10;x=-20980000;
#10;x=-20970000;
#10;x=-20960000;
#10;x=-20950000;
#10;x=-20940000;
#10;x=-20930000;
#10;x=-20920000;
#10;x=-20910000;
#10;x=-20900000;
#10;x=-20890000;
#10;x=-20880000;
#10;x=-20870000;
#10;x=-20860000;
#10;x=-20850000;
#10;x=-20840000;
#10;x=-20830000;
#10;x=-20820000;
#10;x=-20810000;
#10;x=-20800000;
#10;x=-20790000;
#10;x=-20780000;
#10;x=-20770000;
#10;x=-20760000;
#10;x=-20750000;
#10;x=-20740000;
#10;x=-20730000;
#10;x=-20720000;
#10;x=-20710000;
#10;x=-20700000;
#10;x=-20690000;
#10;x=-20680000;
#10;x=-20670000;
#10;x=-20660000;
#10;x=-20650000;
#10;x=-20640000;
#10;x=-20630000;
#10;x=-20620000;
#10;x=-20610000;
#10;x=-20600000;
#10;x=-20590000;
#10;x=-20580000;
#10;x=-20570000;
#10;x=-20560000;
#10;x=-20550000;
#10;x=-20540000;
#10;x=-20530000;
#10;x=-20520000;
#10;x=-20510000;
#10;x=-20500000;
#10;x=-20490000;
#10;x=-20480000;
#10;x=-20470000;
#10;x=-20460000;
#10;x=-20450000;
#10;x=-20440000;
#10;x=-20430000;
#10;x=-20420000;
#10;x=-20410000;
#10;x=-20400000;
#10;x=-20390000;
#10;x=-20380000;
#10;x=-20370000;
#10;x=-20360000;
#10;x=-20350000;
#10;x=-20340000;
#10;x=-20330000;
#10;x=-20320000;
#10;x=-20310000;
#10;x=-20300000;
#10;x=-20290000;
#10;x=-20280000;
#10;x=-20270000;
#10;x=-20260000;
#10;x=-20250000;
#10;x=-20240000;
#10;x=-20230000;
#10;x=-20220000;
#10;x=-20210000;
#10;x=-20200000;
#10;x=-20190000;
#10;x=-20180000;
#10;x=-20170000;
#10;x=-20160000;
#10;x=-20150000;
#10;x=-20140000;
#10;x=-20130000;
#10;x=-20120000;
#10;x=-20110000;
#10;x=-20100000;
#10;x=-20090000;
#10;x=-20080000;
#10;x=-20070000;
#10;x=-20060000;
#10;x=-20050000;
#10;x=-20040000;
#10;x=-20030000;
#10;x=-20020000;
#10;x=-20010000;
#10;x=-20000000;
#10;x=-19990000;
#10;x=-19980000;
#10;x=-19970000;
#10;x=-19960000;
#10;x=-19950000;
#10;x=-19940000;
#10;x=-19930000;
#10;x=-19920000;
#10;x=-19910000;
#10;x=-19900000;
#10;x=-19890000;
#10;x=-19880000;
#10;x=-19870000;
#10;x=-19860000;
#10;x=-19850000;
#10;x=-19840000;
#10;x=-19830000;
#10;x=-19820000;
#10;x=-19810000;
#10;x=-19800000;
#10;x=-19790000;
#10;x=-19780000;
#10;x=-19770000;
#10;x=-19760000;
#10;x=-19750000;
#10;x=-19740000;
#10;x=-19730000;
#10;x=-19720000;
#10;x=-19710000;
#10;x=-19700000;
#10;x=-19690000;
#10;x=-19680000;
#10;x=-19670000;
#10;x=-19660000;
#10;x=-19650000;
#10;x=-19640000;
#10;x=-19630000;
#10;x=-19620000;
#10;x=-19610000;
#10;x=-19600000;
#10;x=-19590000;
#10;x=-19580000;
#10;x=-19570000;
#10;x=-19560000;
#10;x=-19550000;
#10;x=-19540000;
#10;x=-19530000;
#10;x=-19520000;
#10;x=-19510000;
#10;x=-19500000;
#10;x=-19490000;
#10;x=-19480000;
#10;x=-19470000;
#10;x=-19460000;
#10;x=-19450000;
#10;x=-19440000;
#10;x=-19430000;
#10;x=-19420000;
#10;x=-19410000;
#10;x=-19400000;
#10;x=-19390000;
#10;x=-19380000;
#10;x=-19370000;
#10;x=-19360000;
#10;x=-19350000;
#10;x=-19340000;
#10;x=-19330000;
#10;x=-19320000;
#10;x=-19310000;
#10;x=-19300000;
#10;x=-19290000;
#10;x=-19280000;
#10;x=-19270000;
#10;x=-19260000;
#10;x=-19250000;
#10;x=-19240000;
#10;x=-19230000;
#10;x=-19220000;
#10;x=-19210000;
#10;x=-19200000;
#10;x=-19190000;
#10;x=-19180000;
#10;x=-19170000;
#10;x=-19160000;
#10;x=-19150000;
#10;x=-19140000;
#10;x=-19130000;
#10;x=-19120000;
#10;x=-19110000;
#10;x=-19100000;
#10;x=-19090000;
#10;x=-19080000;
#10;x=-19070000;
#10;x=-19060000;
#10;x=-19050000;
#10;x=-19040000;
#10;x=-19030000;
#10;x=-19020000;
#10;x=-19010000;
#10;x=-19000000;
#10;x=-18990000;
#10;x=-18980000;
#10;x=-18970000;
#10;x=-18960000;
#10;x=-18950000;
#10;x=-18940000;
#10;x=-18930000;
#10;x=-18920000;
#10;x=-18910000;
#10;x=-18900000;
#10;x=-18890000;
#10;x=-18880000;
#10;x=-18870000;
#10;x=-18860000;
#10;x=-18850000;
#10;x=-18840000;
#10;x=-18830000;
#10;x=-18820000;
#10;x=-18810000;
#10;x=-18800000;
#10;x=-18790000;
#10;x=-18780000;
#10;x=-18770000;
#10;x=-18760000;
#10;x=-18750000;
#10;x=-18740000;
#10;x=-18730000;
#10;x=-18720000;
#10;x=-18710000;
#10;x=-18700000;
#10;x=-18690000;
#10;x=-18680000;
#10;x=-18670000;
#10;x=-18660000;
#10;x=-18650000;
#10;x=-18640000;
#10;x=-18630000;
#10;x=-18620000;
#10;x=-18610000;
#10;x=-18600000;
#10;x=-18590000;
#10;x=-18580000;
#10;x=-18570000;
#10;x=-18560000;
#10;x=-18550000;
#10;x=-18540000;
#10;x=-18530000;
#10;x=-18520000;
#10;x=-18510000;
#10;x=-18500000;
#10;x=-18490000;
#10;x=-18480000;
#10;x=-18470000;
#10;x=-18460000;
#10;x=-18450000;
#10;x=-18440000;
#10;x=-18430000;
#10;x=-18420000;
#10;x=-18410000;
#10;x=-18400000;
#10;x=-18390000;
#10;x=-18380000;
#10;x=-18370000;
#10;x=-18360000;
#10;x=-18350000;
#10;x=-18340000;
#10;x=-18330000;
#10;x=-18320000;
#10;x=-18310000;
#10;x=-18300000;
#10;x=-18290000;
#10;x=-18280000;
#10;x=-18270000;
#10;x=-18260000;
#10;x=-18250000;
#10;x=-18240000;
#10;x=-18230000;
#10;x=-18220000;
#10;x=-18210000;
#10;x=-18200000;
#10;x=-18190000;
#10;x=-18180000;
#10;x=-18170000;
#10;x=-18160000;
#10;x=-18150000;
#10;x=-18140000;
#10;x=-18130000;
#10;x=-18120000;
#10;x=-18110000;
#10;x=-18100000;
#10;x=-18090000;
#10;x=-18080000;
#10;x=-18070000;
#10;x=-18060000;
#10;x=-18050000;
#10;x=-18040000;
#10;x=-18030000;
#10;x=-18020000;
#10;x=-18010000;
#10;x=-18000000;
#10;x=-17990000;
#10;x=-17980000;
#10;x=-17970000;
#10;x=-17960000;
#10;x=-17950000;
#10;x=-17940000;
#10;x=-17930000;
#10;x=-17920000;
#10;x=-17910000;
#10;x=-17900000;
#10;x=-17890000;
#10;x=-17880000;
#10;x=-17870000;
#10;x=-17860000;
#10;x=-17850000;
#10;x=-17840000;
#10;x=-17830000;
#10;x=-17820000;
#10;x=-17810000;
#10;x=-17800000;
#10;x=-17790000;
#10;x=-17780000;
#10;x=-17770000;
#10;x=-17760000;
#10;x=-17750000;
#10;x=-17740000;
#10;x=-17730000;
#10;x=-17720000;
#10;x=-17710000;
#10;x=-17700000;
#10;x=-17690000;
#10;x=-17680000;
#10;x=-17670000;
#10;x=-17660000;
#10;x=-17650000;
#10;x=-17640000;
#10;x=-17630000;
#10;x=-17620000;
#10;x=-17610000;
#10;x=-17600000;
#10;x=-17590000;
#10;x=-17580000;
#10;x=-17570000;
#10;x=-17560000;
#10;x=-17550000;
#10;x=-17540000;
#10;x=-17530000;
#10;x=-17520000;
#10;x=-17510000;
#10;x=-17500000;
#10;x=-17490000;
#10;x=-17480000;
#10;x=-17470000;
#10;x=-17460000;
#10;x=-17450000;
#10;x=-17440000;
#10;x=-17430000;
#10;x=-17420000;
#10;x=-17410000;
#10;x=-17400000;
#10;x=-17390000;
#10;x=-17380000;
#10;x=-17370000;
#10;x=-17360000;
#10;x=-17350000;
#10;x=-17340000;
#10;x=-17330000;
#10;x=-17320000;
#10;x=-17310000;
#10;x=-17300000;
#10;x=-17290000;
#10;x=-17280000;
#10;x=-17270000;
#10;x=-17260000;
#10;x=-17250000;
#10;x=-17240000;
#10;x=-17230000;
#10;x=-17220000;
#10;x=-17210000;
#10;x=-17200000;
#10;x=-17190000;
#10;x=-17180000;
#10;x=-17170000;
#10;x=-17160000;
#10;x=-17150000;
#10;x=-17140000;
#10;x=-17130000;
#10;x=-17120000;
#10;x=-17110000;
#10;x=-17100000;
#10;x=-17090000;
#10;x=-17080000;
#10;x=-17070000;
#10;x=-17060000;
#10;x=-17050000;
#10;x=-17040000;
#10;x=-17030000;
#10;x=-17020000;
#10;x=-17010000;
#10;x=-17000000;
#10;x=-16990000;
#10;x=-16980000;
#10;x=-16970000;
#10;x=-16960000;
#10;x=-16950000;
#10;x=-16940000;
#10;x=-16930000;
#10;x=-16920000;
#10;x=-16910000;
#10;x=-16900000;
#10;x=-16890000;
#10;x=-16880000;
#10;x=-16870000;
#10;x=-16860000;
#10;x=-16850000;
#10;x=-16840000;
#10;x=-16830000;
#10;x=-16820000;
#10;x=-16810000;
#10;x=-16800000;
#10;x=-16790000;
#10;x=-16780000;
#10;x=-16770000;
#10;x=-16760000;
#10;x=-16750000;
#10;x=-16740000;
#10;x=-16730000;
#10;x=-16720000;
#10;x=-16710000;
#10;x=-16700000;
#10;x=-16690000;
#10;x=-16680000;
#10;x=-16670000;
#10;x=-16660000;
#10;x=-16650000;
#10;x=-16640000;
#10;x=-16630000;
#10;x=-16620000;
#10;x=-16610000;
#10;x=-16600000;
#10;x=-16590000;
#10;x=-16580000;
#10;x=-16570000;
#10;x=-16560000;
#10;x=-16550000;
#10;x=-16540000;
#10;x=-16530000;
#10;x=-16520000;
#10;x=-16510000;
#10;x=-16500000;
#10;x=-16490000;
#10;x=-16480000;
#10;x=-16470000;
#10;x=-16460000;
#10;x=-16450000;
#10;x=-16440000;
#10;x=-16430000;
#10;x=-16420000;
#10;x=-16410000;
#10;x=-16400000;
#10;x=-16390000;
#10;x=-16380000;
#10;x=-16370000;
#10;x=-16360000;
#10;x=-16350000;
#10;x=-16340000;
#10;x=-16330000;
#10;x=-16320000;
#10;x=-16310000;
#10;x=-16300000;
#10;x=-16290000;
#10;x=-16280000;
#10;x=-16270000;
#10;x=-16260000;
#10;x=-16250000;
#10;x=-16240000;
#10;x=-16230000;
#10;x=-16220000;
#10;x=-16210000;
#10;x=-16200000;
#10;x=-16190000;
#10;x=-16180000;
#10;x=-16170000;
#10;x=-16160000;
#10;x=-16150000;
#10;x=-16140000;
#10;x=-16130000;
#10;x=-16120000;
#10;x=-16110000;
#10;x=-16100000;
#10;x=-16090000;
#10;x=-16080000;
#10;x=-16070000;
#10;x=-16060000;
#10;x=-16050000;
#10;x=-16040000;
#10;x=-16030000;
#10;x=-16020000;
#10;x=-16010000;
#10;x=-16000000;
#10;x=-15990000;
#10;x=-15980000;
#10;x=-15970000;
#10;x=-15960000;
#10;x=-15950000;
#10;x=-15940000;
#10;x=-15930000;
#10;x=-15920000;
#10;x=-15910000;
#10;x=-15900000;
#10;x=-15890000;
#10;x=-15880000;
#10;x=-15870000;
#10;x=-15860000;
#10;x=-15850000;
#10;x=-15840000;
#10;x=-15830000;
#10;x=-15820000;
#10;x=-15810000;
#10;x=-15800000;
#10;x=-15790000;
#10;x=-15780000;
#10;x=-15770000;
#10;x=-15760000;
#10;x=-15750000;
#10;x=-15740000;
#10;x=-15730000;
#10;x=-15720000;
#10;x=-15710000;
#10;x=-15700000;
#10;x=-15690000;
#10;x=-15680000;
#10;x=-15670000;
#10;x=-15660000;
#10;x=-15650000;
#10;x=-15640000;
#10;x=-15630000;
#10;x=-15620000;
#10;x=-15610000;
#10;x=-15600000;
#10;x=-15590000;
#10;x=-15580000;
#10;x=-15570000;
#10;x=-15560000;
#10;x=-15550000;
#10;x=-15540000;
#10;x=-15530000;
#10;x=-15520000;
#10;x=-15510000;
#10;x=-15500000;
#10;x=-15490000;
#10;x=-15480000;
#10;x=-15470000;
#10;x=-15460000;
#10;x=-15450000;
#10;x=-15440000;
#10;x=-15430000;
#10;x=-15420000;
#10;x=-15410000;
#10;x=-15400000;
#10;x=-15390000;
#10;x=-15380000;
#10;x=-15370000;
#10;x=-15360000;
#10;x=-15350000;
#10;x=-15340000;
#10;x=-15330000;
#10;x=-15320000;
#10;x=-15310000;
#10;x=-15300000;
#10;x=-15290000;
#10;x=-15280000;
#10;x=-15270000;
#10;x=-15260000;
#10;x=-15250000;
#10;x=-15240000;
#10;x=-15230000;
#10;x=-15220000;
#10;x=-15210000;
#10;x=-15200000;
#10;x=-15190000;
#10;x=-15180000;
#10;x=-15170000;
#10;x=-15160000;
#10;x=-15150000;
#10;x=-15140000;
#10;x=-15130000;
#10;x=-15120000;
#10;x=-15110000;
#10;x=-15100000;
#10;x=-15090000;
#10;x=-15080000;
#10;x=-15070000;
#10;x=-15060000;
#10;x=-15050000;
#10;x=-15040000;
#10;x=-15030000;
#10;x=-15020000;
#10;x=-15010000;
#10;x=-15000000;
#10;x=-14990000;
#10;x=-14980000;
#10;x=-14970000;
#10;x=-14960000;
#10;x=-14950000;
#10;x=-14940000;
#10;x=-14930000;
#10;x=-14920000;
#10;x=-14910000;
#10;x=-14900000;
#10;x=-14890000;
#10;x=-14880000;
#10;x=-14870000;
#10;x=-14860000;
#10;x=-14850000;
#10;x=-14840000;
#10;x=-14830000;
#10;x=-14820000;
#10;x=-14810000;
#10;x=-14800000;
#10;x=-14790000;
#10;x=-14780000;
#10;x=-14770000;
#10;x=-14760000;
#10;x=-14750000;
#10;x=-14740000;
#10;x=-14730000;
#10;x=-14720000;
#10;x=-14710000;
#10;x=-14700000;
#10;x=-14690000;
#10;x=-14680000;
#10;x=-14670000;
#10;x=-14660000;
#10;x=-14650000;
#10;x=-14640000;
#10;x=-14630000;
#10;x=-14620000;
#10;x=-14610000;
#10;x=-14600000;
#10;x=-14590000;
#10;x=-14580000;
#10;x=-14570000;
#10;x=-14560000;
#10;x=-14550000;
#10;x=-14540000;
#10;x=-14530000;
#10;x=-14520000;
#10;x=-14510000;
#10;x=-14500000;
#10;x=-14490000;
#10;x=-14480000;
#10;x=-14470000;
#10;x=-14460000;
#10;x=-14450000;
#10;x=-14440000;
#10;x=-14430000;
#10;x=-14420000;
#10;x=-14410000;
#10;x=-14400000;
#10;x=-14390000;
#10;x=-14380000;
#10;x=-14370000;
#10;x=-14360000;
#10;x=-14350000;
#10;x=-14340000;
#10;x=-14330000;
#10;x=-14320000;
#10;x=-14310000;
#10;x=-14300000;
#10;x=-14290000;
#10;x=-14280000;
#10;x=-14270000;
#10;x=-14260000;
#10;x=-14250000;
#10;x=-14240000;
#10;x=-14230000;
#10;x=-14220000;
#10;x=-14210000;
#10;x=-14200000;
#10;x=-14190000;
#10;x=-14180000;
#10;x=-14170000;
#10;x=-14160000;
#10;x=-14150000;
#10;x=-14140000;
#10;x=-14130000;
#10;x=-14120000;
#10;x=-14110000;
#10;x=-14100000;
#10;x=-14090000;
#10;x=-14080000;
#10;x=-14070000;
#10;x=-14060000;
#10;x=-14050000;
#10;x=-14040000;
#10;x=-14030000;
#10;x=-14020000;
#10;x=-14010000;
#10;x=-14000000;
#10;x=-13990000;
#10;x=-13980000;
#10;x=-13970000;
#10;x=-13960000;
#10;x=-13950000;
#10;x=-13940000;
#10;x=-13930000;
#10;x=-13920000;
#10;x=-13910000;
#10;x=-13900000;
#10;x=-13890000;
#10;x=-13880000;
#10;x=-13870000;
#10;x=-13860000;
#10;x=-13850000;
#10;x=-13840000;
#10;x=-13830000;
#10;x=-13820000;
#10;x=-13810000;
#10;x=-13800000;
#10;x=-13790000;
#10;x=-13780000;
#10;x=-13770000;
#10;x=-13760000;
#10;x=-13750000;
#10;x=-13740000;
#10;x=-13730000;
#10;x=-13720000;
#10;x=-13710000;
#10;x=-13700000;
#10;x=-13690000;
#10;x=-13680000;
#10;x=-13670000;
#10;x=-13660000;
#10;x=-13650000;
#10;x=-13640000;
#10;x=-13630000;
#10;x=-13620000;
#10;x=-13610000;
#10;x=-13600000;
#10;x=-13590000;
#10;x=-13580000;
#10;x=-13570000;
#10;x=-13560000;
#10;x=-13550000;
#10;x=-13540000;
#10;x=-13530000;
#10;x=-13520000;
#10;x=-13510000;
#10;x=-13500000;
#10;x=-13490000;
#10;x=-13480000;
#10;x=-13470000;
#10;x=-13460000;
#10;x=-13450000;
#10;x=-13440000;
#10;x=-13430000;
#10;x=-13420000;
#10;x=-13410000;
#10;x=-13400000;
#10;x=-13390000;
#10;x=-13380000;
#10;x=-13370000;
#10;x=-13360000;
#10;x=-13350000;
#10;x=-13340000;
#10;x=-13330000;
#10;x=-13320000;
#10;x=-13310000;
#10;x=-13300000;
#10;x=-13290000;
#10;x=-13280000;
#10;x=-13270000;
#10;x=-13260000;
#10;x=-13250000;
#10;x=-13240000;
#10;x=-13230000;
#10;x=-13220000;
#10;x=-13210000;
#10;x=-13200000;
#10;x=-13190000;
#10;x=-13180000;
#10;x=-13170000;
#10;x=-13160000;
#10;x=-13150000;
#10;x=-13140000;
#10;x=-13130000;
#10;x=-13120000;
#10;x=-13110000;
#10;x=-13100000;
#10;x=-13090000;
#10;x=-13080000;
#10;x=-13070000;
#10;x=-13060000;
#10;x=-13050000;
#10;x=-13040000;
#10;x=-13030000;
#10;x=-13020000;
#10;x=-13010000;
#10;x=-13000000;
#10;x=-12990000;
#10;x=-12980000;
#10;x=-12970000;
#10;x=-12960000;
#10;x=-12950000;
#10;x=-12940000;
#10;x=-12930000;
#10;x=-12920000;
#10;x=-12910000;
#10;x=-12900000;
#10;x=-12890000;
#10;x=-12880000;
#10;x=-12870000;
#10;x=-12860000;
#10;x=-12850000;
#10;x=-12840000;
#10;x=-12830000;
#10;x=-12820000;
#10;x=-12810000;
#10;x=-12800000;
#10;x=-12790000;
#10;x=-12780000;
#10;x=-12770000;
#10;x=-12760000;
#10;x=-12750000;
#10;x=-12740000;
#10;x=-12730000;
#10;x=-12720000;
#10;x=-12710000;
#10;x=-12700000;
#10;x=-12690000;
#10;x=-12680000;
#10;x=-12670000;
#10;x=-12660000;
#10;x=-12650000;
#10;x=-12640000;
#10;x=-12630000;
#10;x=-12620000;
#10;x=-12610000;
#10;x=-12600000;
#10;x=-12590000;
#10;x=-12580000;
#10;x=-12570000;
#10;x=-12560000;
#10;x=-12550000;
#10;x=-12540000;
#10;x=-12530000;
#10;x=-12520000;
#10;x=-12510000;
#10;x=-12500000;
#10;x=-12490000;
#10;x=-12480000;
#10;x=-12470000;
#10;x=-12460000;
#10;x=-12450000;
#10;x=-12440000;
#10;x=-12430000;
#10;x=-12420000;
#10;x=-12410000;
#10;x=-12400000;
#10;x=-12390000;
#10;x=-12380000;
#10;x=-12370000;
#10;x=-12360000;
#10;x=-12350000;
#10;x=-12340000;
#10;x=-12330000;
#10;x=-12320000;
#10;x=-12310000;
#10;x=-12300000;
#10;x=-12290000;
#10;x=-12280000;
#10;x=-12270000;
#10;x=-12260000;
#10;x=-12250000;
#10;x=-12240000;
#10;x=-12230000;
#10;x=-12220000;
#10;x=-12210000;
#10;x=-12200000;
#10;x=-12190000;
#10;x=-12180000;
#10;x=-12170000;
#10;x=-12160000;
#10;x=-12150000;
#10;x=-12140000;
#10;x=-12130000;
#10;x=-12120000;
#10;x=-12110000;
#10;x=-12100000;
#10;x=-12090000;
#10;x=-12080000;
#10;x=-12070000;
#10;x=-12060000;
#10;x=-12050000;
#10;x=-12040000;
#10;x=-12030000;
#10;x=-12020000;
#10;x=-12010000;
#10;x=-12000000;
#10;x=-11990000;
#10;x=-11980000;
#10;x=-11970000;
#10;x=-11960000;
#10;x=-11950000;
#10;x=-11940000;
#10;x=-11930000;
#10;x=-11920000;
#10;x=-11910000;
#10;x=-11900000;
#10;x=-11890000;
#10;x=-11880000;
#10;x=-11870000;
#10;x=-11860000;
#10;x=-11850000;
#10;x=-11840000;
#10;x=-11830000;
#10;x=-11820000;
#10;x=-11810000;
#10;x=-11800000;
#10;x=-11790000;
#10;x=-11780000;
#10;x=-11770000;
#10;x=-11760000;
#10;x=-11750000;
#10;x=-11740000;
#10;x=-11730000;
#10;x=-11720000;
#10;x=-11710000;
#10;x=-11700000;
#10;x=-11690000;
#10;x=-11680000;
#10;x=-11670000;
#10;x=-11660000;
#10;x=-11650000;
#10;x=-11640000;
#10;x=-11630000;
#10;x=-11620000;
#10;x=-11610000;
#10;x=-11600000;
#10;x=-11590000;
#10;x=-11580000;
#10;x=-11570000;
#10;x=-11560000;
#10;x=-11550000;
#10;x=-11540000;
#10;x=-11530000;
#10;x=-11520000;
#10;x=-11510000;
#10;x=-11500000;
#10;x=-11490000;
#10;x=-11480000;
#10;x=-11470000;
#10;x=-11460000;
#10;x=-11450000;
#10;x=-11440000;
#10;x=-11430000;
#10;x=-11420000;
#10;x=-11410000;
#10;x=-11400000;
#10;x=-11390000;
#10;x=-11380000;
#10;x=-11370000;
#10;x=-11360000;
#10;x=-11350000;
#10;x=-11340000;
#10;x=-11330000;
#10;x=-11320000;
#10;x=-11310000;
#10;x=-11300000;
#10;x=-11290000;
#10;x=-11280000;
#10;x=-11270000;
#10;x=-11260000;
#10;x=-11250000;
#10;x=-11240000;
#10;x=-11230000;
#10;x=-11220000;
#10;x=-11210000;
#10;x=-11200000;
#10;x=-11190000;
#10;x=-11180000;
#10;x=-11170000;
#10;x=-11160000;
#10;x=-11150000;
#10;x=-11140000;
#10;x=-11130000;
#10;x=-11120000;
#10;x=-11110000;
#10;x=-11100000;
#10;x=-11090000;
#10;x=-11080000;
#10;x=-11070000;
#10;x=-11060000;
#10;x=-11050000;
#10;x=-11040000;
#10;x=-11030000;
#10;x=-11020000;
#10;x=-11010000;
#10;x=-11000000;
#10;x=-10990000;
#10;x=-10980000;
#10;x=-10970000;
#10;x=-10960000;
#10;x=-10950000;
#10;x=-10940000;
#10;x=-10930000;
#10;x=-10920000;
#10;x=-10910000;
#10;x=-10900000;
#10;x=-10890000;
#10;x=-10880000;
#10;x=-10870000;
#10;x=-10860000;
#10;x=-10850000;
#10;x=-10840000;
#10;x=-10830000;
#10;x=-10820000;
#10;x=-10810000;
#10;x=-10800000;
#10;x=-10790000;
#10;x=-10780000;
#10;x=-10770000;
#10;x=-10760000;
#10;x=-10750000;
#10;x=-10740000;
#10;x=-10730000;
#10;x=-10720000;
#10;x=-10710000;
#10;x=-10700000;
#10;x=-10690000;
#10;x=-10680000;
#10;x=-10670000;
#10;x=-10660000;
#10;x=-10650000;
#10;x=-10640000;
#10;x=-10630000;
#10;x=-10620000;
#10;x=-10610000;
#10;x=-10600000;
#10;x=-10590000;
#10;x=-10580000;
#10;x=-10570000;
#10;x=-10560000;
#10;x=-10550000;
#10;x=-10540000;
#10;x=-10530000;
#10;x=-10520000;
#10;x=-10510000;
#10;x=-10500000;
#10;x=-10490000;
#10;x=-10480000;
#10;x=-10470000;
#10;x=-10460000;
#10;x=-10450000;
#10;x=-10440000;
#10;x=-10430000;
#10;x=-10420000;
#10;x=-10410000;
#10;x=-10400000;
#10;x=-10390000;
#10;x=-10380000;
#10;x=-10370000;
#10;x=-10360000;
#10;x=-10350000;
#10;x=-10340000;
#10;x=-10330000;
#10;x=-10320000;
#10;x=-10310000;
#10;x=-10300000;
#10;x=-10290000;
#10;x=-10280000;
#10;x=-10270000;
#10;x=-10260000;
#10;x=-10250000;
#10;x=-10240000;
#10;x=-10230000;
#10;x=-10220000;
#10;x=-10210000;
#10;x=-10200000;
#10;x=-10190000;
#10;x=-10180000;
#10;x=-10170000;
#10;x=-10160000;
#10;x=-10150000;
#10;x=-10140000;
#10;x=-10130000;
#10;x=-10120000;
#10;x=-10110000;
#10;x=-10100000;
#10;x=-10090000;
#10;x=-10080000;
#10;x=-10070000;
#10;x=-10060000;
#10;x=-10050000;
#10;x=-10040000;
#10;x=-10030000;
#10;x=-10020000;
#10;x=-10010000;
#10;x=-10000000;
#10;x=-9990000;
#10;x=-9980000;
#10;x=-9970000;
#10;x=-9960000;
#10;x=-9950000;
#10;x=-9940000;
#10;x=-9930000;
#10;x=-9920000;
#10;x=-9910000;
#10;x=-9900000;
#10;x=-9890000;
#10;x=-9880000;
#10;x=-9870000;
#10;x=-9860000;
#10;x=-9850000;
#10;x=-9840000;
#10;x=-9830000;
#10;x=-9820000;
#10;x=-9810000;
#10;x=-9800000;
#10;x=-9790000;
#10;x=-9780000;
#10;x=-9770000;
#10;x=-9760000;
#10;x=-9750000;
#10;x=-9740000;
#10;x=-9730000;
#10;x=-9720000;
#10;x=-9710000;
#10;x=-9700000;
#10;x=-9690000;
#10;x=-9680000;
#10;x=-9670000;
#10;x=-9660000;
#10;x=-9650000;
#10;x=-9640000;
#10;x=-9630000;
#10;x=-9620000;
#10;x=-9610000;
#10;x=-9600000;
#10;x=-9590000;
#10;x=-9580000;
#10;x=-9570000;
#10;x=-9560000;
#10;x=-9550000;
#10;x=-9540000;
#10;x=-9530000;
#10;x=-9520000;
#10;x=-9510000;
#10;x=-9500000;
#10;x=-9490000;
#10;x=-9480000;
#10;x=-9470000;
#10;x=-9460000;
#10;x=-9450000;
#10;x=-9440000;
#10;x=-9430000;
#10;x=-9420000;
#10;x=-9410000;
#10;x=-9400000;
#10;x=-9390000;
#10;x=-9380000;
#10;x=-9370000;
#10;x=-9360000;
#10;x=-9350000;
#10;x=-9340000;
#10;x=-9330000;
#10;x=-9320000;
#10;x=-9310000;
#10;x=-9300000;
#10;x=-9290000;
#10;x=-9280000;
#10;x=-9270000;
#10;x=-9260000;
#10;x=-9250000;
#10;x=-9240000;
#10;x=-9230000;
#10;x=-9220000;
#10;x=-9210000;
#10;x=-9200000;
#10;x=-9190000;
#10;x=-9180000;
#10;x=-9170000;
#10;x=-9160000;
#10;x=-9150000;
#10;x=-9140000;
#10;x=-9130000;
#10;x=-9120000;
#10;x=-9110000;
#10;x=-9100000;
#10;x=-9090000;
#10;x=-9080000;
#10;x=-9070000;
#10;x=-9060000;
#10;x=-9050000;
#10;x=-9040000;
#10;x=-9030000;
#10;x=-9020000;
#10;x=-9010000;
#10;x=-9000000;
#10;x=-8990000;
#10;x=-8980000;
#10;x=-8970000;
#10;x=-8960000;
#10;x=-8950000;
#10;x=-8940000;
#10;x=-8930000;
#10;x=-8920000;
#10;x=-8910000;
#10;x=-8900000;
#10;x=-8890000;
#10;x=-8880000;
#10;x=-8870000;
#10;x=-8860000;
#10;x=-8850000;
#10;x=-8840000;
#10;x=-8830000;
#10;x=-8820000;
#10;x=-8810000;
#10;x=-8800000;
#10;x=-8790000;
#10;x=-8780000;
#10;x=-8770000;
#10;x=-8760000;
#10;x=-8750000;
#10;x=-8740000;
#10;x=-8730000;
#10;x=-8720000;
#10;x=-8710000;
#10;x=-8700000;
#10;x=-8690000;
#10;x=-8680000;
#10;x=-8670000;
#10;x=-8660000;
#10;x=-8650000;
#10;x=-8640000;
#10;x=-8630000;
#10;x=-8620000;
#10;x=-8610000;
#10;x=-8600000;
#10;x=-8590000;
#10;x=-8580000;
#10;x=-8570000;
#10;x=-8560000;
#10;x=-8550000;
#10;x=-8540000;
#10;x=-8530000;
#10;x=-8520000;
#10;x=-8510000;
#10;x=-8500000;
#10;x=-8490000;
#10;x=-8480000;
#10;x=-8470000;
#10;x=-8460000;
#10;x=-8450000;
#10;x=-8440000;
#10;x=-8430000;
#10;x=-8420000;
#10;x=-8410000;
#10;x=-8400000;
#10;x=-8390000;
#10;x=-8380000;
#10;x=-8370000;
#10;x=-8360000;
#10;x=-8350000;
#10;x=-8340000;
#10;x=-8330000;
#10;x=-8320000;
#10;x=-8310000;
#10;x=-8300000;
#10;x=-8290000;
#10;x=-8280000;
#10;x=-8270000;
#10;x=-8260000;
#10;x=-8250000;
#10;x=-8240000;
#10;x=-8230000;
#10;x=-8220000;
#10;x=-8210000;
#10;x=-8200000;
#10;x=-8190000;
#10;x=-8180000;
#10;x=-8170000;
#10;x=-8160000;
#10;x=-8150000;
#10;x=-8140000;
#10;x=-8130000;
#10;x=-8120000;
#10;x=-8110000;
#10;x=-8100000;
#10;x=-8090000;
#10;x=-8080000;
#10;x=-8070000;
#10;x=-8060000;
#10;x=-8050000;
#10;x=-8040000;
#10;x=-8030000;
#10;x=-8020000;
#10;x=-8010000;
#10;x=-8000000;
#10;x=-7990000;
#10;x=-7980000;
#10;x=-7970000;
#10;x=-7960000;
#10;x=-7950000;
#10;x=-7940000;
#10;x=-7930000;
#10;x=-7920000;
#10;x=-7910000;
#10;x=-7900000;
#10;x=-7890000;
#10;x=-7880000;
#10;x=-7870000;
#10;x=-7860000;
#10;x=-7850000;
#10;x=-7840000;
#10;x=-7830000;
#10;x=-7820000;
#10;x=-7810000;
#10;x=-7800000;
#10;x=-7790000;
#10;x=-7780000;
#10;x=-7770000;
#10;x=-7760000;
#10;x=-7750000;
#10;x=-7740000;
#10;x=-7730000;
#10;x=-7720000;
#10;x=-7710000;
#10;x=-7700000;
#10;x=-7690000;
#10;x=-7680000;
#10;x=-7670000;
#10;x=-7660000;
#10;x=-7650000;
#10;x=-7640000;
#10;x=-7630000;
#10;x=-7620000;
#10;x=-7610000;
#10;x=-7600000;
#10;x=-7590000;
#10;x=-7580000;
#10;x=-7570000;
#10;x=-7560000;
#10;x=-7550000;
#10;x=-7540000;
#10;x=-7530000;
#10;x=-7520000;
#10;x=-7510000;
#10;x=-7500000;
#10;x=-7490000;
#10;x=-7480000;
#10;x=-7470000;
#10;x=-7460000;
#10;x=-7450000;
#10;x=-7440000;
#10;x=-7430000;
#10;x=-7420000;
#10;x=-7410000;
#10;x=-7400000;
#10;x=-7390000;
#10;x=-7380000;
#10;x=-7370000;
#10;x=-7360000;
#10;x=-7350000;
#10;x=-7340000;
#10;x=-7330000;
#10;x=-7320000;
#10;x=-7310000;
#10;x=-7300000;
#10;x=-7290000;
#10;x=-7280000;
#10;x=-7270000;
#10;x=-7260000;
#10;x=-7250000;
#10;x=-7240000;
#10;x=-7230000;
#10;x=-7220000;
#10;x=-7210000;
#10;x=-7200000;
#10;x=-7190000;
#10;x=-7180000;
#10;x=-7170000;
#10;x=-7160000;
#10;x=-7150000;
#10;x=-7140000;
#10;x=-7130000;
#10;x=-7120000;
#10;x=-7110000;
#10;x=-7100000;
#10;x=-7090000;
#10;x=-7080000;
#10;x=-7070000;
#10;x=-7060000;
#10;x=-7050000;
#10;x=-7040000;
#10;x=-7030000;
#10;x=-7020000;
#10;x=-7010000;
#10;x=-7000000;
#10;x=-6990000;
#10;x=-6980000;
#10;x=-6970000;
#10;x=-6960000;
#10;x=-6950000;
#10;x=-6940000;
#10;x=-6930000;
#10;x=-6920000;
#10;x=-6910000;
#10;x=-6900000;
#10;x=-6890000;
#10;x=-6880000;
#10;x=-6870000;
#10;x=-6860000;
#10;x=-6850000;
#10;x=-6840000;
#10;x=-6830000;
#10;x=-6820000;
#10;x=-6810000;
#10;x=-6800000;
#10;x=-6790000;
#10;x=-6780000;
#10;x=-6770000;
#10;x=-6760000;
#10;x=-6750000;
#10;x=-6740000;
#10;x=-6730000;
#10;x=-6720000;
#10;x=-6710000;
#10;x=-6700000;
#10;x=-6690000;
#10;x=-6680000;
#10;x=-6670000;
#10;x=-6660000;
#10;x=-6650000;
#10;x=-6640000;
#10;x=-6630000;
#10;x=-6620000;
#10;x=-6610000;
#10;x=-6600000;
#10;x=-6590000;
#10;x=-6580000;
#10;x=-6570000;
#10;x=-6560000;
#10;x=-6550000;
#10;x=-6540000;
#10;x=-6530000;
#10;x=-6520000;
#10;x=-6510000;
#10;x=-6500000;
#10;x=-6490000;
#10;x=-6480000;
#10;x=-6470000;
#10;x=-6460000;
#10;x=-6450000;
#10;x=-6440000;
#10;x=-6430000;
#10;x=-6420000;
#10;x=-6410000;
#10;x=-6400000;
#10;x=-6390000;
#10;x=-6380000;
#10;x=-6370000;
#10;x=-6360000;
#10;x=-6350000;
#10;x=-6340000;
#10;x=-6330000;
#10;x=-6320000;
#10;x=-6310000;
#10;x=-6300000;
#10;x=-6290000;
#10;x=-6280000;
#10;x=-6270000;
#10;x=-6260000;
#10;x=-6250000;
#10;x=-6240000;
#10;x=-6230000;
#10;x=-6220000;
#10;x=-6210000;
#10;x=-6200000;
#10;x=-6190000;
#10;x=-6180000;
#10;x=-6170000;
#10;x=-6160000;
#10;x=-6150000;
#10;x=-6140000;
#10;x=-6130000;
#10;x=-6120000;
#10;x=-6110000;
#10;x=-6100000;
#10;x=-6090000;
#10;x=-6080000;
#10;x=-6070000;
#10;x=-6060000;
#10;x=-6050000;
#10;x=-6040000;
#10;x=-6030000;
#10;x=-6020000;
#10;x=-6010000;
#10;x=-6000000;
#10;x=-5990000;
#10;x=-5980000;
#10;x=-5970000;
#10;x=-5960000;
#10;x=-5950000;
#10;x=-5940000;
#10;x=-5930000;
#10;x=-5920000;
#10;x=-5910000;
#10;x=-5900000;
#10;x=-5890000;
#10;x=-5880000;
#10;x=-5870000;
#10;x=-5860000;
#10;x=-5850000;
#10;x=-5840000;
#10;x=-5830000;
#10;x=-5820000;
#10;x=-5810000;
#10;x=-5800000;
#10;x=-5790000;
#10;x=-5780000;
#10;x=-5770000;
#10;x=-5760000;
#10;x=-5750000;
#10;x=-5740000;
#10;x=-5730000;
#10;x=-5720000;
#10;x=-5710000;
#10;x=-5700000;
#10;x=-5690000;
#10;x=-5680000;
#10;x=-5670000;
#10;x=-5660000;
#10;x=-5650000;
#10;x=-5640000;
#10;x=-5630000;
#10;x=-5620000;
#10;x=-5610000;
#10;x=-5600000;
#10;x=-5590000;
#10;x=-5580000;
#10;x=-5570000;
#10;x=-5560000;
#10;x=-5550000;
#10;x=-5540000;
#10;x=-5530000;
#10;x=-5520000;
#10;x=-5510000;
#10;x=-5500000;
#10;x=-5490000;
#10;x=-5480000;
#10;x=-5470000;
#10;x=-5460000;
#10;x=-5450000;
#10;x=-5440000;
#10;x=-5430000;
#10;x=-5420000;
#10;x=-5410000;
#10;x=-5400000;
#10;x=-5390000;
#10;x=-5380000;
#10;x=-5370000;
#10;x=-5360000;
#10;x=-5350000;
#10;x=-5340000;
#10;x=-5330000;
#10;x=-5320000;
#10;x=-5310000;
#10;x=-5300000;
#10;x=-5290000;
#10;x=-5280000;
#10;x=-5270000;
#10;x=-5260000;
#10;x=-5250000;
#10;x=-5240000;
#10;x=-5230000;
#10;x=-5220000;
#10;x=-5210000;
#10;x=-5200000;
#10;x=-5190000;
#10;x=-5180000;
#10;x=-5170000;
#10;x=-5160000;
#10;x=-5150000;
#10;x=-5140000;
#10;x=-5130000;
#10;x=-5120000;
#10;x=-5110000;
#10;x=-5100000;
#10;x=-5090000;
#10;x=-5080000;
#10;x=-5070000;
#10;x=-5060000;
#10;x=-5050000;
#10;x=-5040000;
#10;x=-5030000;
#10;x=-5020000;
#10;x=-5010000;
#10;x=-5000000;
#10;x=-4990000;
#10;x=-4980000;
#10;x=-4970000;
#10;x=-4960000;
#10;x=-4950000;
#10;x=-4940000;
#10;x=-4930000;
#10;x=-4920000;
#10;x=-4910000;
#10;x=-4900000;
#10;x=-4890000;
#10;x=-4880000;
#10;x=-4870000;
#10;x=-4860000;
#10;x=-4850000;
#10;x=-4840000;
#10;x=-4830000;
#10;x=-4820000;
#10;x=-4810000;
#10;x=-4800000;
#10;x=-4790000;
#10;x=-4780000;
#10;x=-4770000;
#10;x=-4760000;
#10;x=-4750000;
#10;x=-4740000;
#10;x=-4730000;
#10;x=-4720000;
#10;x=-4710000;
#10;x=-4700000;
#10;x=-4690000;
#10;x=-4680000;
#10;x=-4670000;
#10;x=-4660000;
#10;x=-4650000;
#10;x=-4640000;
#10;x=-4630000;
#10;x=-4620000;
#10;x=-4610000;
#10;x=-4600000;
#10;x=-4590000;
#10;x=-4580000;
#10;x=-4570000;
#10;x=-4560000;
#10;x=-4550000;
#10;x=-4540000;
#10;x=-4530000;
#10;x=-4520000;
#10;x=-4510000;
#10;x=-4500000;
#10;x=-4490000;
#10;x=-4480000;
#10;x=-4470000;
#10;x=-4460000;
#10;x=-4450000;
#10;x=-4440000;
#10;x=-4430000;
#10;x=-4420000;
#10;x=-4410000;
#10;x=-4400000;
#10;x=-4390000;
#10;x=-4380000;
#10;x=-4370000;
#10;x=-4360000;
#10;x=-4350000;
#10;x=-4340000;
#10;x=-4330000;
#10;x=-4320000;
#10;x=-4310000;
#10;x=-4300000;
#10;x=-4290000;
#10;x=-4280000;
#10;x=-4270000;
#10;x=-4260000;
#10;x=-4250000;
#10;x=-4240000;
#10;x=-4230000;
#10;x=-4220000;
#10;x=-4210000;
#10;x=-4200000;
#10;x=-4190000;
#10;x=-4180000;
#10;x=-4170000;
#10;x=-4160000;
#10;x=-4150000;
#10;x=-4140000;
#10;x=-4130000;
#10;x=-4120000;
#10;x=-4110000;
#10;x=-4100000;
#10;x=-4090000;
#10;x=-4080000;
#10;x=-4070000;
#10;x=-4060000;
#10;x=-4050000;
#10;x=-4040000;
#10;x=-4030000;
#10;x=-4020000;
#10;x=-4010000;
#10;x=-4000000;
#10;x=-3990000;
#10;x=-3980000;
#10;x=-3970000;
#10;x=-3960000;
#10;x=-3950000;
#10;x=-3940000;
#10;x=-3930000;
#10;x=-3920000;
#10;x=-3910000;
#10;x=-3900000;
#10;x=-3890000;
#10;x=-3880000;
#10;x=-3870000;
#10;x=-3860000;
#10;x=-3850000;
#10;x=-3840000;
#10;x=-3830000;
#10;x=-3820000;
#10;x=-3810000;
#10;x=-3800000;
#10;x=-3790000;
#10;x=-3780000;
#10;x=-3770000;
#10;x=-3760000;
#10;x=-3750000;
#10;x=-3740000;
#10;x=-3730000;
#10;x=-3720000;
#10;x=-3710000;
#10;x=-3700000;
#10;x=-3690000;
#10;x=-3680000;
#10;x=-3670000;
#10;x=-3660000;
#10;x=-3650000;
#10;x=-3640000;
#10;x=-3630000;
#10;x=-3620000;
#10;x=-3610000;
#10;x=-3600000;
#10;x=-3590000;
#10;x=-3580000;
#10;x=-3570000;
#10;x=-3560000;
#10;x=-3550000;
#10;x=-3540000;
#10;x=-3530000;
#10;x=-3520000;
#10;x=-3510000;
#10;x=-3500000;
#10;x=-3490000;
#10;x=-3480000;
#10;x=-3470000;
#10;x=-3460000;
#10;x=-3450000;
#10;x=-3440000;
#10;x=-3430000;
#10;x=-3420000;
#10;x=-3410000;
#10;x=-3400000;
#10;x=-3390000;
#10;x=-3380000;
#10;x=-3370000;
#10;x=-3360000;
#10;x=-3350000;
#10;x=-3340000;
#10;x=-3330000;
#10;x=-3320000;
#10;x=-3310000;
#10;x=-3300000;
#10;x=-3290000;
#10;x=-3280000;
#10;x=-3270000;
#10;x=-3260000;
#10;x=-3250000;
#10;x=-3240000;
#10;x=-3230000;
#10;x=-3220000;
#10;x=-3210000;
#10;x=-3200000;
#10;x=-3190000;
#10;x=-3180000;
#10;x=-3170000;
#10;x=-3160000;
#10;x=-3150000;
#10;x=-3140000;
#10;x=-3130000;
#10;x=-3120000;
#10;x=-3110000;
#10;x=-3100000;
#10;x=-3090000;
#10;x=-3080000;
#10;x=-3070000;
#10;x=-3060000;
#10;x=-3050000;
#10;x=-3040000;
#10;x=-3030000;
#10;x=-3020000;
#10;x=-3010000;
#10;x=-3000000;
#10;x=-2990000;
#10;x=-2980000;
#10;x=-2970000;
#10;x=-2960000;
#10;x=-2950000;
#10;x=-2940000;
#10;x=-2930000;
#10;x=-2920000;
#10;x=-2910000;
#10;x=-2900000;
#10;x=-2890000;
#10;x=-2880000;
#10;x=-2870000;
#10;x=-2860000;
#10;x=-2850000;
#10;x=-2840000;
#10;x=-2830000;
#10;x=-2820000;
#10;x=-2810000;
#10;x=-2800000;
#10;x=-2790000;
#10;x=-2780000;
#10;x=-2770000;
#10;x=-2760000;
#10;x=-2750000;
#10;x=-2740000;
#10;x=-2730000;
#10;x=-2720000;
#10;x=-2710000;
#10;x=-2700000;
#10;x=-2690000;
#10;x=-2680000;
#10;x=-2670000;
#10;x=-2660000;
#10;x=-2650000;
#10;x=-2640000;
#10;x=-2630000;
#10;x=-2620000;
#10;x=-2610000;
#10;x=-2600000;
#10;x=-2590000;
#10;x=-2580000;
#10;x=-2570000;
#10;x=-2560000;
#10;x=-2550000;
#10;x=-2540000;
#10;x=-2530000;
#10;x=-2520000;
#10;x=-2510000;
#10;x=-2500000;
#10;x=-2490000;
#10;x=-2480000;
#10;x=-2470000;
#10;x=-2460000;
#10;x=-2450000;
#10;x=-2440000;
#10;x=-2430000;
#10;x=-2420000;
#10;x=-2410000;
#10;x=-2400000;
#10;x=-2390000;
#10;x=-2380000;
#10;x=-2370000;
#10;x=-2360000;
#10;x=-2350000;
#10;x=-2340000;
#10;x=-2330000;
#10;x=-2320000;
#10;x=-2310000;
#10;x=-2300000;
#10;x=-2290000;
#10;x=-2280000;
#10;x=-2270000;
#10;x=-2260000;
#10;x=-2250000;
#10;x=-2240000;
#10;x=-2230000;
#10;x=-2220000;
#10;x=-2210000;
#10;x=-2200000;
#10;x=-2190000;
#10;x=-2180000;
#10;x=-2170000;
#10;x=-2160000;
#10;x=-2150000;
#10;x=-2140000;
#10;x=-2130000;
#10;x=-2120000;
#10;x=-2110000;
#10;x=-2100000;
#10;x=-2090000;
#10;x=-2080000;
#10;x=-2070000;
#10;x=-2060000;
#10;x=-2050000;
#10;x=-2040000;
#10;x=-2030000;
#10;x=-2020000;
#10;x=-2010000;
#10;x=-2000000;
#10;x=-1990000;
#10;x=-1980000;
#10;x=-1970000;
#10;x=-1960000;
#10;x=-1950000;
#10;x=-1940000;
#10;x=-1930000;
#10;x=-1920000;
#10;x=-1910000;
#10;x=-1900000;
#10;x=-1890000;
#10;x=-1880000;
#10;x=-1870000;
#10;x=-1860000;
#10;x=-1850000;
#10;x=-1840000;
#10;x=-1830000;
#10;x=-1820000;
#10;x=-1810000;
#10;x=-1800000;
#10;x=-1790000;
#10;x=-1780000;
#10;x=-1770000;
#10;x=-1760000;
#10;x=-1750000;
#10;x=-1740000;
#10;x=-1730000;
#10;x=-1720000;
#10;x=-1710000;
#10;x=-1700000;
#10;x=-1690000;
#10;x=-1680000;
#10;x=-1670000;
#10;x=-1660000;
#10;x=-1650000;
#10;x=-1640000;
#10;x=-1630000;
#10;x=-1620000;
#10;x=-1610000;
#10;x=-1600000;
#10;x=-1590000;
#10;x=-1580000;
#10;x=-1570000;
#10;x=-1560000;
#10;x=-1550000;
#10;x=-1540000;
#10;x=-1530000;
#10;x=-1520000;
#10;x=-1510000;
#10;x=-1500000;
#10;x=-1490000;
#10;x=-1480000;
#10;x=-1470000;
#10;x=-1460000;
#10;x=-1450000;
#10;x=-1440000;
#10;x=-1430000;
#10;x=-1420000;
#10;x=-1410000;
#10;x=-1400000;
#10;x=-1390000;
#10;x=-1380000;
#10;x=-1370000;
#10;x=-1360000;
#10;x=-1350000;
#10;x=-1340000;
#10;x=-1330000;
#10;x=-1320000;
#10;x=-1310000;
#10;x=-1300000;
#10;x=-1290000;
#10;x=-1280000;
#10;x=-1270000;
#10;x=-1260000;
#10;x=-1250000;
#10;x=-1240000;
#10;x=-1230000;
#10;x=-1220000;
#10;x=-1210000;
#10;x=-1200000;
#10;x=-1190000;
#10;x=-1180000;
#10;x=-1170000;
#10;x=-1160000;
#10;x=-1150000;
#10;x=-1140000;
#10;x=-1130000;
#10;x=-1120000;
#10;x=-1110000;
#10;x=-1100000;
#10;x=-1090000;
#10;x=-1080000;
#10;x=-1070000;
#10;x=-1060000;
#10;x=-1050000;
#10;x=-1040000;
#10;x=-1030000;
#10;x=-1020000;
#10;x=-1010000;
#10;x=-1000000;
#10;x=-990000;
#10;x=-980000;
#10;x=-970000;
#10;x=-960000;
#10;x=-950000;
#10;x=-940000;
#10;x=-930000;
#10;x=-920000;
#10;x=-910000;
#10;x=-900000;
#10;x=-890000;
#10;x=-880000;
#10;x=-870000;
#10;x=-860000;
#10;x=-850000;
#10;x=-840000;
#10;x=-830000;
#10;x=-820000;
#10;x=-810000;
#10;x=-800000;
#10;x=-790000;
#10;x=-780000;
#10;x=-770000;
#10;x=-760000;
#10;x=-750000;
#10;x=-740000;
#10;x=-730000;
#10;x=-720000;
#10;x=-710000;
#10;x=-700000;
#10;x=-690000;
#10;x=-680000;
#10;x=-670000;
#10;x=-660000;
#10;x=-650000;
#10;x=-640000;
#10;x=-630000;
#10;x=-620000;
#10;x=-610000;
#10;x=-600000;
#10;x=-590000;
#10;x=-580000;
#10;x=-570000;
#10;x=-560000;
#10;x=-550000;
#10;x=-540000;
#10;x=-530000;
#10;x=-520000;
#10;x=-510000;
#10;x=-500000;
#10;x=-490000;
#10;x=-480000;
#10;x=-470000;
#10;x=-460000;
#10;x=-450000;
#10;x=-440000;
#10;x=-430000;
#10;x=-420000;
#10;x=-410000;
#10;x=-400000;
#10;x=-390000;
#10;x=-380000;
#10;x=-370000;
#10;x=-360000;
#10;x=-350000;
#10;x=-340000;
#10;x=-330000;
#10;x=-320000;
#10;x=-310000;
#10;x=-300000;
#10;x=-290000;
#10;x=-280000;
#10;x=-270000;
#10;x=-260000;
#10;x=-250000;
#10;x=-240000;
#10;x=-230000;
#10;x=-220000;
#10;x=-210000;
#10;x=-200000;
#10;x=-190000;
#10;x=-180000;
#10;x=-170000;
#10;x=-160000;
#10;x=-150000;
#10;x=-140000;
#10;x=-130000;
#10;x=-120000;
#10;x=-110000;
#10;x=-100000;
#10;x=-90000;
#10;x=-80000;
#10;x=-70000;
#10;x=-60000;
#10;x=-50000;
#10;x=-40000;
#10;x=-30000;
#10;x=-20000;
#10;x=-10000;
#10;x=0;
#10;x=10000;
#10;x=20000;
#10;x=30000;
#10;x=40000;
#10;x=50000;
#10;x=60000;
#10;x=70000;
#10;x=80000;
#10;x=90000;
#10;x=100000;
#10;x=110000;
#10;x=120000;
#10;x=130000;
#10;x=140000;
#10;x=150000;
#10;x=160000;
#10;x=170000;
#10;x=180000;
#10;x=190000;
#10;x=200000;
#10;x=210000;
#10;x=220000;
#10;x=230000;
#10;x=240000;
#10;x=250000;
#10;x=260000;
#10;x=270000;
#10;x=280000;
#10;x=290000;
#10;x=300000;
#10;x=310000;
#10;x=320000;
#10;x=330000;
#10;x=340000;
#10;x=350000;
#10;x=360000;
#10;x=370000;
#10;x=380000;
#10;x=390000;
#10;x=400000;
#10;x=410000;
#10;x=420000;
#10;x=430000;
#10;x=440000;
#10;x=450000;
#10;x=460000;
#10;x=470000;
#10;x=480000;
#10;x=490000;
#10;x=500000;
#10;x=510000;
#10;x=520000;
#10;x=530000;
#10;x=540000;
#10;x=550000;
#10;x=560000;
#10;x=570000;
#10;x=580000;
#10;x=590000;
#10;x=600000;
#10;x=610000;
#10;x=620000;
#10;x=630000;
#10;x=640000;
#10;x=650000;
#10;x=660000;
#10;x=670000;
#10;x=680000;
#10;x=690000;
#10;x=700000;
#10;x=710000;
#10;x=720000;
#10;x=730000;
#10;x=740000;
#10;x=750000;
#10;x=760000;
#10;x=770000;
#10;x=780000;
#10;x=790000;
#10;x=800000;
#10;x=810000;
#10;x=820000;
#10;x=830000;
#10;x=840000;
#10;x=850000;
#10;x=860000;
#10;x=870000;
#10;x=880000;
#10;x=890000;
#10;x=900000;
#10;x=910000;
#10;x=920000;
#10;x=930000;
#10;x=940000;
#10;x=950000;
#10;x=960000;
#10;x=970000;
#10;x=980000;
#10;x=990000;
#10;x=1000000;
#10;x=1010000;
#10;x=1020000;
#10;x=1030000;
#10;x=1040000;
#10;x=1050000;
#10;x=1060000;
#10;x=1070000;
#10;x=1080000;
#10;x=1090000;
#10;x=1100000;
#10;x=1110000;
#10;x=1120000;
#10;x=1130000;
#10;x=1140000;
#10;x=1150000;
#10;x=1160000;
#10;x=1170000;
#10;x=1180000;
#10;x=1190000;
#10;x=1200000;
#10;x=1210000;
#10;x=1220000;
#10;x=1230000;
#10;x=1240000;
#10;x=1250000;
#10;x=1260000;
#10;x=1270000;
#10;x=1280000;
#10;x=1290000;
#10;x=1300000;
#10;x=1310000;
#10;x=1320000;
#10;x=1330000;
#10;x=1340000;
#10;x=1350000;
#10;x=1360000;
#10;x=1370000;
#10;x=1380000;
#10;x=1390000;
#10;x=1400000;
#10;x=1410000;
#10;x=1420000;
#10;x=1430000;
#10;x=1440000;
#10;x=1450000;
#10;x=1460000;
#10;x=1470000;
#10;x=1480000;
#10;x=1490000;
#10;x=1500000;
#10;x=1510000;
#10;x=1520000;
#10;x=1530000;
#10;x=1540000;
#10;x=1550000;
#10;x=1560000;
#10;x=1570000;
#10;x=1580000;
#10;x=1590000;
#10;x=1600000;
#10;x=1610000;
#10;x=1620000;
#10;x=1630000;
#10;x=1640000;
#10;x=1650000;
#10;x=1660000;
#10;x=1670000;
#10;x=1680000;
#10;x=1690000;
#10;x=1700000;
#10;x=1710000;
#10;x=1720000;
#10;x=1730000;
#10;x=1740000;
#10;x=1750000;
#10;x=1760000;
#10;x=1770000;
#10;x=1780000;
#10;x=1790000;
#10;x=1800000;
#10;x=1810000;
#10;x=1820000;
#10;x=1830000;
#10;x=1840000;
#10;x=1850000;
#10;x=1860000;
#10;x=1870000;
#10;x=1880000;
#10;x=1890000;
#10;x=1900000;
#10;x=1910000;
#10;x=1920000;
#10;x=1930000;
#10;x=1940000;
#10;x=1950000;
#10;x=1960000;
#10;x=1970000;
#10;x=1980000;
#10;x=1990000;
#10;x=2000000;
#10;x=2010000;
#10;x=2020000;
#10;x=2030000;
#10;x=2040000;
#10;x=2050000;
#10;x=2060000;
#10;x=2070000;
#10;x=2080000;
#10;x=2090000;
#10;x=2100000;
#10;x=2110000;
#10;x=2120000;
#10;x=2130000;
#10;x=2140000;
#10;x=2150000;
#10;x=2160000;
#10;x=2170000;
#10;x=2180000;
#10;x=2190000;
#10;x=2200000;
#10;x=2210000;
#10;x=2220000;
#10;x=2230000;
#10;x=2240000;
#10;x=2250000;
#10;x=2260000;
#10;x=2270000;
#10;x=2280000;
#10;x=2290000;
#10;x=2300000;
#10;x=2310000;
#10;x=2320000;
#10;x=2330000;
#10;x=2340000;
#10;x=2350000;
#10;x=2360000;
#10;x=2370000;
#10;x=2380000;
#10;x=2390000;
#10;x=2400000;
#10;x=2410000;
#10;x=2420000;
#10;x=2430000;
#10;x=2440000;
#10;x=2450000;
#10;x=2460000;
#10;x=2470000;
#10;x=2480000;
#10;x=2490000;
#10;x=2500000;
#10;x=2510000;
#10;x=2520000;
#10;x=2530000;
#10;x=2540000;
#10;x=2550000;
#10;x=2560000;
#10;x=2570000;
#10;x=2580000;
#10;x=2590000;
#10;x=2600000;
#10;x=2610000;
#10;x=2620000;
#10;x=2630000;
#10;x=2640000;
#10;x=2650000;
#10;x=2660000;
#10;x=2670000;
#10;x=2680000;
#10;x=2690000;
#10;x=2700000;
#10;x=2710000;
#10;x=2720000;
#10;x=2730000;
#10;x=2740000;
#10;x=2750000;
#10;x=2760000;
#10;x=2770000;
#10;x=2780000;
#10;x=2790000;
#10;x=2800000;
#10;x=2810000;
#10;x=2820000;
#10;x=2830000;
#10;x=2840000;
#10;x=2850000;
#10;x=2860000;
#10;x=2870000;
#10;x=2880000;
#10;x=2890000;
#10;x=2900000;
#10;x=2910000;
#10;x=2920000;
#10;x=2930000;
#10;x=2940000;
#10;x=2950000;
#10;x=2960000;
#10;x=2970000;
#10;x=2980000;
#10;x=2990000;
#10;x=3000000;
#10;x=3010000;
#10;x=3020000;
#10;x=3030000;
#10;x=3040000;
#10;x=3050000;
#10;x=3060000;
#10;x=3070000;
#10;x=3080000;
#10;x=3090000;
#10;x=3100000;
#10;x=3110000;
#10;x=3120000;
#10;x=3130000;
#10;x=3140000;
#10;x=3150000;
#10;x=3160000;
#10;x=3170000;
#10;x=3180000;
#10;x=3190000;
#10;x=3200000;
#10;x=3210000;
#10;x=3220000;
#10;x=3230000;
#10;x=3240000;
#10;x=3250000;
#10;x=3260000;
#10;x=3270000;
#10;x=3280000;
#10;x=3290000;
#10;x=3300000;
#10;x=3310000;
#10;x=3320000;
#10;x=3330000;
#10;x=3340000;
#10;x=3350000;
#10;x=3360000;
#10;x=3370000;
#10;x=3380000;
#10;x=3390000;
#10;x=3400000;
#10;x=3410000;
#10;x=3420000;
#10;x=3430000;
#10;x=3440000;
#10;x=3450000;
#10;x=3460000;
#10;x=3470000;
#10;x=3480000;
#10;x=3490000;
#10;x=3500000;
#10;x=3510000;
#10;x=3520000;
#10;x=3530000;
#10;x=3540000;
#10;x=3550000;
#10;x=3560000;
#10;x=3570000;
#10;x=3580000;
#10;x=3590000;
#10;x=3600000;
#10;x=3610000;
#10;x=3620000;
#10;x=3630000;
#10;x=3640000;
#10;x=3650000;
#10;x=3660000;
#10;x=3670000;
#10;x=3680000;
#10;x=3690000;
#10;x=3700000;
#10;x=3710000;
#10;x=3720000;
#10;x=3730000;
#10;x=3740000;
#10;x=3750000;
#10;x=3760000;
#10;x=3770000;
#10;x=3780000;
#10;x=3790000;
#10;x=3800000;
#10;x=3810000;
#10;x=3820000;
#10;x=3830000;
#10;x=3840000;
#10;x=3850000;
#10;x=3860000;
#10;x=3870000;
#10;x=3880000;
#10;x=3890000;
#10;x=3900000;
#10;x=3910000;
#10;x=3920000;
#10;x=3930000;
#10;x=3940000;
#10;x=3950000;
#10;x=3960000;
#10;x=3970000;
#10;x=3980000;
#10;x=3990000;
#10;x=4000000;
#10;x=4010000;
#10;x=4020000;
#10;x=4030000;
#10;x=4040000;
#10;x=4050000;
#10;x=4060000;
#10;x=4070000;
#10;x=4080000;
#10;x=4090000;
#10;x=4100000;
#10;x=4110000;
#10;x=4120000;
#10;x=4130000;
#10;x=4140000;
#10;x=4150000;
#10;x=4160000;
#10;x=4170000;
#10;x=4180000;
#10;x=4190000;
#10;x=4200000;
#10;x=4210000;
#10;x=4220000;
#10;x=4230000;
#10;x=4240000;
#10;x=4250000;
#10;x=4260000;
#10;x=4270000;
#10;x=4280000;
#10;x=4290000;
#10;x=4300000;
#10;x=4310000;
#10;x=4320000;
#10;x=4330000;
#10;x=4340000;
#10;x=4350000;
#10;x=4360000;
#10;x=4370000;
#10;x=4380000;
#10;x=4390000;
#10;x=4400000;
#10;x=4410000;
#10;x=4420000;
#10;x=4430000;
#10;x=4440000;
#10;x=4450000;
#10;x=4460000;
#10;x=4470000;
#10;x=4480000;
#10;x=4490000;
#10;x=4500000;
#10;x=4510000;
#10;x=4520000;
#10;x=4530000;
#10;x=4540000;
#10;x=4550000;
#10;x=4560000;
#10;x=4570000;
#10;x=4580000;
#10;x=4590000;
#10;x=4600000;
#10;x=4610000;
#10;x=4620000;
#10;x=4630000;
#10;x=4640000;
#10;x=4650000;
#10;x=4660000;
#10;x=4670000;
#10;x=4680000;
#10;x=4690000;
#10;x=4700000;
#10;x=4710000;
#10;x=4720000;
#10;x=4730000;
#10;x=4740000;
#10;x=4750000;
#10;x=4760000;
#10;x=4770000;
#10;x=4780000;
#10;x=4790000;
#10;x=4800000;
#10;x=4810000;
#10;x=4820000;
#10;x=4830000;
#10;x=4840000;
#10;x=4850000;
#10;x=4860000;
#10;x=4870000;
#10;x=4880000;
#10;x=4890000;
#10;x=4900000;
#10;x=4910000;
#10;x=4920000;
#10;x=4930000;
#10;x=4940000;
#10;x=4950000;
#10;x=4960000;
#10;x=4970000;
#10;x=4980000;
#10;x=4990000;
#10;x=5000000;
#10;x=5010000;
#10;x=5020000;
#10;x=5030000;
#10;x=5040000;
#10;x=5050000;
#10;x=5060000;
#10;x=5070000;
#10;x=5080000;
#10;x=5090000;
#10;x=5100000;
#10;x=5110000;
#10;x=5120000;
#10;x=5130000;
#10;x=5140000;
#10;x=5150000;
#10;x=5160000;
#10;x=5170000;
#10;x=5180000;
#10;x=5190000;
#10;x=5200000;
#10;x=5210000;
#10;x=5220000;
#10;x=5230000;
#10;x=5240000;
#10;x=5250000;
#10;x=5260000;
#10;x=5270000;
#10;x=5280000;
#10;x=5290000;
#10;x=5300000;
#10;x=5310000;
#10;x=5320000;
#10;x=5330000;
#10;x=5340000;
#10;x=5350000;
#10;x=5360000;
#10;x=5370000;
#10;x=5380000;
#10;x=5390000;
#10;x=5400000;
#10;x=5410000;
#10;x=5420000;
#10;x=5430000;
#10;x=5440000;
#10;x=5450000;
#10;x=5460000;
#10;x=5470000;
#10;x=5480000;
#10;x=5490000;
#10;x=5500000;
#10;x=5510000;
#10;x=5520000;
#10;x=5530000;
#10;x=5540000;
#10;x=5550000;
#10;x=5560000;
#10;x=5570000;
#10;x=5580000;
#10;x=5590000;
#10;x=5600000;
#10;x=5610000;
#10;x=5620000;
#10;x=5630000;
#10;x=5640000;
#10;x=5650000;
#10;x=5660000;
#10;x=5670000;
#10;x=5680000;
#10;x=5690000;
#10;x=5700000;
#10;x=5710000;
#10;x=5720000;
#10;x=5730000;
#10;x=5740000;
#10;x=5750000;
#10;x=5760000;
#10;x=5770000;
#10;x=5780000;
#10;x=5790000;
#10;x=5800000;
#10;x=5810000;
#10;x=5820000;
#10;x=5830000;
#10;x=5840000;
#10;x=5850000;
#10;x=5860000;
#10;x=5870000;
#10;x=5880000;
#10;x=5890000;
#10;x=5900000;
#10;x=5910000;
#10;x=5920000;
#10;x=5930000;
#10;x=5940000;
#10;x=5950000;
#10;x=5960000;
#10;x=5970000;
#10;x=5980000;
#10;x=5990000;
#10;x=6000000;
#10;x=6010000;
#10;x=6020000;
#10;x=6030000;
#10;x=6040000;
#10;x=6050000;
#10;x=6060000;
#10;x=6070000;
#10;x=6080000;
#10;x=6090000;
#10;x=6100000;
#10;x=6110000;
#10;x=6120000;
#10;x=6130000;
#10;x=6140000;
#10;x=6150000;
#10;x=6160000;
#10;x=6170000;
#10;x=6180000;
#10;x=6190000;
#10;x=6200000;
#10;x=6210000;
#10;x=6220000;
#10;x=6230000;
#10;x=6240000;
#10;x=6250000;
#10;x=6260000;
#10;x=6270000;
#10;x=6280000;
#10;x=6290000;
#10;x=6300000;
#10;x=6310000;
#10;x=6320000;
#10;x=6330000;
#10;x=6340000;
#10;x=6350000;
#10;x=6360000;
#10;x=6370000;
#10;x=6380000;
#10;x=6390000;
#10;x=6400000;
#10;x=6410000;
#10;x=6420000;
#10;x=6430000;
#10;x=6440000;
#10;x=6450000;
#10;x=6460000;
#10;x=6470000;
#10;x=6480000;
#10;x=6490000;
#10;x=6500000;
#10;x=6510000;
#10;x=6520000;
#10;x=6530000;
#10;x=6540000;
#10;x=6550000;
#10;x=6560000;
#10;x=6570000;
#10;x=6580000;
#10;x=6590000;
#10;x=6600000;
#10;x=6610000;
#10;x=6620000;
#10;x=6630000;
#10;x=6640000;
#10;x=6650000;
#10;x=6660000;
#10;x=6670000;
#10;x=6680000;
#10;x=6690000;
#10;x=6700000;
#10;x=6710000;
#10;x=6720000;
#10;x=6730000;
#10;x=6740000;
#10;x=6750000;
#10;x=6760000;
#10;x=6770000;
#10;x=6780000;
#10;x=6790000;
#10;x=6800000;
#10;x=6810000;
#10;x=6820000;
#10;x=6830000;
#10;x=6840000;
#10;x=6850000;
#10;x=6860000;
#10;x=6870000;
#10;x=6880000;
#10;x=6890000;
#10;x=6900000;
#10;x=6910000;
#10;x=6920000;
#10;x=6930000;
#10;x=6940000;
#10;x=6950000;
#10;x=6960000;
#10;x=6970000;
#10;x=6980000;
#10;x=6990000;
#10;x=7000000;
#10;x=7010000;
#10;x=7020000;
#10;x=7030000;
#10;x=7040000;
#10;x=7050000;
#10;x=7060000;
#10;x=7070000;
#10;x=7080000;
#10;x=7090000;
#10;x=7100000;
#10;x=7110000;
#10;x=7120000;
#10;x=7130000;
#10;x=7140000;
#10;x=7150000;
#10;x=7160000;
#10;x=7170000;
#10;x=7180000;
#10;x=7190000;
#10;x=7200000;
#10;x=7210000;
#10;x=7220000;
#10;x=7230000;
#10;x=7240000;
#10;x=7250000;
#10;x=7260000;
#10;x=7270000;
#10;x=7280000;
#10;x=7290000;
#10;x=7300000;
#10;x=7310000;
#10;x=7320000;
#10;x=7330000;
#10;x=7340000;
#10;x=7350000;
#10;x=7360000;
#10;x=7370000;
#10;x=7380000;
#10;x=7390000;
#10;x=7400000;
#10;x=7410000;
#10;x=7420000;
#10;x=7430000;
#10;x=7440000;
#10;x=7450000;
#10;x=7460000;
#10;x=7470000;
#10;x=7480000;
#10;x=7490000;
#10;x=7500000;
#10;x=7510000;
#10;x=7520000;
#10;x=7530000;
#10;x=7540000;
#10;x=7550000;
#10;x=7560000;
#10;x=7570000;
#10;x=7580000;
#10;x=7590000;
#10;x=7600000;
#10;x=7610000;
#10;x=7620000;
#10;x=7630000;
#10;x=7640000;
#10;x=7650000;
#10;x=7660000;
#10;x=7670000;
#10;x=7680000;
#10;x=7690000;
#10;x=7700000;
#10;x=7710000;
#10;x=7720000;
#10;x=7730000;
#10;x=7740000;
#10;x=7750000;
#10;x=7760000;
#10;x=7770000;
#10;x=7780000;
#10;x=7790000;
#10;x=7800000;
#10;x=7810000;
#10;x=7820000;
#10;x=7830000;
#10;x=7840000;
#10;x=7850000;
#10;x=7860000;
#10;x=7870000;
#10;x=7880000;
#10;x=7890000;
#10;x=7900000;
#10;x=7910000;
#10;x=7920000;
#10;x=7930000;
#10;x=7940000;
#10;x=7950000;
#10;x=7960000;
#10;x=7970000;
#10;x=7980000;
#10;x=7990000;
#10;x=8000000;
#10;x=8010000;
#10;x=8020000;
#10;x=8030000;
#10;x=8040000;
#10;x=8050000;
#10;x=8060000;
#10;x=8070000;
#10;x=8080000;
#10;x=8090000;
#10;x=8100000;
#10;x=8110000;
#10;x=8120000;
#10;x=8130000;
#10;x=8140000;
#10;x=8150000;
#10;x=8160000;
#10;x=8170000;
#10;x=8180000;
#10;x=8190000;
#10;x=8200000;
#10;x=8210000;
#10;x=8220000;
#10;x=8230000;
#10;x=8240000;
#10;x=8250000;
#10;x=8260000;
#10;x=8270000;
#10;x=8280000;
#10;x=8290000;
#10;x=8300000;
#10;x=8310000;
#10;x=8320000;
#10;x=8330000;
#10;x=8340000;
#10;x=8350000;
#10;x=8360000;
#10;x=8370000;
#10;x=8380000;
#10;x=8390000;
#10;x=8400000;
#10;x=8410000;
#10;x=8420000;
#10;x=8430000;
#10;x=8440000;
#10;x=8450000;
#10;x=8460000;
#10;x=8470000;
#10;x=8480000;
#10;x=8490000;
#10;x=8500000;
#10;x=8510000;
#10;x=8520000;
#10;x=8530000;
#10;x=8540000;
#10;x=8550000;
#10;x=8560000;
#10;x=8570000;
#10;x=8580000;
#10;x=8590000;
#10;x=8600000;
#10;x=8610000;
#10;x=8620000;
#10;x=8630000;
#10;x=8640000;
#10;x=8650000;
#10;x=8660000;
#10;x=8670000;
#10;x=8680000;
#10;x=8690000;
#10;x=8700000;
#10;x=8710000;
#10;x=8720000;
#10;x=8730000;
#10;x=8740000;
#10;x=8750000;
#10;x=8760000;
#10;x=8770000;
#10;x=8780000;
#10;x=8790000;
#10;x=8800000;
#10;x=8810000;
#10;x=8820000;
#10;x=8830000;
#10;x=8840000;
#10;x=8850000;
#10;x=8860000;
#10;x=8870000;
#10;x=8880000;
#10;x=8890000;
#10;x=8900000;
#10;x=8910000;
#10;x=8920000;
#10;x=8930000;
#10;x=8940000;
#10;x=8950000;
#10;x=8960000;
#10;x=8970000;
#10;x=8980000;
#10;x=8990000;
#10;x=9000000;
#10;x=9010000;
#10;x=9020000;
#10;x=9030000;
#10;x=9040000;
#10;x=9050000;
#10;x=9060000;
#10;x=9070000;
#10;x=9080000;
#10;x=9090000;
#10;x=9100000;
#10;x=9110000;
#10;x=9120000;
#10;x=9130000;
#10;x=9140000;
#10;x=9150000;
#10;x=9160000;
#10;x=9170000;
#10;x=9180000;
#10;x=9190000;
#10;x=9200000;
#10;x=9210000;
#10;x=9220000;
#10;x=9230000;
#10;x=9240000;
#10;x=9250000;
#10;x=9260000;
#10;x=9270000;
#10;x=9280000;
#10;x=9290000;
#10;x=9300000;
#10;x=9310000;
#10;x=9320000;
#10;x=9330000;
#10;x=9340000;
#10;x=9350000;
#10;x=9360000;
#10;x=9370000;
#10;x=9380000;
#10;x=9390000;
#10;x=9400000;
#10;x=9410000;
#10;x=9420000;
#10;x=9430000;
#10;x=9440000;
#10;x=9450000;
#10;x=9460000;
#10;x=9470000;
#10;x=9480000;
#10;x=9490000;
#10;x=9500000;
#10;x=9510000;
#10;x=9520000;
#10;x=9530000;
#10;x=9540000;
#10;x=9550000;
#10;x=9560000;
#10;x=9570000;
#10;x=9580000;
#10;x=9590000;
#10;x=9600000;
#10;x=9610000;
#10;x=9620000;
#10;x=9630000;
#10;x=9640000;
#10;x=9650000;
#10;x=9660000;
#10;x=9670000;
#10;x=9680000;
#10;x=9690000;
#10;x=9700000;
#10;x=9710000;
#10;x=9720000;
#10;x=9730000;
#10;x=9740000;
#10;x=9750000;
#10;x=9760000;
#10;x=9770000;
#10;x=9780000;
#10;x=9790000;
#10;x=9800000;
#10;x=9810000;
#10;x=9820000;
#10;x=9830000;
#10;x=9840000;
#10;x=9850000;
#10;x=9860000;
#10;x=9870000;
#10;x=9880000;
#10;x=9890000;
#10;x=9900000;
#10;x=9910000;
#10;x=9920000;
#10;x=9930000;
#10;x=9940000;
#10;x=9950000;
#10;x=9960000;
#10;x=9970000;
#10;x=9980000;
#10;x=9990000;
#10;x=10000000;
#10;x=10010000;
#10;x=10020000;
#10;x=10030000;
#10;x=10040000;
#10;x=10050000;
#10;x=10060000;
#10;x=10070000;
#10;x=10080000;
#10;x=10090000;
#10;x=10100000;
#10;x=10110000;
#10;x=10120000;
#10;x=10130000;
#10;x=10140000;
#10;x=10150000;
#10;x=10160000;
#10;x=10170000;
#10;x=10180000;
#10;x=10190000;
#10;x=10200000;
#10;x=10210000;
#10;x=10220000;
#10;x=10230000;
#10;x=10240000;
#10;x=10250000;
#10;x=10260000;
#10;x=10270000;
#10;x=10280000;
#10;x=10290000;
#10;x=10300000;
#10;x=10310000;
#10;x=10320000;
#10;x=10330000;
#10;x=10340000;
#10;x=10350000;
#10;x=10360000;
#10;x=10370000;
#10;x=10380000;
#10;x=10390000;
#10;x=10400000;
#10;x=10410000;
#10;x=10420000;
#10;x=10430000;
#10;x=10440000;
#10;x=10450000;
#10;x=10460000;
#10;x=10470000;
#10;x=10480000;
#10;x=10490000;
#10;x=10500000;
#10;x=10510000;
#10;x=10520000;
#10;x=10530000;
#10;x=10540000;
#10;x=10550000;
#10;x=10560000;
#10;x=10570000;
#10;x=10580000;
#10;x=10590000;
#10;x=10600000;
#10;x=10610000;
#10;x=10620000;
#10;x=10630000;
#10;x=10640000;
#10;x=10650000;
#10;x=10660000;
#10;x=10670000;
#10;x=10680000;
#10;x=10690000;
#10;x=10700000;
#10;x=10710000;
#10;x=10720000;
#10;x=10730000;
#10;x=10740000;
#10;x=10750000;
#10;x=10760000;
#10;x=10770000;
#10;x=10780000;
#10;x=10790000;
#10;x=10800000;
#10;x=10810000;
#10;x=10820000;
#10;x=10830000;
#10;x=10840000;
#10;x=10850000;
#10;x=10860000;
#10;x=10870000;
#10;x=10880000;
#10;x=10890000;
#10;x=10900000;
#10;x=10910000;
#10;x=10920000;
#10;x=10930000;
#10;x=10940000;
#10;x=10950000;
#10;x=10960000;
#10;x=10970000;
#10;x=10980000;
#10;x=10990000;
#10;x=11000000;
#10;x=11010000;
#10;x=11020000;
#10;x=11030000;
#10;x=11040000;
#10;x=11050000;
#10;x=11060000;
#10;x=11070000;
#10;x=11080000;
#10;x=11090000;
#10;x=11100000;
#10;x=11110000;
#10;x=11120000;
#10;x=11130000;
#10;x=11140000;
#10;x=11150000;
#10;x=11160000;
#10;x=11170000;
#10;x=11180000;
#10;x=11190000;
#10;x=11200000;
#10;x=11210000;
#10;x=11220000;
#10;x=11230000;
#10;x=11240000;
#10;x=11250000;
#10;x=11260000;
#10;x=11270000;
#10;x=11280000;
#10;x=11290000;
#10;x=11300000;
#10;x=11310000;
#10;x=11320000;
#10;x=11330000;
#10;x=11340000;
#10;x=11350000;
#10;x=11360000;
#10;x=11370000;
#10;x=11380000;
#10;x=11390000;
#10;x=11400000;
#10;x=11410000;
#10;x=11420000;
#10;x=11430000;
#10;x=11440000;
#10;x=11450000;
#10;x=11460000;
#10;x=11470000;
#10;x=11480000;
#10;x=11490000;
#10;x=11500000;
#10;x=11510000;
#10;x=11520000;
#10;x=11530000;
#10;x=11540000;
#10;x=11550000;
#10;x=11560000;
#10;x=11570000;
#10;x=11580000;
#10;x=11590000;
#10;x=11600000;
#10;x=11610000;
#10;x=11620000;
#10;x=11630000;
#10;x=11640000;
#10;x=11650000;
#10;x=11660000;
#10;x=11670000;
#10;x=11680000;
#10;x=11690000;
#10;x=11700000;
#10;x=11710000;
#10;x=11720000;
#10;x=11730000;
#10;x=11740000;
#10;x=11750000;
#10;x=11760000;
#10;x=11770000;
#10;x=11780000;
#10;x=11790000;
#10;x=11800000;
#10;x=11810000;
#10;x=11820000;
#10;x=11830000;
#10;x=11840000;
#10;x=11850000;
#10;x=11860000;
#10;x=11870000;
#10;x=11880000;
#10;x=11890000;
#10;x=11900000;
#10;x=11910000;
#10;x=11920000;
#10;x=11930000;
#10;x=11940000;
#10;x=11950000;
#10;x=11960000;
#10;x=11970000;
#10;x=11980000;
#10;x=11990000;
#10;x=12000000;
#10;x=12010000;
#10;x=12020000;
#10;x=12030000;
#10;x=12040000;
#10;x=12050000;
#10;x=12060000;
#10;x=12070000;
#10;x=12080000;
#10;x=12090000;
#10;x=12100000;
#10;x=12110000;
#10;x=12120000;
#10;x=12130000;
#10;x=12140000;
#10;x=12150000;
#10;x=12160000;
#10;x=12170000;
#10;x=12180000;
#10;x=12190000;
#10;x=12200000;
#10;x=12210000;
#10;x=12220000;
#10;x=12230000;
#10;x=12240000;
#10;x=12250000;
#10;x=12260000;
#10;x=12270000;
#10;x=12280000;
#10;x=12290000;
#10;x=12300000;
#10;x=12310000;
#10;x=12320000;
#10;x=12330000;
#10;x=12340000;
#10;x=12350000;
#10;x=12360000;
#10;x=12370000;
#10;x=12380000;
#10;x=12390000;
#10;x=12400000;
#10;x=12410000;
#10;x=12420000;
#10;x=12430000;
#10;x=12440000;
#10;x=12450000;
#10;x=12460000;
#10;x=12470000;
#10;x=12480000;
#10;x=12490000;
#10;x=12500000;
#10;x=12510000;
#10;x=12520000;
#10;x=12530000;
#10;x=12540000;
#10;x=12550000;
#10;x=12560000;
#10;x=12570000;
#10;x=12580000;
#10;x=12590000;
#10;x=12600000;
#10;x=12610000;
#10;x=12620000;
#10;x=12630000;
#10;x=12640000;
#10;x=12650000;
#10;x=12660000;
#10;x=12670000;
#10;x=12680000;
#10;x=12690000;
#10;x=12700000;
#10;x=12710000;
#10;x=12720000;
#10;x=12730000;
#10;x=12740000;
#10;x=12750000;
#10;x=12760000;
#10;x=12770000;
#10;x=12780000;
#10;x=12790000;
#10;x=12800000;
#10;x=12810000;
#10;x=12820000;
#10;x=12830000;
#10;x=12840000;
#10;x=12850000;
#10;x=12860000;
#10;x=12870000;
#10;x=12880000;
#10;x=12890000;
#10;x=12900000;
#10;x=12910000;
#10;x=12920000;
#10;x=12930000;
#10;x=12940000;
#10;x=12950000;
#10;x=12960000;
#10;x=12970000;
#10;x=12980000;
#10;x=12990000;
#10;x=13000000;
#10;x=13010000;
#10;x=13020000;
#10;x=13030000;
#10;x=13040000;
#10;x=13050000;
#10;x=13060000;
#10;x=13070000;
#10;x=13080000;
#10;x=13090000;
#10;x=13100000;
#10;x=13110000;
#10;x=13120000;
#10;x=13130000;
#10;x=13140000;
#10;x=13150000;
#10;x=13160000;
#10;x=13170000;
#10;x=13180000;
#10;x=13190000;
#10;x=13200000;
#10;x=13210000;
#10;x=13220000;
#10;x=13230000;
#10;x=13240000;
#10;x=13250000;
#10;x=13260000;
#10;x=13270000;
#10;x=13280000;
#10;x=13290000;
#10;x=13300000;
#10;x=13310000;
#10;x=13320000;
#10;x=13330000;
#10;x=13340000;
#10;x=13350000;
#10;x=13360000;
#10;x=13370000;
#10;x=13380000;
#10;x=13390000;
#10;x=13400000;
#10;x=13410000;
#10;x=13420000;
#10;x=13430000;
#10;x=13440000;
#10;x=13450000;
#10;x=13460000;
#10;x=13470000;
#10;x=13480000;
#10;x=13490000;
#10;x=13500000;
#10;x=13510000;
#10;x=13520000;
#10;x=13530000;
#10;x=13540000;
#10;x=13550000;
#10;x=13560000;
#10;x=13570000;
#10;x=13580000;
#10;x=13590000;
#10;x=13600000;
#10;x=13610000;
#10;x=13620000;
#10;x=13630000;
#10;x=13640000;
#10;x=13650000;
#10;x=13660000;
#10;x=13670000;
#10;x=13680000;
#10;x=13690000;
#10;x=13700000;
#10;x=13710000;
#10;x=13720000;
#10;x=13730000;
#10;x=13740000;
#10;x=13750000;
#10;x=13760000;
#10;x=13770000;
#10;x=13780000;
#10;x=13790000;
#10;x=13800000;
#10;x=13810000;
#10;x=13820000;
#10;x=13830000;
#10;x=13840000;
#10;x=13850000;
#10;x=13860000;
#10;x=13870000;
#10;x=13880000;
#10;x=13890000;
#10;x=13900000;
#10;x=13910000;
#10;x=13920000;
#10;x=13930000;
#10;x=13940000;
#10;x=13950000;
#10;x=13960000;
#10;x=13970000;
#10;x=13980000;
#10;x=13990000;
#10;x=14000000;
#10;x=14010000;
#10;x=14020000;
#10;x=14030000;
#10;x=14040000;
#10;x=14050000;
#10;x=14060000;
#10;x=14070000;
#10;x=14080000;
#10;x=14090000;
#10;x=14100000;
#10;x=14110000;
#10;x=14120000;
#10;x=14130000;
#10;x=14140000;
#10;x=14150000;
#10;x=14160000;
#10;x=14170000;
#10;x=14180000;
#10;x=14190000;
#10;x=14200000;
#10;x=14210000;
#10;x=14220000;
#10;x=14230000;
#10;x=14240000;
#10;x=14250000;
#10;x=14260000;
#10;x=14270000;
#10;x=14280000;
#10;x=14290000;
#10;x=14300000;
#10;x=14310000;
#10;x=14320000;
#10;x=14330000;
#10;x=14340000;
#10;x=14350000;
#10;x=14360000;
#10;x=14370000;
#10;x=14380000;
#10;x=14390000;
#10;x=14400000;
#10;x=14410000;
#10;x=14420000;
#10;x=14430000;
#10;x=14440000;
#10;x=14450000;
#10;x=14460000;
#10;x=14470000;
#10;x=14480000;
#10;x=14490000;
#10;x=14500000;
#10;x=14510000;
#10;x=14520000;
#10;x=14530000;
#10;x=14540000;
#10;x=14550000;
#10;x=14560000;
#10;x=14570000;
#10;x=14580000;
#10;x=14590000;
#10;x=14600000;
#10;x=14610000;
#10;x=14620000;
#10;x=14630000;
#10;x=14640000;
#10;x=14650000;
#10;x=14660000;
#10;x=14670000;
#10;x=14680000;
#10;x=14690000;
#10;x=14700000;
#10;x=14710000;
#10;x=14720000;
#10;x=14730000;
#10;x=14740000;
#10;x=14750000;
#10;x=14760000;
#10;x=14770000;
#10;x=14780000;
#10;x=14790000;
#10;x=14800000;
#10;x=14810000;
#10;x=14820000;
#10;x=14830000;
#10;x=14840000;
#10;x=14850000;
#10;x=14860000;
#10;x=14870000;
#10;x=14880000;
#10;x=14890000;
#10;x=14900000;
#10;x=14910000;
#10;x=14920000;
#10;x=14930000;
#10;x=14940000;
#10;x=14950000;
#10;x=14960000;
#10;x=14970000;
#10;x=14980000;
#10;x=14990000;
#10;x=15000000;
#10;x=15010000;
#10;x=15020000;
#10;x=15030000;
#10;x=15040000;
#10;x=15050000;
#10;x=15060000;
#10;x=15070000;
#10;x=15080000;
#10;x=15090000;
#10;x=15100000;
#10;x=15110000;
#10;x=15120000;
#10;x=15130000;
#10;x=15140000;
#10;x=15150000;
#10;x=15160000;
#10;x=15170000;
#10;x=15180000;
#10;x=15190000;
#10;x=15200000;
#10;x=15210000;
#10;x=15220000;
#10;x=15230000;
#10;x=15240000;
#10;x=15250000;
#10;x=15260000;
#10;x=15270000;
#10;x=15280000;
#10;x=15290000;
#10;x=15300000;
#10;x=15310000;
#10;x=15320000;
#10;x=15330000;
#10;x=15340000;
#10;x=15350000;
#10;x=15360000;
#10;x=15370000;
#10;x=15380000;
#10;x=15390000;
#10;x=15400000;
#10;x=15410000;
#10;x=15420000;
#10;x=15430000;
#10;x=15440000;
#10;x=15450000;
#10;x=15460000;
#10;x=15470000;
#10;x=15480000;
#10;x=15490000;
#10;x=15500000;
#10;x=15510000;
#10;x=15520000;
#10;x=15530000;
#10;x=15540000;
#10;x=15550000;
#10;x=15560000;
#10;x=15570000;
#10;x=15580000;
#10;x=15590000;
#10;x=15600000;
#10;x=15610000;
#10;x=15620000;
#10;x=15630000;
#10;x=15640000;
#10;x=15650000;
#10;x=15660000;
#10;x=15670000;
#10;x=15680000;
#10;x=15690000;
#10;x=15700000;
#10;x=15710000;
#10;x=15720000;
#10;x=15730000;
#10;x=15740000;
#10;x=15750000;
#10;x=15760000;
#10;x=15770000;
#10;x=15780000;
#10;x=15790000;
#10;x=15800000;
#10;x=15810000;
#10;x=15820000;
#10;x=15830000;
#10;x=15840000;
#10;x=15850000;
#10;x=15860000;
#10;x=15870000;
#10;x=15880000;
#10;x=15890000;
#10;x=15900000;
#10;x=15910000;
#10;x=15920000;
#10;x=15930000;
#10;x=15940000;
#10;x=15950000;
#10;x=15960000;
#10;x=15970000;
#10;x=15980000;
#10;x=15990000;
#10;x=16000000;
#10;x=16010000;
#10;x=16020000;
#10;x=16030000;
#10;x=16040000;
#10;x=16050000;
#10;x=16060000;
#10;x=16070000;
#10;x=16080000;
#10;x=16090000;
#10;x=16100000;
#10;x=16110000;
#10;x=16120000;
#10;x=16130000;
#10;x=16140000;
#10;x=16150000;
#10;x=16160000;
#10;x=16170000;
#10;x=16180000;
#10;x=16190000;
#10;x=16200000;
#10;x=16210000;
#10;x=16220000;
#10;x=16230000;
#10;x=16240000;
#10;x=16250000;
#10;x=16260000;
#10;x=16270000;
#10;x=16280000;
#10;x=16290000;
#10;x=16300000;
#10;x=16310000;
#10;x=16320000;
#10;x=16330000;
#10;x=16340000;
#10;x=16350000;
#10;x=16360000;
#10;x=16370000;
#10;x=16380000;
#10;x=16390000;
#10;x=16400000;
#10;x=16410000;
#10;x=16420000;
#10;x=16430000;
#10;x=16440000;
#10;x=16450000;
#10;x=16460000;
#10;x=16470000;
#10;x=16480000;
#10;x=16490000;
#10;x=16500000;
#10;x=16510000;
#10;x=16520000;
#10;x=16530000;
#10;x=16540000;
#10;x=16550000;
#10;x=16560000;
#10;x=16570000;
#10;x=16580000;
#10;x=16590000;
#10;x=16600000;
#10;x=16610000;
#10;x=16620000;
#10;x=16630000;
#10;x=16640000;
#10;x=16650000;
#10;x=16660000;
#10;x=16670000;
#10;x=16680000;
#10;x=16690000;
#10;x=16700000;
#10;x=16710000;
#10;x=16720000;
#10;x=16730000;
#10;x=16740000;
#10;x=16750000;
#10;x=16760000;
#10;x=16770000;
#10;x=16780000;
#10;x=16790000;
#10;x=16800000;
#10;x=16810000;
#10;x=16820000;
#10;x=16830000;
#10;x=16840000;
#10;x=16850000;
#10;x=16860000;
#10;x=16870000;
#10;x=16880000;
#10;x=16890000;
#10;x=16900000;
#10;x=16910000;
#10;x=16920000;
#10;x=16930000;
#10;x=16940000;
#10;x=16950000;
#10;x=16960000;
#10;x=16970000;
#10;x=16980000;
#10;x=16990000;
#10;x=17000000;
#10;x=17010000;
#10;x=17020000;
#10;x=17030000;
#10;x=17040000;
#10;x=17050000;
#10;x=17060000;
#10;x=17070000;
#10;x=17080000;
#10;x=17090000;
#10;x=17100000;
#10;x=17110000;
#10;x=17120000;
#10;x=17130000;
#10;x=17140000;
#10;x=17150000;
#10;x=17160000;
#10;x=17170000;
#10;x=17180000;
#10;x=17190000;
#10;x=17200000;
#10;x=17210000;
#10;x=17220000;
#10;x=17230000;
#10;x=17240000;
#10;x=17250000;
#10;x=17260000;
#10;x=17270000;
#10;x=17280000;
#10;x=17290000;
#10;x=17300000;
#10;x=17310000;
#10;x=17320000;
#10;x=17330000;
#10;x=17340000;
#10;x=17350000;
#10;x=17360000;
#10;x=17370000;
#10;x=17380000;
#10;x=17390000;
#10;x=17400000;
#10;x=17410000;
#10;x=17420000;
#10;x=17430000;
#10;x=17440000;
#10;x=17450000;
#10;x=17460000;
#10;x=17470000;
#10;x=17480000;
#10;x=17490000;
#10;x=17500000;
#10;x=17510000;
#10;x=17520000;
#10;x=17530000;
#10;x=17540000;
#10;x=17550000;
#10;x=17560000;
#10;x=17570000;
#10;x=17580000;
#10;x=17590000;
#10;x=17600000;
#10;x=17610000;
#10;x=17620000;
#10;x=17630000;
#10;x=17640000;
#10;x=17650000;
#10;x=17660000;
#10;x=17670000;
#10;x=17680000;
#10;x=17690000;
#10;x=17700000;
#10;x=17710000;
#10;x=17720000;
#10;x=17730000;
#10;x=17740000;
#10;x=17750000;
#10;x=17760000;
#10;x=17770000;
#10;x=17780000;
#10;x=17790000;
#10;x=17800000;
#10;x=17810000;
#10;x=17820000;
#10;x=17830000;
#10;x=17840000;
#10;x=17850000;
#10;x=17860000;
#10;x=17870000;
#10;x=17880000;
#10;x=17890000;
#10;x=17900000;
#10;x=17910000;
#10;x=17920000;
#10;x=17930000;
#10;x=17940000;
#10;x=17950000;
#10;x=17960000;
#10;x=17970000;
#10;x=17980000;
#10;x=17990000;
#10;x=18000000;
#10;x=18010000;
#10;x=18020000;
#10;x=18030000;
#10;x=18040000;
#10;x=18050000;
#10;x=18060000;
#10;x=18070000;
#10;x=18080000;
#10;x=18090000;
#10;x=18100000;
#10;x=18110000;
#10;x=18120000;
#10;x=18130000;
#10;x=18140000;
#10;x=18150000;
#10;x=18160000;
#10;x=18170000;
#10;x=18180000;
#10;x=18190000;
#10;x=18200000;
#10;x=18210000;
#10;x=18220000;
#10;x=18230000;
#10;x=18240000;
#10;x=18250000;
#10;x=18260000;
#10;x=18270000;
#10;x=18280000;
#10;x=18290000;
#10;x=18300000;
#10;x=18310000;
#10;x=18320000;
#10;x=18330000;
#10;x=18340000;
#10;x=18350000;
#10;x=18360000;
#10;x=18370000;
#10;x=18380000;
#10;x=18390000;
#10;x=18400000;
#10;x=18410000;
#10;x=18420000;
#10;x=18430000;
#10;x=18440000;
#10;x=18450000;
#10;x=18460000;
#10;x=18470000;
#10;x=18480000;
#10;x=18490000;
#10;x=18500000;
#10;x=18510000;
#10;x=18520000;
#10;x=18530000;
#10;x=18540000;
#10;x=18550000;
#10;x=18560000;
#10;x=18570000;
#10;x=18580000;
#10;x=18590000;
#10;x=18600000;
#10;x=18610000;
#10;x=18620000;
#10;x=18630000;
#10;x=18640000;
#10;x=18650000;
#10;x=18660000;
#10;x=18670000;
#10;x=18680000;
#10;x=18690000;
#10;x=18700000;
#10;x=18710000;
#10;x=18720000;
#10;x=18730000;
#10;x=18740000;
#10;x=18750000;
#10;x=18760000;
#10;x=18770000;
#10;x=18780000;
#10;x=18790000;
#10;x=18800000;
#10;x=18810000;
#10;x=18820000;
#10;x=18830000;
#10;x=18840000;
#10;x=18850000;
#10;x=18860000;
#10;x=18870000;
#10;x=18880000;
#10;x=18890000;
#10;x=18900000;
#10;x=18910000;
#10;x=18920000;
#10;x=18930000;
#10;x=18940000;
#10;x=18950000;
#10;x=18960000;
#10;x=18970000;
#10;x=18980000;
#10;x=18990000;
#10;x=19000000;
#10;x=19010000;
#10;x=19020000;
#10;x=19030000;
#10;x=19040000;
#10;x=19050000;
#10;x=19060000;
#10;x=19070000;
#10;x=19080000;
#10;x=19090000;
#10;x=19100000;
#10;x=19110000;
#10;x=19120000;
#10;x=19130000;
#10;x=19140000;
#10;x=19150000;
#10;x=19160000;
#10;x=19170000;
#10;x=19180000;
#10;x=19190000;
#10;x=19200000;
#10;x=19210000;
#10;x=19220000;
#10;x=19230000;
#10;x=19240000;
#10;x=19250000;
#10;x=19260000;
#10;x=19270000;
#10;x=19280000;
#10;x=19290000;
#10;x=19300000;
#10;x=19310000;
#10;x=19320000;
#10;x=19330000;
#10;x=19340000;
#10;x=19350000;
#10;x=19360000;
#10;x=19370000;
#10;x=19380000;
#10;x=19390000;
#10;x=19400000;
#10;x=19410000;
#10;x=19420000;
#10;x=19430000;
#10;x=19440000;
#10;x=19450000;
#10;x=19460000;
#10;x=19470000;
#10;x=19480000;
#10;x=19490000;
#10;x=19500000;
#10;x=19510000;
#10;x=19520000;
#10;x=19530000;
#10;x=19540000;
#10;x=19550000;
#10;x=19560000;
#10;x=19570000;
#10;x=19580000;
#10;x=19590000;
#10;x=19600000;
#10;x=19610000;
#10;x=19620000;
#10;x=19630000;
#10;x=19640000;
#10;x=19650000;
#10;x=19660000;
#10;x=19670000;
#10;x=19680000;
#10;x=19690000;
#10;x=19700000;
#10;x=19710000;
#10;x=19720000;
#10;x=19730000;
#10;x=19740000;
#10;x=19750000;
#10;x=19760000;
#10;x=19770000;
#10;x=19780000;
#10;x=19790000;
#10;x=19800000;
#10;x=19810000;
#10;x=19820000;
#10;x=19830000;
#10;x=19840000;
#10;x=19850000;
#10;x=19860000;
#10;x=19870000;
#10;x=19880000;
#10;x=19890000;
#10;x=19900000;
#10;x=19910000;
#10;x=19920000;
#10;x=19930000;
#10;x=19940000;
#10;x=19950000;
#10;x=19960000;
#10;x=19970000;
#10;x=19980000;
#10;x=19990000;
#10;x=20000000;
#10;x=20010000;
#10;x=20020000;
#10;x=20030000;
#10;x=20040000;
#10;x=20050000;
#10;x=20060000;
#10;x=20070000;
#10;x=20080000;
#10;x=20090000;
#10;x=20100000;
#10;x=20110000;
#10;x=20120000;
#10;x=20130000;
#10;x=20140000;
#10;x=20150000;
#10;x=20160000;
#10;x=20170000;
#10;x=20180000;
#10;x=20190000;
#10;x=20200000;
#10;x=20210000;
#10;x=20220000;
#10;x=20230000;
#10;x=20240000;
#10;x=20250000;
#10;x=20260000;
#10;x=20270000;
#10;x=20280000;
#10;x=20290000;
#10;x=20300000;
#10;x=20310000;
#10;x=20320000;
#10;x=20330000;
#10;x=20340000;
#10;x=20350000;
#10;x=20360000;
#10;x=20370000;
#10;x=20380000;
#10;x=20390000;
#10;x=20400000;
#10;x=20410000;
#10;x=20420000;
#10;x=20430000;
#10;x=20440000;
#10;x=20450000;
#10;x=20460000;
#10;x=20470000;
#10;x=20480000;
#10;x=20490000;
#10;x=20500000;
#10;x=20510000;
#10;x=20520000;
#10;x=20530000;
#10;x=20540000;
#10;x=20550000;
#10;x=20560000;
#10;x=20570000;
#10;x=20580000;
#10;x=20590000;
#10;x=20600000;
#10;x=20610000;
#10;x=20620000;
#10;x=20630000;
#10;x=20640000;
#10;x=20650000;
#10;x=20660000;
#10;x=20670000;
#10;x=20680000;
#10;x=20690000;
#10;x=20700000;
#10;x=20710000;
#10;x=20720000;
#10;x=20730000;
#10;x=20740000;
#10;x=20750000;
#10;x=20760000;
#10;x=20770000;
#10;x=20780000;
#10;x=20790000;
#10;x=20800000;
#10;x=20810000;
#10;x=20820000;
#10;x=20830000;
#10;x=20840000;
#10;x=20850000;
#10;x=20860000;
#10;x=20870000;
#10;x=20880000;
#10;x=20890000;
#10;x=20900000;
#10;x=20910000;
#10;x=20920000;
#10;x=20930000;
#10;x=20940000;
#10;x=20950000;
#10;x=20960000;
#10;x=20970000;
#10;x=20980000;
#10;x=20990000;
#10;x=21000000;
#10;x=21010000;
#10;x=21020000;
#10;x=21030000;
#10;x=21040000;
#10;x=21050000;
#10;x=21060000;
#10;x=21070000;
#10;x=21080000;
#10;x=21090000;
#10;x=21100000;
#10;x=21110000;
#10;x=21120000;
#10;x=21130000;
#10;x=21140000;
#10;x=21150000;
#10;x=21160000;
#10;x=21170000;
#10;x=21180000;
#10;x=21190000;
#10;x=21200000;
#10;x=21210000;
#10;x=21220000;
#10;x=21230000;
#10;x=21240000;
#10;x=21250000;
#10;x=21260000;
#10;x=21270000;
#10;x=21280000;
#10;x=21290000;
#10;x=21300000;
#10;x=21310000;
#10;x=21320000;
#10;x=21330000;
#10;x=21340000;
#10;x=21350000;
#10;x=21360000;
#10;x=21370000;
#10;x=21380000;
#10;x=21390000;
#10;x=21400000;
#10;x=21410000;
#10;x=21420000;
#10;x=21430000;
#10;x=21440000;
#10;x=21450000;
#10;x=21460000;
#10;x=21470000;
#10;x=21480000;
#10;x=21490000;
#10;x=21500000;
#10;x=21510000;
#10;x=21520000;
#10;x=21530000;
#10;x=21540000;
#10;x=21550000;
#10;x=21560000;
#10;x=21570000;
#10;x=21580000;
#10;x=21590000;
#10;x=21600000;
#10;x=21610000;
#10;x=21620000;
#10;x=21630000;
#10;x=21640000;
#10;x=21650000;
#10;x=21660000;
#10;x=21670000;
#10;x=21680000;
#10;x=21690000;
#10;x=21700000;
#10;x=21710000;
#10;x=21720000;
#10;x=21730000;
#10;x=21740000;
#10;x=21750000;
#10;x=21760000;
#10;x=21770000;
#10;x=21780000;
#10;x=21790000;
#10;x=21800000;
#10;x=21810000;
#10;x=21820000;
#10;x=21830000;
#10;x=21840000;
#10;x=21850000;
#10;x=21860000;
#10;x=21870000;
#10;x=21880000;
#10;x=21890000;
#10;x=21900000;
#10;x=21910000;
#10;x=21920000;
#10;x=21930000;
#10;x=21940000;
#10;x=21950000;
#10;x=21960000;
#10;x=21970000;
#10;x=21980000;
#10;x=21990000;
#10;x=22000000;
#10;x=22010000;
#10;x=22020000;
#10;x=22030000;
#10;x=22040000;
#10;x=22050000;
#10;x=22060000;
#10;x=22070000;
#10;x=22080000;
#10;x=22090000;
#10;x=22100000;
#10;x=22110000;
#10;x=22120000;
#10;x=22130000;
#10;x=22140000;
#10;x=22150000;
#10;x=22160000;
#10;x=22170000;
#10;x=22180000;
#10;x=22190000;
#10;x=22200000;
#10;x=22210000;
#10;x=22220000;
#10;x=22230000;
#10;x=22240000;
#10;x=22250000;
#10;x=22260000;
#10;x=22270000;
#10;x=22280000;
#10;x=22290000;
#10;x=22300000;
#10;x=22310000;
#10;x=22320000;
#10;x=22330000;
#10;x=22340000;
#10;x=22350000;
#10;x=22360000;
#10;x=22370000;
#10;x=22380000;
#10;x=22390000;
#10;x=22400000;
#10;x=22410000;
#10;x=22420000;
#10;x=22430000;
#10;x=22440000;
#10;x=22450000;
#10;x=22460000;
#10;x=22470000;
#10;x=22480000;
#10;x=22490000;
#10;x=22500000;
#10;x=22510000;
#10;x=22520000;
#10;x=22530000;
#10;x=22540000;
#10;x=22550000;
#10;x=22560000;
#10;x=22570000;
#10;x=22580000;
#10;x=22590000;
#10;x=22600000;
#10;x=22610000;
#10;x=22620000;
#10;x=22630000;
#10;x=22640000;
#10;x=22650000;
#10;x=22660000;
#10;x=22670000;
#10;x=22680000;
#10;x=22690000;
#10;x=22700000;
#10;x=22710000;
#10;x=22720000;
#10;x=22730000;
#10;x=22740000;
#10;x=22750000;
#10;x=22760000;
#10;x=22770000;
#10;x=22780000;
#10;x=22790000;
#10;x=22800000;
#10;x=22810000;
#10;x=22820000;
#10;x=22830000;
#10;x=22840000;
#10;x=22850000;
#10;x=22860000;
#10;x=22870000;
#10;x=22880000;
#10;x=22890000;
#10;x=22900000;
#10;x=22910000;
#10;x=22920000;
#10;x=22930000;
#10;x=22940000;
#10;x=22950000;
#10;x=22960000;
#10;x=22970000;
#10;x=22980000;
#10;x=22990000;
#10;x=23000000;
#10;x=23010000;
#10;x=23020000;
#10;x=23030000;
#10;x=23040000;
#10;x=23050000;
#10;x=23060000;
#10;x=23070000;
#10;x=23080000;
#10;x=23090000;
#10;x=23100000;
#10;x=23110000;
#10;x=23120000;
#10;x=23130000;
#10;x=23140000;
#10;x=23150000;
#10;x=23160000;
#10;x=23170000;
#10;x=23180000;
#10;x=23190000;
#10;x=23200000;
#10;x=23210000;
#10;x=23220000;
#10;x=23230000;
#10;x=23240000;
#10;x=23250000;
#10;x=23260000;
#10;x=23270000;
#10;x=23280000;
#10;x=23290000;
#10;x=23300000;
#10;x=23310000;
#10;x=23320000;
#10;x=23330000;
#10;x=23340000;
#10;x=23350000;
#10;x=23360000;
#10;x=23370000;
#10;x=23380000;
#10;x=23390000;
#10;x=23400000;
#10;x=23410000;
#10;x=23420000;
#10;x=23430000;
#10;x=23440000;
#10;x=23450000;
#10;x=23460000;
#10;x=23470000;
#10;x=23480000;
#10;x=23490000;
#10;x=23500000;
#10;x=23510000;
#10;x=23520000;
#10;x=23530000;
#10;x=23540000;
#10;x=23550000;
#10;x=23560000;
#10;x=23570000;
#10;x=23580000;
#10;x=23590000;
#10;x=23600000;
#10;x=23610000;
#10;x=23620000;
#10;x=23630000;
#10;x=23640000;
#10;x=23650000;
#10;x=23660000;
#10;x=23670000;
#10;x=23680000;
#10;x=23690000;
#10;x=23700000;
#10;x=23710000;
#10;x=23720000;
#10;x=23730000;
#10;x=23740000;
#10;x=23750000;
#10;x=23760000;
#10;x=23770000;
#10;x=23780000;
#10;x=23790000;
#10;x=23800000;
#10;x=23810000;
#10;x=23820000;
#10;x=23830000;
#10;x=23840000;
#10;x=23850000;
#10;x=23860000;
#10;x=23870000;
#10;x=23880000;
#10;x=23890000;
#10;x=23900000;
#10;x=23910000;
#10;x=23920000;
#10;x=23930000;
#10;x=23940000;
#10;x=23950000;
#10;x=23960000;
#10;x=23970000;
#10;x=23980000;
#10;x=23990000;
#10;x=24000000;
#10;x=24010000;
#10;x=24020000;
#10;x=24030000;
#10;x=24040000;
#10;x=24050000;
#10;x=24060000;
#10;x=24070000;
#10;x=24080000;
#10;x=24090000;
#10;x=24100000;
#10;x=24110000;
#10;x=24120000;
#10;x=24130000;
#10;x=24140000;
#10;x=24150000;
#10;x=24160000;
#10;x=24170000;
#10;x=24180000;
#10;x=24190000;
#10;x=24200000;
#10;x=24210000;
#10;x=24220000;
#10;x=24230000;
#10;x=24240000;
#10;x=24250000;
#10;x=24260000;
#10;x=24270000;
#10;x=24280000;
#10;x=24290000;
#10;x=24300000;
#10;x=24310000;
#10;x=24320000;
#10;x=24330000;
#10;x=24340000;
#10;x=24350000;
#10;x=24360000;
#10;x=24370000;
#10;x=24380000;
#10;x=24390000;
#10;x=24400000;
#10;x=24410000;
#10;x=24420000;
#10;x=24430000;
#10;x=24440000;
#10;x=24450000;
#10;x=24460000;
#10;x=24470000;
#10;x=24480000;
#10;x=24490000;
#10;x=24500000;
#10;x=24510000;
#10;x=24520000;
#10;x=24530000;
#10;x=24540000;
#10;x=24550000;
#10;x=24560000;
#10;x=24570000;
#10;x=24580000;
#10;x=24590000;
#10;x=24600000;
#10;x=24610000;
#10;x=24620000;
#10;x=24630000;
#10;x=24640000;
#10;x=24650000;
#10;x=24660000;
#10;x=24670000;
#10;x=24680000;
#10;x=24690000;
#10;x=24700000;
#10;x=24710000;
#10;x=24720000;
#10;x=24730000;
#10;x=24740000;
#10;x=24750000;
#10;x=24760000;
#10;x=24770000;
#10;x=24780000;
#10;x=24790000;
#10;x=24800000;
#10;x=24810000;
#10;x=24820000;
#10;x=24830000;
#10;x=24840000;
#10;x=24850000;
#10;x=24860000;
#10;x=24870000;
#10;x=24880000;
#10;x=24890000;
#10;x=24900000;
#10;x=24910000;
#10;x=24920000;
#10;x=24930000;
#10;x=24940000;
#10;x=24950000;
#10;x=24960000;
#10;x=24970000;
#10;x=24980000;
#10;x=24990000;
#10;x=25000000;
#10;x=25010000;
#10;x=25020000;
#10;x=25030000;
#10;x=25040000;
#10;x=25050000;
#10;x=25060000;
#10;x=25070000;
#10;x=25080000;
#10;x=25090000;
#10;x=25100000;
#10;x=25110000;
#10;x=25120000;
#10;x=25130000;
#10;x=25140000;
#10;x=25150000;
#10;x=25160000;
#10;x=25170000;
#10;x=25180000;
#10;x=25190000;
#10;x=25200000;
#10;x=25210000;
#10;x=25220000;
#10;x=25230000;
#10;x=25240000;
#10;x=25250000;
#10;x=25260000;
#10;x=25270000;
#10;x=25280000;
#10;x=25290000;
#10;x=25300000;
#10;x=25310000;
#10;x=25320000;
#10;x=25330000;
#10;x=25340000;
#10;x=25350000;
#10;x=25360000;
#10;x=25370000;
#10;x=25380000;
#10;x=25390000;
#10;x=25400000;
#10;x=25410000;
#10;x=25420000;
#10;x=25430000;
#10;x=25440000;
#10;x=25450000;
#10;x=25460000;
#10;x=25470000;
#10;x=25480000;
#10;x=25490000;
#10;x=25500000;
#10;x=25510000;
#10;x=25520000;
#10;x=25530000;
#10;x=25540000;
#10;x=25550000;
#10;x=25560000;
#10;x=25570000;
#10;x=25580000;
#10;x=25590000;
#10;x=25600000;
#10;x=25610000;
#10;x=25620000;
#10;x=25630000;
#10;x=25640000;
#10;x=25650000;
#10;x=25660000;
#10;x=25670000;
#10;x=25680000;
#10;x=25690000;
#10;x=25700000;
#10;x=25710000;
#10;x=25720000;
#10;x=25730000;
#10;x=25740000;
#10;x=25750000;
#10;x=25760000;
#10;x=25770000;
#10;x=25780000;
#10;x=25790000;
#10;x=25800000;
#10;x=25810000;
#10;x=25820000;
#10;x=25830000;
#10;x=25840000;
#10;x=25850000;
#10;x=25860000;
#10;x=25870000;
#10;x=25880000;
#10;x=25890000;
#10;x=25900000;
#10;x=25910000;
#10;x=25920000;
#10;x=25930000;
#10;x=25940000;
#10;x=25950000;
#10;x=25960000;
#10;x=25970000;
#10;x=25980000;
#10;x=25990000;
#10;x=26000000;
#10;x=26010000;
#10;x=26020000;
#10;x=26030000;
#10;x=26040000;
#10;x=26050000;
#10;x=26060000;
#10;x=26070000;
#10;x=26080000;
#10;x=26090000;
#10;x=26100000;
#10;x=26110000;
#10;x=26120000;
#10;x=26130000;
#10;x=26140000;
#10;x=26150000;
#10;x=26160000;
#10;x=26170000;
#10;x=26180000;
#10;x=26190000;
#10;x=26200000;
#10;x=26210000;
#10;x=26220000;
#10;x=26230000;
#10;x=26240000;
#10;x=26250000;
#10;x=26260000;
#10;x=26270000;
#10;x=26280000;
#10;x=26290000;
#10;x=26300000;
#10;x=26310000;
#10;x=26320000;
#10;x=26330000;
#10;x=26340000;
#10;x=26350000;
#10;x=26360000;
#10;x=26370000;
#10;x=26380000;
#10;x=26390000;
#10;x=26400000;
#10;x=26410000;
#10;x=26420000;
#10;x=26430000;
#10;x=26440000;
#10;x=26450000;
#10;x=26460000;
#10;x=26470000;
#10;x=26480000;
#10;x=26490000;
#10;x=26500000;
#10;x=26510000;
#10;x=26520000;
#10;x=26530000;
#10;x=26540000;
#10;x=26550000;
#10;x=26560000;
#10;x=26570000;
#10;x=26580000;
#10;x=26590000;
#10;x=26600000;
#10;x=26610000;
#10;x=26620000;
#10;x=26630000;
#10;x=26640000;
#10;x=26650000;
#10;x=26660000;
#10;x=26670000;
#10;x=26680000;
#10;x=26690000;
#10;x=26700000;
#10;x=26710000;
#10;x=26720000;
#10;x=26730000;
#10;x=26740000;
#10;x=26750000;
#10;x=26760000;
#10;x=26770000;
#10;x=26780000;
#10;x=26790000;
#10;x=26800000;
#10;x=26810000;
#10;x=26820000;
#10;x=26830000;
#10;x=26840000;
#10;x=26850000;
#10;x=26860000;
#10;x=26870000;
#10;x=26880000;
#10;x=26890000;
#10;x=26900000;
#10;x=26910000;
#10;x=26920000;
#10;x=26930000;
#10;x=26940000;
#10;x=26950000;
#10;x=26960000;
#10;x=26970000;
#10;x=26980000;
#10;x=26990000;
#10;x=27000000;
#10;x=27010000;
#10;x=27020000;
#10;x=27030000;
#10;x=27040000;
#10;x=27050000;
#10;x=27060000;
#10;x=27070000;
#10;x=27080000;
#10;x=27090000;
#10;x=27100000;
#10;x=27110000;
#10;x=27120000;
#10;x=27130000;
#10;x=27140000;
#10;x=27150000;
#10;x=27160000;
#10;x=27170000;
#10;x=27180000;
#10;x=27190000;
#10;x=27200000;
#10;x=27210000;
#10;x=27220000;
#10;x=27230000;
#10;x=27240000;
#10;x=27250000;
#10;x=27260000;
#10;x=27270000;
#10;x=27280000;
#10;x=27290000;
#10;x=27300000;
#10;x=27310000;
#10;x=27320000;
#10;x=27330000;
#10;x=27340000;
#10;x=27350000;
#10;x=27360000;
#10;x=27370000;
#10;x=27380000;
#10;x=27390000;
#10;x=27400000;
#10;x=27410000;
#10;x=27420000;
#10;x=27430000;
#10;x=27440000;
#10;x=27450000;
#10;x=27460000;
#10;x=27470000;
#10;x=27480000;
#10;x=27490000;
#10;x=27500000;
#10;x=27510000;
#10;x=27520000;
#10;x=27530000;
#10;x=27540000;
#10;x=27550000;
#10;x=27560000;
#10;x=27570000;
#10;x=27580000;
#10;x=27590000;
#10;x=27600000;
#10;x=27610000;
#10;x=27620000;
#10;x=27630000;
#10;x=27640000;
#10;x=27650000;
#10;x=27660000;
#10;x=27670000;
#10;x=27680000;
#10;x=27690000;
#10;x=27700000;
#10;x=27710000;
#10;x=27720000;
#10;x=27730000;
#10;x=27740000;
#10;x=27750000;
#10;x=27760000;
#10;x=27770000;
#10;x=27780000;
#10;x=27790000;
#10;x=27800000;
#10;x=27810000;
#10;x=27820000;
#10;x=27830000;
#10;x=27840000;
#10;x=27850000;
#10;x=27860000;
#10;x=27870000;
#10;x=27880000;
#10;x=27890000;
#10;x=27900000;
#10;x=27910000;
#10;x=27920000;
#10;x=27930000;
#10;x=27940000;
#10;x=27950000;
#10;x=27960000;
#10;x=27970000;
#10;x=27980000;
#10;x=27990000;
#10;x=28000000;
#10;x=28010000;
#10;x=28020000;
#10;x=28030000;
#10;x=28040000;
#10;x=28050000;
#10;x=28060000;
#10;x=28070000;
#10;x=28080000;
#10;x=28090000;
#10;x=28100000;
#10;x=28110000;
#10;x=28120000;
#10;x=28130000;
#10;x=28140000;
#10;x=28150000;
#10;x=28160000;
#10;x=28170000;
#10;x=28180000;
#10;x=28190000;
#10;x=28200000;
#10;x=28210000;
#10;x=28220000;
#10;x=28230000;
#10;x=28240000;
#10;x=28250000;
#10;x=28260000;
#10;x=28270000;
#10;x=28280000;
#10;x=28290000;
#10;x=28300000;
#10;x=28310000;
#10;x=28320000;
#10;x=28330000;
#10;x=28340000;
#10;x=28350000;
#10;x=28360000;
#10;x=28370000;
#10;x=28380000;
#10;x=28390000;
#10;x=28400000;
#10;x=28410000;
#10;x=28420000;
#10;x=28430000;
#10;x=28440000;
#10;x=28450000;
#10;x=28460000;
#10;x=28470000;
#10;x=28480000;
#10;x=28490000;
#10;x=28500000;
#10;x=28510000;
#10;x=28520000;
#10;x=28530000;
#10;x=28540000;
#10;x=28550000;
#10;x=28560000;
#10;x=28570000;
#10;x=28580000;
#10;x=28590000;
#10;x=28600000;
#10;x=28610000;
#10;x=28620000;
#10;x=28630000;
#10;x=28640000;
#10;x=28650000;
#10;x=28660000;
#10;x=28670000;
#10;x=28680000;
#10;x=28690000;
#10;x=28700000;
#10;x=28710000;
#10;x=28720000;
#10;x=28730000;
#10;x=28740000;
#10;x=28750000;
#10;x=28760000;
#10;x=28770000;
#10;x=28780000;
#10;x=28790000;
#10;x=28800000;
#10;x=28810000;
#10;x=28820000;
#10;x=28830000;
#10;x=28840000;
#10;x=28850000;
#10;x=28860000;
#10;x=28870000;
#10;x=28880000;
#10;x=28890000;
#10;x=28900000;
#10;x=28910000;
#10;x=28920000;
#10;x=28930000;
#10;x=28940000;
#10;x=28950000;
#10;x=28960000;
#10;x=28970000;
#10;x=28980000;
#10;x=28990000;
#10;x=29000000;
#10;x=29010000;
#10;x=29020000;
#10;x=29030000;
#10;x=29040000;
#10;x=29050000;
#10;x=29060000;
#10;x=29070000;
#10;x=29080000;
#10;x=29090000;
#10;x=29100000;
#10;x=29110000;
#10;x=29120000;
#10;x=29130000;
#10;x=29140000;
#10;x=29150000;
#10;x=29160000;
#10;x=29170000;
#10;x=29180000;
#10;x=29190000;
#10;x=29200000;
#10;x=29210000;
#10;x=29220000;
#10;x=29230000;
#10;x=29240000;
#10;x=29250000;
#10;x=29260000;
#10;x=29270000;
#10;x=29280000;
#10;x=29290000;
#10;x=29300000;
#10;x=29310000;
#10;x=29320000;
#10;x=29330000;
#10;x=29340000;
#10;x=29350000;
#10;x=29360000;
#10;x=29370000;
#10;x=29380000;
#10;x=29390000;
#10;x=29400000;
#10;x=29410000;
#10;x=29420000;
#10;x=29430000;
#10;x=29440000;
#10;x=29450000;
#10;x=29460000;
#10;x=29470000;
#10;x=29480000;
#10;x=29490000;
#10;x=29500000;
#10;x=29510000;
#10;x=29520000;
#10;x=29530000;
#10;x=29540000;
#10;x=29550000;
#10;x=29560000;
#10;x=29570000;
#10;x=29580000;
#10;x=29590000;
#10;x=29600000;
#10;x=29610000;
#10;x=29620000;
#10;x=29630000;
#10;x=29640000;
#10;x=29650000;
#10;x=29660000;
#10;x=29670000;
#10;x=29680000;
#10;x=29690000;
#10;x=29700000;
#10;x=29710000;
#10;x=29720000;
#10;x=29730000;
#10;x=29740000;
#10;x=29750000;
#10;x=29760000;
#10;x=29770000;
#10;x=29780000;
#10;x=29790000;
#10;x=29800000;
#10;x=29810000;
#10;x=29820000;
#10;x=29830000;
#10;x=29840000;
#10;x=29850000;
#10;x=29860000;
#10;x=29870000;
#10;x=29880000;
#10;x=29890000;
#10;x=29900000;
#10;x=29910000;
#10;x=29920000;
#10;x=29930000;
#10;x=29940000;
#10;x=29950000;
#10;x=29960000;
#10;x=29970000;
#10;x=29980000;
#10;x=29990000;
#10;x=30000000;
#10;x=30010000;
#10;x=30020000;
#10;x=30030000;
#10;x=30040000;
#10;x=30050000;
#10;x=30060000;
#10;x=30070000;
#10;x=30080000;
#10;x=30090000;
#10;x=30100000;
#10;x=30110000;
#10;x=30120000;
#10;x=30130000;
#10;x=30140000;
#10;x=30150000;
#10;x=30160000;
#10;x=30170000;
#10;x=30180000;
#10;x=30190000;
#10;x=30200000;
#10;x=30210000;
#10;x=30220000;
#10;x=30230000;
#10;x=30240000;
#10;x=30250000;
#10;x=30260000;
#10;x=30270000;
#10;x=30280000;
#10;x=30290000;
#10;x=30300000;
#10;x=30310000;
#10;x=30320000;
#10;x=30330000;
#10;x=30340000;
#10;x=30350000;
#10;x=30360000;
#10;x=30370000;
#10;x=30380000;
#10;x=30390000;
#10;x=30400000;
#10;x=30410000;
#10;x=30420000;
#10;x=30430000;
#10;x=30440000;
#10;x=30450000;
#10;x=30460000;
#10;x=30470000;
#10;x=30480000;
#10;x=30490000;
#10;x=30500000;
#10;x=30510000;
#10;x=30520000;
#10;x=30530000;
#10;x=30540000;
#10;x=30550000;
#10;x=30560000;
#10;x=30570000;
#10;x=30580000;
#10;x=30590000;
#10;x=30600000;
#10;x=30610000;
#10;x=30620000;
#10;x=30630000;
#10;x=30640000;
#10;x=30650000;
#10;x=30660000;
#10;x=30670000;
#10;x=30680000;
#10;x=30690000;
#10;x=30700000;
#10;x=30710000;
#10;x=30720000;
#10;x=30730000;
#10;x=30740000;
#10;x=30750000;
#10;x=30760000;
#10;x=30770000;
#10;x=30780000;
#10;x=30790000;
#10;x=30800000;
#10;x=30810000;
#10;x=30820000;
#10;x=30830000;
#10;x=30840000;
#10;x=30850000;
#10;x=30860000;
#10;x=30870000;
#10;x=30880000;
#10;x=30890000;
#10;x=30900000;
#10;x=30910000;
#10;x=30920000;
#10;x=30930000;
#10;x=30940000;
#10;x=30950000;
#10;x=30960000;
#10;x=30970000;
#10;x=30980000;
#10;x=30990000;
#10;x=31000000;
#10;x=31010000;
#10;x=31020000;
#10;x=31030000;
#10;x=31040000;
#10;x=31050000;
#10;x=31060000;
#10;x=31070000;
#10;x=31080000;
#10;x=31090000;
#10;x=31100000;
#10;x=31110000;
#10;x=31120000;
#10;x=31130000;
#10;x=31140000;
#10;x=31150000;
#10;x=31160000;
#10;x=31170000;
#10;x=31180000;
#10;x=31190000;
#10;x=31200000;
#10;x=31210000;
#10;x=31220000;
#10;x=31230000;
#10;x=31240000;
#10;x=31250000;
#10;x=31260000;
#10;x=31270000;
#10;x=31280000;
#10;x=31290000;
#10;x=31300000;
#10;x=31310000;
#10;x=31320000;
#10;x=31330000;
#10;x=31340000;
#10;x=31350000;
#10;x=31360000;
#10;x=31370000;
#10;x=31380000;
#10;x=31390000;
#10;x=31400000;
#10;x=31410000;
#10;x=31420000;
#10;x=31430000;
#10;x=31440000;
#10;x=31450000;
#10;x=31460000;
#10;x=31470000;
#10;x=31480000;
#10;x=31490000;
#10;x=31500000;
#10;x=31510000;
#10;x=31520000;
#10;x=31530000;
#10;x=31540000;
#10;x=31550000;
#10;x=31560000;
#10;x=31570000;
#10;x=31580000;
#10;x=31590000;
#10;x=31600000;
#10;x=31610000;
#10;x=31620000;
#10;x=31630000;
#10;x=31640000;
#10;x=31650000;
#10;x=31660000;
#10;x=31670000;
#10;x=31680000;
#10;x=31690000;
#10;x=31700000;
#10;x=31710000;
#10;x=31720000;
#10;x=31730000;
#10;x=31740000;
#10;x=31750000;
#10;x=31760000;
#10;x=31770000;
#10;x=31780000;
#10;x=31790000;
#10;x=31800000;
#10;x=31810000;
#10;x=31820000;
#10;x=31830000;
#10;x=31840000;
#10;x=31850000;
#10;x=31860000;
#10;x=31870000;
#10;x=31880000;
#10;x=31890000;
#10;x=31900000;
#10;x=31910000;
#10;x=31920000;
#10;x=31930000;
#10;x=31940000;
#10;x=31950000;
#10;x=31960000;
#10;x=31970000;
#10;x=31980000;
#10;x=31990000;
#10;x=32000000;
#10;x=32010000;
#10;x=32020000;
#10;x=32030000;
#10;x=32040000;
#10;x=32050000;
#10;x=32060000;
#10;x=32070000;
#10;x=32080000;
#10;x=32090000;
#10;x=32100000;
#10;x=32110000;
#10;x=32120000;
#10;x=32130000;
#10;x=32140000;
#10;x=32150000;
#10;x=32160000;
#10;x=32170000;
#10;x=32180000;
#10;x=32190000;
#10;x=32200000;
#10;x=32210000;
#10;x=32220000;
#10;x=32230000;
#10;x=32240000;
#10;x=32250000;
#10;x=32260000;
#10;x=32270000;
#10;x=32280000;
#10;x=32290000;
#10;x=32300000;
#10;x=32310000;
#10;x=32320000;
#10;x=32330000;
#10;x=32340000;
#10;x=32350000;
#10;x=32360000;
#10;x=32370000;
#10;x=32380000;
#10;x=32390000;
#10;x=32400000;
#10;x=32410000;
#10;x=32420000;
#10;x=32430000;
#10;x=32440000;
#10;x=32450000;
#10;x=32460000;
#10;x=32470000;
#10;x=32480000;
#10;x=32490000;
#10;x=32500000;
#10;x=32510000;
#10;x=32520000;
#10;x=32530000;
#10;x=32540000;
#10;x=32550000;
#10;x=32560000;
#10;x=32570000;
#10;x=32580000;
#10;x=32590000;
#10;x=32600000;
#10;x=32610000;
#10;x=32620000;
#10;x=32630000;
#10;x=32640000;
#10;x=32650000;
#10;x=32660000;
#10;x=32670000;
#10;x=32680000;
#10;x=32690000;
#10;x=32700000;
#10;x=32710000;
#10;x=32720000;
#10;x=32730000;
#10;x=32740000;
#10;x=32750000;
#10;x=32760000;
#10;x=32770000;
#10;x=32780000;
#10;x=32790000;
#10;x=32800000;
#10;x=32810000;
#10;x=32820000;
#10;x=32830000;
#10;x=32840000;
#10;x=32850000;
#10;x=32860000;
#10;x=32870000;
#10;x=32880000;
#10;x=32890000;
#10;x=32900000;
#10;x=32910000;
#10;x=32920000;
#10;x=32930000;
#10;x=32940000;
#10;x=32950000;
#10;x=32960000;
#10;x=32970000;
#10;x=32980000;
#10;x=32990000;
#10;x=33000000;
#10;x=33010000;
#10;x=33020000;
#10;x=33030000;
#10;x=33040000;
#10;x=33050000;
#10;x=33060000;
#10;x=33070000;
#10;x=33080000;
#10;x=33090000;
#10;x=33100000;
#10;x=33110000;
#10;x=33120000;
#10;x=33130000;
#10;x=33140000;
#10;x=33150000;
#10;x=33160000;
#10;x=33170000;
#10;x=33180000;
#10;x=33190000;
#10;x=33200000;
#10;x=33210000;
#10;x=33220000;
#10;x=33230000;
#10;x=33240000;
#10;x=33250000;
#10;x=33260000;
#10;x=33270000;
#10;x=33280000;
#10;x=33290000;
#10;x=33300000;
#10;x=33310000;
#10;x=33320000;
#10;x=33330000;
#10;x=33340000;
#10;x=33350000;
#10;x=33360000;
#10;x=33370000;
#10;x=33380000;
#10;x=33390000;
#10;x=33400000;
#10;x=33410000;
#10;x=33420000;
#10;x=33430000;
#10;x=33440000;
#10;x=33450000;
#10;x=33460000;
#10;x=33470000;
#10;x=33480000;
#10;x=33490000;
#10;x=33500000;
#10;x=33510000;
#10;x=33520000;
#10;x=33530000;
#10;x=33540000;
#10;x=33550000;
#10;x=33560000;
#10;x=33570000;
#10;x=33580000;
#10;x=33590000;
#10;x=33600000;
#10;x=33610000;
#10;x=33620000;
#10;x=33630000;
#10;x=33640000;
#10;x=33650000;
#10;x=33660000;
#10;x=33670000;
#10;x=33680000;
#10;x=33690000;
#10;x=33700000;
#10;x=33710000;
#10;x=33720000;
#10;x=33730000;
#10;x=33740000;
#10;x=33750000;
#10;x=33760000;
#10;x=33770000;
#10;x=33780000;
#10;x=33790000;
#10;x=33800000;
#10;x=33810000;
#10;x=33820000;
#10;x=33830000;
#10;x=33840000;
#10;x=33850000;
#10;x=33860000;
#10;x=33870000;
#10;x=33880000;
#10;x=33890000;
#10;x=33900000;
#10;x=33910000;
#10;x=33920000;
#10;x=33930000;
#10;x=33940000;
#10;x=33950000;
#10;x=33960000;
#10;x=33970000;
#10;x=33980000;
#10;x=33990000;
#10;x=34000000;
#10;x=34010000;
#10;x=34020000;
#10;x=34030000;
#10;x=34040000;
#10;x=34050000;
#10;x=34060000;
#10;x=34070000;
#10;x=34080000;
#10;x=34090000;
#10;x=34100000;
#10;x=34110000;
#10;x=34120000;
#10;x=34130000;
#10;x=34140000;
#10;x=34150000;
#10;x=34160000;
#10;x=34170000;
#10;x=34180000;
#10;x=34190000;
#10;x=34200000;
#10;x=34210000;
#10;x=34220000;
#10;x=34230000;
#10;x=34240000;
#10;x=34250000;
#10;x=34260000;
#10;x=34270000;
#10;x=34280000;
#10;x=34290000;
#10;x=34300000;
#10;x=34310000;
#10;x=34320000;
#10;x=34330000;
#10;x=34340000;
#10;x=34350000;
#10;x=34360000;
#10;x=34370000;
#10;x=34380000;
#10;x=34390000;
#10;x=34400000;
#10;x=34410000;
#10;x=34420000;
#10;x=34430000;
#10;x=34440000;
#10;x=34450000;
#10;x=34460000;
#10;x=34470000;
#10;x=34480000;
#10;x=34490000;
#10;x=34500000;
#10;x=34510000;
#10;x=34520000;
#10;x=34530000;
#10;x=34540000;
#10;x=34550000;
#10;x=34560000;
#10;x=34570000;
#10;x=34580000;
#10;x=34590000;
#10;x=34600000;
#10;x=34610000;
#10;x=34620000;
#10;x=34630000;
#10;x=34640000;
#10;x=34650000;
#10;x=34660000;
#10;x=34670000;
#10;x=34680000;
#10;x=34690000;
#10;x=34700000;
#10;x=34710000;
#10;x=34720000;
#10;x=34730000;
#10;x=34740000;
#10;x=34750000;
#10;x=34760000;
#10;x=34770000;
#10;x=34780000;
#10;x=34790000;
#10;x=34800000;
#10;x=34810000;
#10;x=34820000;
#10;x=34830000;
#10;x=34840000;
#10;x=34850000;
#10;x=34860000;
#10;x=34870000;
#10;x=34880000;
#10;x=34890000;
#10;x=34900000;
#10;x=34910000;
#10;x=34920000;
#10;x=34930000;
#10;x=34940000;
#10;x=34950000;
#10;x=34960000;
#10;x=34970000;
#10;x=34980000;
#10;x=34990000;
#10;x=35000000;
#10;x=35010000;
#10;x=35020000;
#10;x=35030000;
#10;x=35040000;
#10;x=35050000;
#10;x=35060000;
#10;x=35070000;
#10;x=35080000;
#10;x=35090000;
#10;x=35100000;
#10;x=35110000;
#10;x=35120000;
#10;x=35130000;
#10;x=35140000;
#10;x=35150000;
#10;x=35160000;
#10;x=35170000;
#10;x=35180000;
#10;x=35190000;
#10;x=35200000;
#10;x=35210000;
#10;x=35220000;
#10;x=35230000;
#10;x=35240000;
#10;x=35250000;
#10;x=35260000;
#10;x=35270000;
#10;x=35280000;
#10;x=35290000;
#10;x=35300000;
#10;x=35310000;
#10;x=35320000;
#10;x=35330000;
#10;x=35340000;
#10;x=35350000;
#10;x=35360000;
#10;x=35370000;
#10;x=35380000;
#10;x=35390000;
#10;x=35400000;
#10;x=35410000;
#10;x=35420000;
#10;x=35430000;
#10;x=35440000;
#10;x=35450000;
#10;x=35460000;
#10;x=35470000;
#10;x=35480000;
#10;x=35490000;
#10;x=35500000;
#10;x=35510000;
#10;x=35520000;
#10;x=35530000;
#10;x=35540000;
#10;x=35550000;
#10;x=35560000;
#10;x=35570000;
#10;x=35580000;
#10;x=35590000;
#10;x=35600000;
#10;x=35610000;
#10;x=35620000;
#10;x=35630000;
#10;x=35640000;
#10;x=35650000;
#10;x=35660000;
#10;x=35670000;
#10;x=35680000;
#10;x=35690000;
#10;x=35700000;
#10;x=35710000;
#10;x=35720000;
#10;x=35730000;
#10;x=35740000;
#10;x=35750000;
#10;x=35760000;
#10;x=35770000;
#10;x=35780000;
#10;x=35790000;
#10;x=35800000;
#10;x=35810000;
#10;x=35820000;
#10;x=35830000;
#10;x=35840000;
#10;x=35850000;
#10;x=35860000;
#10;x=35870000;
#10;x=35880000;
#10;x=35890000;
#10;x=35900000;
#10;x=35910000;
#10;x=35920000;
#10;x=35930000;
#10;x=35940000;
#10;x=35950000;
#10;x=35960000;
#10;x=35970000;
#10;x=35980000;
#10;x=35990000;
#10;x=36000000;
#10;x=36010000;
#10;x=36020000;
#10;x=36030000;
#10;x=36040000;
#10;x=36050000;
#10;x=36060000;
#10;x=36070000;
#10;x=36080000;
#10;x=36090000;
#10;x=36100000;
#10;x=36110000;
#10;x=36120000;
#10;x=36130000;
#10;x=36140000;
#10;x=36150000;
#10;x=36160000;
#10;x=36170000;
#10;x=36180000;
#10;x=36190000;
#10;x=36200000;
#10;x=36210000;
#10;x=36220000;
#10;x=36230000;
#10;x=36240000;
#10;x=36250000;
#10;x=36260000;
#10;x=36270000;
#10;x=36280000;
#10;x=36290000;
#10;x=36300000;
#10;x=36310000;
#10;x=36320000;
#10;x=36330000;
#10;x=36340000;
#10;x=36350000;
#10;x=36360000;
#10;x=36370000;
#10;x=36380000;
#10;x=36390000;
#10;x=36400000;
#10;x=36410000;
#10;x=36420000;
#10;x=36430000;
#10;x=36440000;
#10;x=36450000;
#10;x=36460000;
#10;x=36470000;
#10;x=36480000;
#10;x=36490000;
#10;x=36500000;
#10;x=36510000;
#10;x=36520000;
#10;x=36530000;
#10;x=36540000;
#10;x=36550000;
#10;x=36560000;
#10;x=36570000;
#10;x=36580000;
#10;x=36590000;
#10;x=36600000;
#10;x=36610000;
#10;x=36620000;
#10;x=36630000;
#10;x=36640000;
#10;x=36650000;
#10;x=36660000;
#10;x=36670000;
#10;x=36680000;
#10;x=36690000;
#10;x=36700000;
#10;x=36710000;
#10;x=36720000;
#10;x=36730000;
#10;x=36740000;
#10;x=36750000;
#10;x=36760000;
#10;x=36770000;
#10;x=36780000;
#10;x=36790000;
#10;x=36800000;
#10;x=36810000;
#10;x=36820000;
#10;x=36830000;
#10;x=36840000;
#10;x=36850000;
#10;x=36860000;
#10;x=36870000;
#10;x=36880000;
#10;x=36890000;
#10;x=36900000;
#10;x=36910000;
#10;x=36920000;
#10;x=36930000;
#10;x=36940000;
#10;x=36950000;
#10;x=36960000;
#10;x=36970000;
#10;x=36980000;
#10;x=36990000;
#10;x=37000000;
#10;x=37010000;
#10;x=37020000;
#10;x=37030000;
#10;x=37040000;
#10;x=37050000;
#10;x=37060000;
#10;x=37070000;
#10;x=37080000;
#10;x=37090000;
#10;x=37100000;
#10;x=37110000;
#10;x=37120000;
#10;x=37130000;
#10;x=37140000;
#10;x=37150000;
#10;x=37160000;
#10;x=37170000;
#10;x=37180000;
#10;x=37190000;
#10;x=37200000;
#10;x=37210000;
#10;x=37220000;
#10;x=37230000;
#10;x=37240000;
#10;x=37250000;
#10;x=37260000;
#10;x=37270000;
#10;x=37280000;
#10;x=37290000;
#10;x=37300000;
#10;x=37310000;
#10;x=37320000;
#10;x=37330000;
#10;x=37340000;
#10;x=37350000;
#10;x=37360000;
#10;x=37370000;
#10;x=37380000;
#10;x=37390000;
#10;x=37400000;
#10;x=37410000;
#10;x=37420000;
#10;x=37430000;
#10;x=37440000;
#10;x=37450000;
#10;x=37460000;
#10;x=37470000;
#10;x=37480000;
#10;x=37490000;
#10;x=37500000;
#10;x=37510000;
#10;x=37520000;
#10;x=37530000;
#10;x=37540000;
#10;x=37550000;
#10;x=37560000;
#10;x=37570000;
#10;x=37580000;
#10;x=37590000;
#10;x=37600000;
#10;x=37610000;
#10;x=37620000;
#10;x=37630000;
#10;x=37640000;
#10;x=37650000;
#10;x=37660000;
#10;x=37670000;
#10;x=37680000;
#10;x=37690000;
#10;x=37700000;
#10;x=37710000;
#10;x=37720000;
#10;x=37730000;
#10;x=37740000;
#10;x=37750000;
#10;x=37760000;
#10;x=37770000;
#10;x=37780000;
#10;x=37790000;
#10;x=37800000;
#10;x=37810000;
#10;x=37820000;
#10;x=37830000;
#10;x=37840000;
#10;x=37850000;
#10;x=37860000;
#10;x=37870000;
#10;x=37880000;
#10;x=37890000;
#10;x=37900000;
#10;x=37910000;
#10;x=37920000;
#10;x=37930000;
#10;x=37940000;
#10;x=37950000;
#10;x=37960000;
#10;x=37970000;
#10;x=37980000;
#10;x=37990000;
#10;x=38000000;
#10;x=38010000;
#10;x=38020000;
#10;x=38030000;
#10;x=38040000;
#10;x=38050000;
#10;x=38060000;
#10;x=38070000;
#10;x=38080000;
#10;x=38090000;
#10;x=38100000;
#10;x=38110000;
#10;x=38120000;
#10;x=38130000;
#10;x=38140000;
#10;x=38150000;
#10;x=38160000;
#10;x=38170000;
#10;x=38180000;
#10;x=38190000;
#10;x=38200000;
#10;x=38210000;
#10;x=38220000;
#10;x=38230000;
#10;x=38240000;
#10;x=38250000;
#10;x=38260000;
#10;x=38270000;
#10;x=38280000;
#10;x=38290000;
#10;x=38300000;
#10;x=38310000;
#10;x=38320000;
#10;x=38330000;
#10;x=38340000;
#10;x=38350000;
#10;x=38360000;
#10;x=38370000;
#10;x=38380000;
#10;x=38390000;
#10;x=38400000;
#10;x=38410000;
#10;x=38420000;
#10;x=38430000;
#10;x=38440000;
#10;x=38450000;
#10;x=38460000;
#10;x=38470000;
#10;x=38480000;
#10;x=38490000;
#10;x=38500000;
#10;x=38510000;
#10;x=38520000;
#10;x=38530000;
#10;x=38540000;
#10;x=38550000;
#10;x=38560000;
#10;x=38570000;
#10;x=38580000;
#10;x=38590000;
#10;x=38600000;
#10;x=38610000;
#10;x=38620000;
#10;x=38630000;
#10;x=38640000;
#10;x=38650000;
#10;x=38660000;
#10;x=38670000;
#10;x=38680000;
#10;x=38690000;
#10;x=38700000;
#10;x=38710000;
#10;x=38720000;
#10;x=38730000;
#10;x=38740000;
#10;x=38750000;
#10;x=38760000;
#10;x=38770000;
#10;x=38780000;
#10;x=38790000;
#10;x=38800000;
#10;x=38810000;
#10;x=38820000;
#10;x=38830000;
#10;x=38840000;
#10;x=38850000;
#10;x=38860000;
#10;x=38870000;
#10;x=38880000;
#10;x=38890000;
#10;x=38900000;
#10;x=38910000;
#10;x=38920000;
#10;x=38930000;
#10;x=38940000;
#10;x=38950000;
#10;x=38960000;
#10;x=38970000;
#10;x=38980000;
#10;x=38990000;
#10;x=39000000;
#10;x=39010000;
#10;x=39020000;
#10;x=39030000;
#10;x=39040000;
#10;x=39050000;
#10;x=39060000;
#10;x=39070000;
#10;x=39080000;
#10;x=39090000;
#10;x=39100000;
#10;x=39110000;
#10;x=39120000;
#10;x=39130000;
#10;x=39140000;
#10;x=39150000;
#10;x=39160000;
#10;x=39170000;
#10;x=39180000;
#10;x=39190000;
#10;x=39200000;
#10;x=39210000;
#10;x=39220000;
#10;x=39230000;
#10;x=39240000;
#10;x=39250000;
#10;x=39260000;
#10;x=39270000;
#10;x=39280000;
#10;x=39290000;
#10;x=39300000;
#10;x=39310000;
#10;x=39320000;
#10;x=39330000;
#10;x=39340000;
#10;x=39350000;
#10;x=39360000;
#10;x=39370000;
#10;x=39380000;
#10;x=39390000;
#10;x=39400000;
#10;x=39410000;
#10;x=39420000;
#10;x=39430000;
#10;x=39440000;
#10;x=39450000;
#10;x=39460000;
#10;x=39470000;
#10;x=39480000;
#10;x=39490000;
#10;x=39500000;
#10;x=39510000;
#10;x=39520000;
#10;x=39530000;
#10;x=39540000;
#10;x=39550000;
#10;x=39560000;
#10;x=39570000;
#10;x=39580000;
#10;x=39590000;
#10;x=39600000;
#10;x=39610000;
#10;x=39620000;
#10;x=39630000;
#10;x=39640000;
#10;x=39650000;
#10;x=39660000;
#10;x=39670000;
#10;x=39680000;
#10;x=39690000;
#10;x=39700000;
#10;x=39710000;
#10;x=39720000;
#10;x=39730000;
#10;x=39740000;
#10;x=39750000;
#10;x=39760000;
#10;x=39770000;
#10;x=39780000;
#10;x=39790000;
#10;x=39800000;
#10;x=39810000;
#10;x=39820000;
#10;x=39830000;
#10;x=39840000;
#10;x=39850000;
#10;x=39860000;
#10;x=39870000;
#10;x=39880000;
#10;x=39890000;
#10;x=39900000;
#10;x=39910000;
#10;x=39920000;
#10;x=39930000;
#10;x=39940000;
#10;x=39950000;
#10;x=39960000;
#10;x=39970000;
#10;x=39980000;
#10;x=39990000;
#10;x=40000000;
#10;x=40010000;
#10;x=40020000;
#10;x=40030000;
#10;x=40040000;
#10;x=40050000;
#10;x=40060000;
#10;x=40070000;
#10;x=40080000;
#10;x=40090000;
#10;x=40100000;
#10;x=40110000;
#10;x=40120000;
#10;x=40130000;
#10;x=40140000;
#10;x=40150000;
#10;x=40160000;
#10;x=40170000;
#10;x=40180000;
#10;x=40190000;
#10;x=40200000;
#10;x=40210000;
#10;x=40220000;
#10;x=40230000;
#10;x=40240000;
#10;x=40250000;
#10;x=40260000;
#10;x=40270000;
#10;x=40280000;
#10;x=40290000;
#10;x=40300000;
#10;x=40310000;
#10;x=40320000;
#10;x=40330000;
#10;x=40340000;
#10;x=40350000;
#10;x=40360000;
#10;x=40370000;
#10;x=40380000;
#10;x=40390000;
#10;x=40400000;
#10;x=40410000;
#10;x=40420000;
#10;x=40430000;
#10;x=40440000;
#10;x=40450000;
#10;x=40460000;
#10;x=40470000;
#10;x=40480000;
#10;x=40490000;
#10;x=40500000;
#10;x=40510000;
#10;x=40520000;
#10;x=40530000;
#10;x=40540000;
#10;x=40550000;
#10;x=40560000;
#10;x=40570000;
#10;x=40580000;
#10;x=40590000;
#10;x=40600000;
#10;x=40610000;
#10;x=40620000;
#10;x=40630000;
#10;x=40640000;
#10;x=40650000;
#10;x=40660000;
#10;x=40670000;
#10;x=40680000;
#10;x=40690000;
#10;x=40700000;
#10;x=40710000;
#10;x=40720000;
#10;x=40730000;
#10;x=40740000;
#10;x=40750000;
#10;x=40760000;
#10;x=40770000;
#10;x=40780000;
#10;x=40790000;
#10;x=40800000;
#10;x=40810000;
#10;x=40820000;
#10;x=40830000;
#10;x=40840000;
#10;x=40850000;
#10;x=40860000;
#10;x=40870000;
#10;x=40880000;
#10;x=40890000;
#10;x=40900000;
#10;x=40910000;
#10;x=40920000;
#10;x=40930000;
#10;x=40940000;
#10;x=40950000;
#10;x=40960000;
#10;x=40970000;
#10;x=40980000;
#10;x=40990000;
#10;x=41000000;
#10;x=41010000;
#10;x=41020000;
#10;x=41030000;
#10;x=41040000;
#10;x=41050000;
#10;x=41060000;
#10;x=41070000;
#10;x=41080000;
#10;x=41090000;
#10;x=41100000;
#10;x=41110000;
#10;x=41120000;
#10;x=41130000;
#10;x=41140000;
#10;x=41150000;
#10;x=41160000;
#10;x=41170000;
#10;x=41180000;
#10;x=41190000;
#10;x=41200000;
#10;x=41210000;
#10;x=41220000;
#10;x=41230000;
#10;x=41240000;
#10;x=41250000;
#10;x=41260000;
#10;x=41270000;
#10;x=41280000;
#10;x=41290000;
#10;x=41300000;
#10;x=41310000;
#10;x=41320000;
#10;x=41330000;
#10;x=41340000;
#10;x=41350000;
#10;x=41360000;
#10;x=41370000;
#10;x=41380000;
#10;x=41390000;
#10;x=41400000;
#10;x=41410000;
#10;x=41420000;
#10;x=41430000;
#10;x=41440000;
#10;x=41450000;
#10;x=41460000;
#10;x=41470000;
#10;x=41480000;
#10;x=41490000;
#10;x=41500000;
#10;x=41510000;
#10;x=41520000;
#10;x=41530000;
#10;x=41540000;
#10;x=41550000;
#10;x=41560000;
#10;x=41570000;
#10;x=41580000;
#10;x=41590000;
#10;x=41600000;
#10;x=41610000;
#10;x=41620000;
#10;x=41630000;
#10;x=41640000;
#10;x=41650000;
#10;x=41660000;
#10;x=41670000;
#10;x=41680000;
#10;x=41690000;
#10;x=41700000;
#10;x=41710000;
#10;x=41720000;
#10;x=41730000;
#10;x=41740000;
#10;x=41750000;
#10;x=41760000;
#10;x=41770000;
#10;x=41780000;
#10;x=41790000;
#10;x=41800000;
#10;x=41810000;
#10;x=41820000;
#10;x=41830000;
#10;x=41840000;
#10;x=41850000;
#10;x=41860000;
#10;x=41870000;
#10;x=41880000;
#10;x=41890000;
#10;x=41900000;
#10;x=41910000;
#10;x=41920000;
#10;x=41930000;
#10;x=41940000;
#10;x=41950000;
#10;x=41960000;
#10;x=41970000;
#10;x=41980000;
#10;x=41990000;
#10;x=42000000;
#10;x=42010000;
#10;x=42020000;
#10;x=42030000;
#10;x=42040000;
#10;x=42050000;
#10;x=42060000;
#10;x=42070000;
#10;x=42080000;
#10;x=42090000;
#10;x=42100000;
#10;x=42110000;
#10;x=42120000;
#10;x=42130000;
#10;x=42140000;
#10;x=42150000;
#10;x=42160000;
#10;x=42170000;
#10;x=42180000;
#10;x=42190000;
#10;x=42200000;
#10;x=42210000;
#10;x=42220000;
#10;x=42230000;
#10;x=42240000;
#10;x=42250000;
#10;x=42260000;
#10;x=42270000;
#10;x=42280000;
#10;x=42290000;
#10;x=42300000;
#10;x=42310000;
#10;x=42320000;
#10;x=42330000;
#10;x=42340000;
#10;x=42350000;
#10;x=42360000;
#10;x=42370000;
#10;x=42380000;
#10;x=42390000;
#10;x=42400000;
#10;x=42410000;
#10;x=42420000;
#10;x=42430000;
#10;x=42440000;
#10;x=42450000;
#10;x=42460000;
#10;x=42470000;
#10;x=42480000;
#10;x=42490000;
#10;x=42500000;
#10;x=42510000;
#10;x=42520000;
#10;x=42530000;
#10;x=42540000;
#10;x=42550000;
#10;x=42560000;
#10;x=42570000;
#10;x=42580000;
#10;x=42590000;
#10;x=42600000;
#10;x=42610000;
#10;x=42620000;
#10;x=42630000;
#10;x=42640000;
#10;x=42650000;
#10;x=42660000;
#10;x=42670000;
#10;x=42680000;
#10;x=42690000;
#10;x=42700000;
#10;x=42710000;
#10;x=42720000;
#10;x=42730000;
#10;x=42740000;
#10;x=42750000;
#10;x=42760000;
#10;x=42770000;
#10;x=42780000;
#10;x=42790000;
#10;x=42800000;
#10;x=42810000;
#10;x=42820000;
#10;x=42830000;
#10;x=42840000;
#10;x=42850000;
#10;x=42860000;
#10;x=42870000;
#10;x=42880000;
#10;x=42890000;
#10;x=42900000;
#10;x=42910000;
#10;x=42920000;
#10;x=42930000;
#10;x=42940000;
#10;x=42950000;
#10;x=42960000;
#10;x=42970000;
#10;x=42980000;
#10;x=42990000;
#10;x=43000000;
#10;x=43010000;
#10;x=43020000;
#10;x=43030000;
#10;x=43040000;
#10;x=43050000;
#10;x=43060000;
#10;x=43070000;
#10;x=43080000;
#10;x=43090000;
#10;x=43100000;
#10;x=43110000;
#10;x=43120000;
#10;x=43130000;
#10;x=43140000;
#10;x=43150000;
#10;x=43160000;
#10;x=43170000;
#10;x=43180000;
#10;x=43190000;
#10;x=43200000;
#10;x=43210000;
#10;x=43220000;
#10;x=43230000;
#10;x=43240000;
#10;x=43250000;
#10;x=43260000;
#10;x=43270000;
#10;x=43280000;
#10;x=43290000;
#10;x=43300000;
#10;x=43310000;
#10;x=43320000;
#10;x=43330000;
#10;x=43340000;
#10;x=43350000;
#10;x=43360000;
#10;x=43370000;
#10;x=43380000;
#10;x=43390000;
#10;x=43400000;
#10;x=43410000;
#10;x=43420000;
#10;x=43430000;
#10;x=43440000;
#10;x=43450000;
#10;x=43460000;
#10;x=43470000;
#10;x=43480000;
#10;x=43490000;
#10;x=43500000;
#10;x=43510000;
#10;x=43520000;
#10;x=43530000;
#10;x=43540000;
#10;x=43550000;
#10;x=43560000;
#10;x=43570000;
#10;x=43580000;
#10;x=43590000;
#10;x=43600000;
#10;x=43610000;
#10;x=43620000;
#10;x=43630000;
#10;x=43640000;
#10;x=43650000;
#10;x=43660000;
#10;x=43670000;
#10;x=43680000;
#10;x=43690000;
#10;x=43700000;
#10;x=43710000;
#10;x=43720000;
#10;x=43730000;
#10;x=43740000;
#10;x=43750000;
#10;x=43760000;
#10;x=43770000;
#10;x=43780000;
#10;x=43790000;
#10;x=43800000;
#10;x=43810000;
#10;x=43820000;
#10;x=43830000;
#10;x=43840000;
#10;x=43850000;
#10;x=43860000;
#10;x=43870000;
#10;x=43880000;
#10;x=43890000;
#10;x=43900000;
#10;x=43910000;
#10;x=43920000;
#10;x=43930000;
#10;x=43940000;
#10;x=43950000;
#10;x=43960000;
#10;x=43970000;
#10;x=43980000;
#10;x=43990000;
#10;x=44000000;
#10;x=44010000;
#10;x=44020000;
#10;x=44030000;
#10;x=44040000;
#10;x=44050000;
#10;x=44060000;
#10;x=44070000;
#10;x=44080000;
#10;x=44090000;
#10;x=44100000;
#10;x=44110000;
#10;x=44120000;
#10;x=44130000;
#10;x=44140000;
#10;x=44150000;
#10;x=44160000;
#10;x=44170000;
#10;x=44180000;
#10;x=44190000;
#10;x=44200000;
#10;x=44210000;
#10;x=44220000;
#10;x=44230000;
#10;x=44240000;
#10;x=44250000;
#10;x=44260000;
#10;x=44270000;
#10;x=44280000;
#10;x=44290000;
#10;x=44300000;
#10;x=44310000;
#10;x=44320000;
#10;x=44330000;
#10;x=44340000;
#10;x=44350000;
#10;x=44360000;
#10;x=44370000;
#10;x=44380000;
#10;x=44390000;
#10;x=44400000;
#10;x=44410000;
#10;x=44420000;
#10;x=44430000;
#10;x=44440000;
#10;x=44450000;
#10;x=44460000;
#10;x=44470000;
#10;x=44480000;
#10;x=44490000;
#10;x=44500000;
#10;x=44510000;
#10;x=44520000;
#10;x=44530000;
#10;x=44540000;
#10;x=44550000;
#10;x=44560000;
#10;x=44570000;
#10;x=44580000;
#10;x=44590000;
#10;x=44600000;
#10;x=44610000;
#10;x=44620000;
#10;x=44630000;
#10;x=44640000;
#10;x=44650000;
#10;x=44660000;
#10;x=44670000;
#10;x=44680000;
#10;x=44690000;
#10;x=44700000;
#10;x=44710000;
#10;x=44720000;
#10;x=44730000;
#10;x=44740000;
#10;x=44750000;
#10;x=44760000;
#10;x=44770000;
#10;x=44780000;
#10;x=44790000;
#10;x=44800000;
#10;x=44810000;
#10;x=44820000;
#10;x=44830000;
#10;x=44840000;
#10;x=44850000;
#10;x=44860000;
#10;x=44870000;
#10;x=44880000;
#10;x=44890000;
#10;x=44900000;
#10;x=44910000;
#10;x=44920000;
#10;x=44930000;
#10;x=44940000;
#10;x=44950000;
#10;x=44960000;
#10;x=44970000;
#10;x=44980000;
#10;x=44990000;
#10;x=45000000;
#10;x=45010000;
#10;x=45020000;
#10;x=45030000;
#10;x=45040000;
#10;x=45050000;
#10;x=45060000;
#10;x=45070000;
#10;x=45080000;
#10;x=45090000;
#10;x=45100000;
#10;x=45110000;
#10;x=45120000;
#10;x=45130000;
#10;x=45140000;
#10;x=45150000;
#10;x=45160000;
#10;x=45170000;
#10;x=45180000;
#10;x=45190000;
#10;x=45200000;
#10;x=45210000;
#10;x=45220000;
#10;x=45230000;
#10;x=45240000;
#10;x=45250000;
#10;x=45260000;
#10;x=45270000;
#10;x=45280000;
#10;x=45290000;
#10;x=45300000;
#10;x=45310000;
#10;x=45320000;
#10;x=45330000;
#10;x=45340000;
#10;x=45350000;
#10;x=45360000;
#10;x=45370000;
#10;x=45380000;
#10;x=45390000;
#10;x=45400000;
#10;x=45410000;
#10;x=45420000;
#10;x=45430000;
#10;x=45440000;
#10;x=45450000;
#10;x=45460000;
#10;x=45470000;
#10;x=45480000;
#10;x=45490000;
#10;x=45500000;
#10;x=45510000;
#10;x=45520000;
#10;x=45530000;
#10;x=45540000;
#10;x=45550000;
#10;x=45560000;
#10;x=45570000;
#10;x=45580000;
#10;x=45590000;
#10;x=45600000;
#10;x=45610000;
#10;x=45620000;
#10;x=45630000;
#10;x=45640000;
#10;x=45650000;
#10;x=45660000;
#10;x=45670000;
#10;x=45680000;
#10;x=45690000;
#10;x=45700000;
#10;x=45710000;
#10;x=45720000;
#10;x=45730000;
#10;x=45740000;
#10;x=45750000;
#10;x=45760000;
#10;x=45770000;
#10;x=45780000;
#10;x=45790000;
#10;x=45800000;
#10;x=45810000;
#10;x=45820000;
#10;x=45830000;
#10;x=45840000;
#10;x=45850000;
#10;x=45860000;
#10;x=45870000;
#10;x=45880000;
#10;x=45890000;
#10;x=45900000;
#10;x=45910000;
#10;x=45920000;
#10;x=45930000;
#10;x=45940000;
#10;x=45950000;
#10;x=45960000;
#10;x=45970000;
#10;x=45980000;
#10;x=45990000;
#10;x=46000000;
#10;x=46010000;
#10;x=46020000;
#10;x=46030000;
#10;x=46040000;
#10;x=46050000;
#10;x=46060000;
#10;x=46070000;
#10;x=46080000;
#10;x=46090000;
#10;x=46100000;
#10;x=46110000;
#10;x=46120000;
#10;x=46130000;
#10;x=46140000;
#10;x=46150000;
#10;x=46160000;
#10;x=46170000;
#10;x=46180000;
#10;x=46190000;
#10;x=46200000;
#10;x=46210000;
#10;x=46220000;
#10;x=46230000;
#10;x=46240000;
#10;x=46250000;
#10;x=46260000;
#10;x=46270000;
#10;x=46280000;
#10;x=46290000;
#10;x=46300000;
#10;x=46310000;
#10;x=46320000;
#10;x=46330000;
#10;x=46340000;
#10;x=46350000;
#10;x=46360000;
#10;x=46370000;
#10;x=46380000;
#10;x=46390000;
#10;x=46400000;
#10;x=46410000;
#10;x=46420000;
#10;x=46430000;
#10;x=46440000;
#10;x=46450000;
#10;x=46460000;
#10;x=46470000;
#10;x=46480000;
#10;x=46490000;
#10;x=46500000;
#10;x=46510000;
#10;x=46520000;
#10;x=46530000;
#10;x=46540000;
#10;x=46550000;
#10;x=46560000;
#10;x=46570000;
#10;x=46580000;
#10;x=46590000;
#10;x=46600000;
#10;x=46610000;
#10;x=46620000;
#10;x=46630000;
#10;x=46640000;
#10;x=46650000;
#10;x=46660000;
#10;x=46670000;
#10;x=46680000;
#10;x=46690000;
#10;x=46700000;
#10;x=46710000;
#10;x=46720000;
#10;x=46730000;
#10;x=46740000;
#10;x=46750000;
#10;x=46760000;
#10;x=46770000;
#10;x=46780000;
#10;x=46790000;
#10;x=46800000;
#10;x=46810000;
#10;x=46820000;
#10;x=46830000;
#10;x=46840000;
#10;x=46850000;
#10;x=46860000;
#10;x=46870000;
#10;x=46880000;
#10;x=46890000;
#10;x=46900000;
#10;x=46910000;
#10;x=46920000;
#10;x=46930000;
#10;x=46940000;
#10;x=46950000;
#10;x=46960000;
#10;x=46970000;
#10;x=46980000;
#10;x=46990000;
#10;x=47000000;
#10;x=47010000;
#10;x=47020000;
#10;x=47030000;
#10;x=47040000;
#10;x=47050000;
#10;x=47060000;
#10;x=47070000;
#10;x=47080000;
#10;x=47090000;
#10;x=47100000;
#10;x=47110000;
#10;x=47120000;
#10;x=47130000;
#10;x=47140000;
#10;x=47150000;
#10;x=47160000;
#10;x=47170000;
#10;x=47180000;
#10;x=47190000;
#10;x=47200000;
#10;x=47210000;
#10;x=47220000;
#10;x=47230000;
#10;x=47240000;
#10;x=47250000;
#10;x=47260000;
#10;x=47270000;
#10;x=47280000;
#10;x=47290000;
#10;x=47300000;
#10;x=47310000;
#10;x=47320000;
#10;x=47330000;
#10;x=47340000;
#10;x=47350000;
#10;x=47360000;
#10;x=47370000;
#10;x=47380000;
#10;x=47390000;
#10;x=47400000;
#10;x=47410000;
#10;x=47420000;
#10;x=47430000;
#10;x=47440000;
#10;x=47450000;
#10;x=47460000;
#10;x=47470000;
#10;x=47480000;
#10;x=47490000;
#10;x=47500000;
#10;x=47510000;
#10;x=47520000;
#10;x=47530000;
#10;x=47540000;
#10;x=47550000;
#10;x=47560000;
#10;x=47570000;
#10;x=47580000;
#10;x=47590000;
#10;x=47600000;
#10;x=47610000;
#10;x=47620000;
#10;x=47630000;
#10;x=47640000;
#10;x=47650000;
#10;x=47660000;
#10;x=47670000;
#10;x=47680000;
#10;x=47690000;
#10;x=47700000;
#10;x=47710000;
#10;x=47720000;
#10;x=47730000;
#10;x=47740000;
#10;x=47750000;
#10;x=47760000;
#10;x=47770000;
#10;x=47780000;
#10;x=47790000;
#10;x=47800000;
#10;x=47810000;
#10;x=47820000;
#10;x=47830000;
#10;x=47840000;
#10;x=47850000;
#10;x=47860000;
#10;x=47870000;
#10;x=47880000;
#10;x=47890000;
#10;x=47900000;
#10;x=47910000;
#10;x=47920000;
#10;x=47930000;
#10;x=47940000;
#10;x=47950000;
#10;x=47960000;
#10;x=47970000;
#10;x=47980000;
#10;x=47990000;
#10;x=48000000;
#10;x=48010000;
#10;x=48020000;
#10;x=48030000;
#10;x=48040000;
#10;x=48050000;
#10;x=48060000;
#10;x=48070000;
#10;x=48080000;
#10;x=48090000;
#10;x=48100000;
#10;x=48110000;
#10;x=48120000;
#10;x=48130000;
#10;x=48140000;
#10;x=48150000;
#10;x=48160000;
#10;x=48170000;
#10;x=48180000;
#10;x=48190000;
#10;x=48200000;
#10;x=48210000;
#10;x=48220000;
#10;x=48230000;
#10;x=48240000;
#10;x=48250000;
#10;x=48260000;
#10;x=48270000;
#10;x=48280000;
#10;x=48290000;
#10;x=48300000;
#10;x=48310000;
#10;x=48320000;
#10;x=48330000;
#10;x=48340000;
#10;x=48350000;
#10;x=48360000;
#10;x=48370000;
#10;x=48380000;
#10;x=48390000;
#10;x=48400000;
#10;x=48410000;
#10;x=48420000;
#10;x=48430000;
#10;x=48440000;
#10;x=48450000;
#10;x=48460000;
#10;x=48470000;
#10;x=48480000;
#10;x=48490000;
#10;x=48500000;
#10;x=48510000;
#10;x=48520000;
#10;x=48530000;
#10;x=48540000;
#10;x=48550000;
#10;x=48560000;
#10;x=48570000;
#10;x=48580000;
#10;x=48590000;
#10;x=48600000;
#10;x=48610000;
#10;x=48620000;
#10;x=48630000;
#10;x=48640000;
#10;x=48650000;
#10;x=48660000;
#10;x=48670000;
#10;x=48680000;
#10;x=48690000;
#10;x=48700000;
#10;x=48710000;
#10;x=48720000;
#10;x=48730000;
#10;x=48740000;
#10;x=48750000;
#10;x=48760000;
#10;x=48770000;
#10;x=48780000;
#10;x=48790000;
#10;x=48800000;
#10;x=48810000;
#10;x=48820000;
#10;x=48830000;
#10;x=48840000;
#10;x=48850000;
#10;x=48860000;
#10;x=48870000;
#10;x=48880000;
#10;x=48890000;
#10;x=48900000;
#10;x=48910000;
#10;x=48920000;
#10;x=48930000;
#10;x=48940000;
#10;x=48950000;
#10;x=48960000;
#10;x=48970000;
#10;x=48980000;
#10;x=48990000;
#10;x=49000000;
#10;x=49010000;
#10;x=49020000;
#10;x=49030000;
#10;x=49040000;
#10;x=49050000;
#10;x=49060000;
#10;x=49070000;
#10;x=49080000;
#10;x=49090000;
#10;x=49100000;
#10;x=49110000;
#10;x=49120000;
#10;x=49130000;
#10;x=49140000;
#10;x=49150000;
#10;x=49160000;
#10;x=49170000;
#10;x=49180000;
#10;x=49190000;
#10;x=49200000;
#10;x=49210000;
#10;x=49220000;
#10;x=49230000;
#10;x=49240000;
#10;x=49250000;
#10;x=49260000;
#10;x=49270000;
#10;x=49280000;
#10;x=49290000;
#10;x=49300000;
#10;x=49310000;
#10;x=49320000;
#10;x=49330000;
#10;x=49340000;
#10;x=49350000;
#10;x=49360000;
#10;x=49370000;
#10;x=49380000;
#10;x=49390000;
#10;x=49400000;
#10;x=49410000;
#10;x=49420000;
#10;x=49430000;
#10;x=49440000;
#10;x=49450000;
#10;x=49460000;
#10;x=49470000;
#10;x=49480000;
#10;x=49490000;
#10;x=49500000;
#10;x=49510000;
#10;x=49520000;
#10;x=49530000;
#10;x=49540000;
#10;x=49550000;
#10;x=49560000;
#10;x=49570000;
#10;x=49580000;
#10;x=49590000;
#10;x=49600000;
#10;x=49610000;
#10;x=49620000;
#10;x=49630000;
#10;x=49640000;
#10;x=49650000;
#10;x=49660000;
#10;x=49670000;
#10;x=49680000;
#10;x=49690000;
#10;x=49700000;
#10;x=49710000;
#10;x=49720000;
#10;x=49730000;
#10;x=49740000;
#10;x=49750000;
#10;x=49760000;
#10;x=49770000;
#10;x=49780000;
#10;x=49790000;
#10;x=49800000;
#10;x=49810000;
#10;x=49820000;
#10;x=49830000;
#10;x=49840000;
#10;x=49850000;
#10;x=49860000;
#10;x=49870000;
#10;x=49880000;
#10;x=49890000;
#10;x=49900000;
#10;x=49910000;
#10;x=49920000;
#10;x=49930000;
#10;x=49940000;
#10;x=49950000;
#10;x=49960000;
#10;x=49970000;
#10;x=49980000;
#10;x=49990000;
#10;x=50000000;
#10;x=50010000;
#10;x=50020000;
#10;x=50030000;
#10;x=50040000;
#10;x=50050000;
#10;x=50060000;
#10;x=50070000;
#10;x=50080000;
#10;x=50090000;
#10;x=50100000;
#10;x=50110000;
#10;x=50120000;
#10;x=50130000;
#10;x=50140000;
#10;x=50150000;
#10;x=50160000;
#10;x=50170000;
#10;x=50180000;
#10;x=50190000;
#10;x=50200000;
#10;x=50210000;
#10;x=50220000;
#10;x=50230000;
#10;x=50240000;
#10;x=50250000;
#10;x=50260000;
#10;x=50270000;
#10;x=50280000;
#10;x=50290000;
#10;x=50300000;
#10;x=50310000;
#10;x=50320000;
#10;x=50330000;
#10;x=50340000;
#10;x=50350000;
#10;x=50360000;
#10;x=50370000;
#10;x=50380000;
#10;x=50390000;
#10;x=50400000;
#10;x=50410000;
#10;x=50420000;
#10;x=50430000;
#10;x=50440000;
#10;x=50450000;
#10;x=50460000;
#10;x=50470000;
#10;x=50480000;
#10;x=50490000;
#10;x=50500000;
#10;x=50510000;
#10;x=50520000;
#10;x=50530000;
#10;x=50540000;
#10;x=50550000;
#10;x=50560000;
#10;x=50570000;
#10;x=50580000;
#10;x=50590000;
#10;x=50600000;
#10;x=50610000;
#10;x=50620000;
#10;x=50630000;
#10;x=50640000;
#10;x=50650000;
#10;x=50660000;
#10;x=50670000;
#10;x=50680000;
#10;x=50690000;
#10;x=50700000;
#10;x=50710000;
#10;x=50720000;
#10;x=50730000;
#10;x=50740000;
#10;x=50750000;
#10;x=50760000;
#10;x=50770000;
#10;x=50780000;
#10;x=50790000;
#10;x=50800000;
#10;x=50810000;
#10;x=50820000;
#10;x=50830000;
#10;x=50840000;
#10;x=50850000;
#10;x=50860000;
#10;x=50870000;
#10;x=50880000;
#10;x=50890000;
#10;x=50900000;
#10;x=50910000;
#10;x=50920000;
#10;x=50930000;
#10;x=50940000;
#10;x=50950000;
#10;x=50960000;
#10;x=50970000;
#10;x=50980000;
#10;x=50990000;
#10;x=51000000;
#10;x=51010000;
#10;x=51020000;
#10;x=51030000;
#10;x=51040000;
#10;x=51050000;
#10;x=51060000;
#10;x=51070000;
#10;x=51080000;
#10;x=51090000;
#10;x=51100000;
#10;x=51110000;
#10;x=51120000;
#10;x=51130000;
#10;x=51140000;
#10;x=51150000;
#10;x=51160000;
#10;x=51170000;
#10;x=51180000;
#10;x=51190000;
#10;x=51200000;
#10;x=51210000;
#10;x=51220000;
#10;x=51230000;
#10;x=51240000;
#10;x=51250000;
#10;x=51260000;
#10;x=51270000;
#10;x=51280000;
#10;x=51290000;
#10;x=51300000;
#10;x=51310000;
#10;x=51320000;
#10;x=51330000;
#10;x=51340000;
#10;x=51350000;
#10;x=51360000;
#10;x=51370000;
#10;x=51380000;
#10;x=51390000;
#10;x=51400000;
#10;x=51410000;
#10;x=51420000;
#10;x=51430000;
#10;x=51440000;
#10;x=51450000;
#10;x=51460000;
#10;x=51470000;
#10;x=51480000;
#10;x=51490000;
#10;x=51500000;
#10;x=51510000;
#10;x=51520000;
#10;x=51530000;
#10;x=51540000;
#10;x=51550000;
#10;x=51560000;
#10;x=51570000;
#10;x=51580000;
#10;x=51590000;
#10;x=51600000;
#10;x=51610000;
#10;x=51620000;
#10;x=51630000;
#10;x=51640000;
#10;x=51650000;
#10;x=51660000;
#10;x=51670000;
#10;x=51680000;
#10;x=51690000;
#10;x=51700000;
#10;x=51710000;
#10;x=51720000;
#10;x=51730000;
#10;x=51740000;
#10;x=51750000;
#10;x=51760000;
#10;x=51770000;
#10;x=51780000;
#10;x=51790000;
#10;x=51800000;
#10;x=51810000;
#10;x=51820000;
#10;x=51830000;
#10;x=51840000;
#10;x=51850000;
#10;x=51860000;
#10;x=51870000;
#10;x=51880000;
#10;x=51890000;
#10;x=51900000;
#10;x=51910000;
#10;x=51920000;
#10;x=51930000;
#10;x=51940000;
#10;x=51950000;
#10;x=51960000;
#10;x=51970000;
#10;x=51980000;
#10;x=51990000;
#10;x=52000000;
#10;x=52010000;
#10;x=52020000;
#10;x=52030000;
#10;x=52040000;
#10;x=52050000;
#10;x=52060000;
#10;x=52070000;
#10;x=52080000;
#10;x=52090000;
#10;x=52100000;
#10;x=52110000;
#10;x=52120000;
#10;x=52130000;
#10;x=52140000;
#10;x=52150000;
#10;x=52160000;
#10;x=52170000;
#10;x=52180000;
#10;x=52190000;
#10;x=52200000;
#10;x=52210000;
#10;x=52220000;
#10;x=52230000;
#10;x=52240000;
#10;x=52250000;
#10;x=52260000;
#10;x=52270000;
#10;x=52280000;
#10;x=52290000;
#10;x=52300000;
#10;x=52310000;
#10;x=52320000;
#10;x=52330000;
#10;x=52340000;
#10;x=52350000;
#10;x=52360000;
#10;x=52370000;
#10;x=52380000;
#10;x=52390000;
#10;x=52400000;
#10;x=52410000;
#10;x=52420000;
#10;x=52430000;
#10;x=52440000;
#10;x=52450000;
#10;x=52460000;
#10;x=52470000;
#10;x=52480000;
#10;x=52490000;
#10;x=52500000;
#10;x=52510000;
#10;x=52520000;
#10;x=52530000;
#10;x=52540000;
#10;x=52550000;
#10;x=52560000;
#10;x=52570000;
#10;x=52580000;
#10;x=52590000;
#10;x=52600000;
#10;x=52610000;
#10;x=52620000;
#10;x=52630000;
#10;x=52640000;
#10;x=52650000;
#10;x=52660000;
#10;x=52670000;
#10;x=52680000;
#10;x=52690000;
#10;x=52700000;
#10;x=52710000;
#10;x=52720000;
#10;x=52730000;
#10;x=52740000;
#10;x=52750000;
#10;x=52760000;
#10;x=52770000;
#10;x=52780000;
#10;x=52790000;
#10;x=52800000;
#10;x=52810000;
#10;x=52820000;
#10;x=52830000;
#10;x=52840000;
#10;x=52850000;
#10;x=52860000;
#10;x=52870000;
#10;x=52880000;
#10;x=52890000;
#10;x=52900000;
#10;x=52910000;
#10;x=52920000;
#10;x=52930000;
#10;x=52940000;
#10;x=52950000;
#10;x=52960000;
#10;x=52970000;
#10;x=52980000;
#10;x=52990000;
#10;x=53000000;
#10;x=53010000;
#10;x=53020000;
#10;x=53030000;
#10;x=53040000;
#10;x=53050000;
#10;x=53060000;
#10;x=53070000;
#10;x=53080000;
#10;x=53090000;
#10;x=53100000;
#10;x=53110000;
#10;x=53120000;
#10;x=53130000;
#10;x=53140000;
#10;x=53150000;
#10;x=53160000;
#10;x=53170000;
#10;x=53180000;
#10;x=53190000;
#10;x=53200000;
#10;x=53210000;
#10;x=53220000;
#10;x=53230000;
#10;x=53240000;
#10;x=53250000;
#10;x=53260000;
#10;x=53270000;
#10;x=53280000;
#10;x=53290000;
#10;x=53300000;
#10;x=53310000;
#10;x=53320000;
#10;x=53330000;
#10;x=53340000;
#10;x=53350000;
#10;x=53360000;
#10;x=53370000;
#10;x=53380000;
#10;x=53390000;
#10;x=53400000;
#10;x=53410000;
#10;x=53420000;
#10;x=53430000;
#10;x=53440000;
#10;x=53450000;
#10;x=53460000;
#10;x=53470000;
#10;x=53480000;
#10;x=53490000;
#10;x=53500000;
#10;x=53510000;
#10;x=53520000;
#10;x=53530000;
#10;x=53540000;
#10;x=53550000;
#10;x=53560000;
#10;x=53570000;
#10;x=53580000;
#10;x=53590000;
#10;x=53600000;
#10;x=53610000;
#10;x=53620000;
#10;x=53630000;
#10;x=53640000;
#10;x=53650000;
#10;x=53660000;
#10;x=53670000;
#10;x=53680000;
#10;x=53690000;
#10;x=53700000;
#10;x=53710000;
#10;x=53720000;
#10;x=53730000;
#10;x=53740000;
#10;x=53750000;
#10;x=53760000;
#10;x=53770000;
#10;x=53780000;
#10;x=53790000;
#10;x=53800000;
#10;x=53810000;
#10;x=53820000;
#10;x=53830000;
#10;x=53840000;
#10;x=53850000;
#10;x=53860000;
#10;x=53870000;
#10;x=53880000;
#10;x=53890000;
#10;x=53900000;
#10;x=53910000;
#10;x=53920000;
#10;x=53930000;
#10;x=53940000;
#10;x=53950000;
#10;x=53960000;
#10;x=53970000;
#10;x=53980000;
#10;x=53990000;
#10;x=54000000;
#10;x=54010000;
#10;x=54020000;
#10;x=54030000;
#10;x=54040000;
#10;x=54050000;
#10;x=54060000;
#10;x=54070000;
#10;x=54080000;
#10;x=54090000;
#10;x=54100000;
#10;x=54110000;
#10;x=54120000;
#10;x=54130000;
#10;x=54140000;
#10;x=54150000;
#10;x=54160000;
#10;x=54170000;
#10;x=54180000;
#10;x=54190000;
#10;x=54200000;
#10;x=54210000;
#10;x=54220000;
#10;x=54230000;
#10;x=54240000;
#10;x=54250000;
#10;x=54260000;
#10;x=54270000;
#10;x=54280000;
#10;x=54290000;
#10;x=54300000;
#10;x=54310000;
#10;x=54320000;
#10;x=54330000;
#10;x=54340000;
#10;x=54350000;
#10;x=54360000;
#10;x=54370000;
#10;x=54380000;
#10;x=54390000;
#10;x=54400000;
#10;x=54410000;
#10;x=54420000;
#10;x=54430000;
#10;x=54440000;
#10;x=54450000;
#10;x=54460000;
#10;x=54470000;
#10;x=54480000;
#10;x=54490000;
#10;x=54500000;
#10;x=54510000;
#10;x=54520000;
#10;x=54530000;
#10;x=54540000;
#10;x=54550000;
#10;x=54560000;
#10;x=54570000;
#10;x=54580000;
#10;x=54590000;
#10;x=54600000;
#10;x=54610000;
#10;x=54620000;
#10;x=54630000;
#10;x=54640000;
#10;x=54650000;
#10;x=54660000;
#10;x=54670000;
#10;x=54680000;
#10;x=54690000;
#10;x=54700000;
#10;x=54710000;
#10;x=54720000;
#10;x=54730000;
#10;x=54740000;
#10;x=54750000;
#10;x=54760000;
#10;x=54770000;
#10;x=54780000;
#10;x=54790000;
#10;x=54800000;
#10;x=54810000;
#10;x=54820000;
#10;x=54830000;
#10;x=54840000;
#10;x=54850000;
#10;x=54860000;
#10;x=54870000;
#10;x=54880000;
#10;x=54890000;
#10;x=54900000;
#10;x=54910000;
#10;x=54920000;
#10;x=54930000;
#10;x=54940000;
#10;x=54950000;
#10;x=54960000;
#10;x=54970000;
#10;x=54980000;
#10;x=54990000;
#10;x=55000000;
#10;x=55010000;
#10;x=55020000;
#10;x=55030000;
#10;x=55040000;
#10;x=55050000;
#10;x=55060000;
#10;x=55070000;
#10;x=55080000;
#10;x=55090000;
#10;x=55100000;
#10;x=55110000;
#10;x=55120000;
#10;x=55130000;
#10;x=55140000;
#10;x=55150000;
#10;x=55160000;
#10;x=55170000;
#10;x=55180000;
#10;x=55190000;
#10;x=55200000;
#10;x=55210000;
#10;x=55220000;
#10;x=55230000;
#10;x=55240000;
#10;x=55250000;
#10;x=55260000;
#10;x=55270000;
#10;x=55280000;
#10;x=55290000;
#10;x=55300000;
#10;x=55310000;
#10;x=55320000;
#10;x=55330000;
#10;x=55340000;
#10;x=55350000;
#10;x=55360000;
#10;x=55370000;
#10;x=55380000;
#10;x=55390000;
#10;x=55400000;
#10;x=55410000;
#10;x=55420000;
#10;x=55430000;
#10;x=55440000;
#10;x=55450000;
#10;x=55460000;
#10;x=55470000;
#10;x=55480000;
#10;x=55490000;
#10;x=55500000;
#10;x=55510000;
#10;x=55520000;
#10;x=55530000;
#10;x=55540000;
#10;x=55550000;
#10;x=55560000;
#10;x=55570000;
#10;x=55580000;
#10;x=55590000;
#10;x=55600000;
#10;x=55610000;
#10;x=55620000;
#10;x=55630000;
#10;x=55640000;
#10;x=55650000;
#10;x=55660000;
#10;x=55670000;
#10;x=55680000;
#10;x=55690000;
#10;x=55700000;
#10;x=55710000;
#10;x=55720000;
#10;x=55730000;
#10;x=55740000;
#10;x=55750000;
#10;x=55760000;
#10;x=55770000;
#10;x=55780000;
#10;x=55790000;
#10;x=55800000;
#10;x=55810000;
#10;x=55820000;
#10;x=55830000;
#10;x=55840000;
#10;x=55850000;
#10;x=55860000;
#10;x=55870000;
#10;x=55880000;
#10;x=55890000;
#10;x=55900000;
#10;x=55910000;
#10;x=55920000;
#10;x=55930000;
#10;x=55940000;
#10;x=55950000;
#10;x=55960000;
#10;x=55970000;
#10;x=55980000;
#10;x=55990000;
#10;x=56000000;
#10;x=56010000;
#10;x=56020000;
#10;x=56030000;
#10;x=56040000;
#10;x=56050000;
#10;x=56060000;
#10;x=56070000;
#10;x=56080000;
#10;x=56090000;
#10;x=56100000;
#10;x=56110000;
#10;x=56120000;
#10;x=56130000;
#10;x=56140000;
#10;x=56150000;
#10;x=56160000;
#10;x=56170000;
#10;x=56180000;
#10;x=56190000;
#10;x=56200000;
#10;x=56210000;
#10;x=56220000;
#10;x=56230000;
#10;x=56240000;
#10;x=56250000;
#10;x=56260000;
#10;x=56270000;
#10;x=56280000;
#10;x=56290000;
#10;x=56300000;
#10;x=56310000;
#10;x=56320000;
#10;x=56330000;
#10;x=56340000;
#10;x=56350000;
#10;x=56360000;
#10;x=56370000;
#10;x=56380000;
#10;x=56390000;
#10;x=56400000;
#10;x=56410000;
#10;x=56420000;
#10;x=56430000;
#10;x=56440000;
#10;x=56450000;
#10;x=56460000;
#10;x=56470000;
#10;x=56480000;
#10;x=56490000;
#10;x=56500000;
#10;x=56510000;
#10;x=56520000;
#10;x=56530000;
#10;x=56540000;
#10;x=56550000;
#10;x=56560000;
#10;x=56570000;
#10;x=56580000;
#10;x=56590000;
#10;x=56600000;
#10;x=56610000;
#10;x=56620000;
#10;x=56630000;
#10;x=56640000;
#10;x=56650000;
#10;x=56660000;
#10;x=56670000;
#10;x=56680000;
#10;x=56690000;
#10;x=56700000;
#10;x=56710000;
#10;x=56720000;
#10;x=56730000;
#10;x=56740000;
#10;x=56750000;
#10;x=56760000;
#10;x=56770000;
#10;x=56780000;
#10;x=56790000;
#10;x=56800000;
#10;x=56810000;
#10;x=56820000;
#10;x=56830000;
#10;x=56840000;
#10;x=56850000;
#10;x=56860000;
#10;x=56870000;
#10;x=56880000;
#10;x=56890000;
#10;x=56900000;
#10;x=56910000;
#10;x=56920000;
#10;x=56930000;
#10;x=56940000;
#10;x=56950000;
#10;x=56960000;
#10;x=56970000;
#10;x=56980000;
#10;x=56990000;
#10;x=57000000;
#10;x=57010000;
#10;x=57020000;
#10;x=57030000;
#10;x=57040000;
#10;x=57050000;
#10;x=57060000;
#10;x=57070000;
#10;x=57080000;
#10;x=57090000;
#10;x=57100000;
#10;x=57110000;
#10;x=57120000;
#10;x=57130000;
#10;x=57140000;
#10;x=57150000;
#10;x=57160000;
#10;x=57170000;
#10;x=57180000;
#10;x=57190000;
#10;x=57200000;
#10;x=57210000;
#10;x=57220000;
#10;x=57230000;
#10;x=57240000;
#10;x=57250000;
#10;x=57260000;
#10;x=57270000;
#10;x=57280000;
#10;x=57290000;
#10;x=57300000;
#10;x=57310000;
#10;x=57320000;
#10;x=57330000;
#10;x=57340000;
#10;x=57350000;
#10;x=57360000;
#10;x=57370000;
#10;x=57380000;
#10;x=57390000;
#10;x=57400000;
#10;x=57410000;
#10;x=57420000;
#10;x=57430000;
#10;x=57440000;
#10;x=57450000;
#10;x=57460000;
#10;x=57470000;
#10;x=57480000;
#10;x=57490000;
#10;x=57500000;
#10;x=57510000;
#10;x=57520000;
#10;x=57530000;
#10;x=57540000;
#10;x=57550000;
#10;x=57560000;
#10;x=57570000;
#10;x=57580000;
#10;x=57590000;
#10;x=57600000;
#10;x=57610000;
#10;x=57620000;
#10;x=57630000;
#10;x=57640000;
#10;x=57650000;
#10;x=57660000;
#10;x=57670000;
#10;x=57680000;
#10;x=57690000;
#10;x=57700000;
#10;x=57710000;
#10;x=57720000;
#10;x=57730000;
#10;x=57740000;
#10;x=57750000;
#10;x=57760000;
#10;x=57770000;
#10;x=57780000;
#10;x=57790000;
#10;x=57800000;
#10;x=57810000;
#10;x=57820000;
#10;x=57830000;
#10;x=57840000;
#10;x=57850000;
#10;x=57860000;
#10;x=57870000;
#10;x=57880000;
#10;x=57890000;
#10;x=57900000;
#10;x=57910000;
#10;x=57920000;
#10;x=57930000;
#10;x=57940000;
#10;x=57950000;
#10;x=57960000;
#10;x=57970000;
#10;x=57980000;
#10;x=57990000;
#10;x=58000000;
#10;x=58010000;
#10;x=58020000;
#10;x=58030000;
#10;x=58040000;
#10;x=58050000;
#10;x=58060000;
#10;x=58070000;
#10;x=58080000;
#10;x=58090000;
#10;x=58100000;
#10;x=58110000;
#10;x=58120000;
#10;x=58130000;
#10;x=58140000;
#10;x=58150000;
#10;x=58160000;
#10;x=58170000;
#10;x=58180000;
#10;x=58190000;
#10;x=58200000;
#10;x=58210000;
#10;x=58220000;
#10;x=58230000;
#10;x=58240000;
#10;x=58250000;
#10;x=58260000;
#10;x=58270000;
#10;x=58280000;
#10;x=58290000;
#10;x=58300000;
#10;x=58310000;
#10;x=58320000;
#10;x=58330000;
#10;x=58340000;
#10;x=58350000;
#10;x=58360000;
#10;x=58370000;
#10;x=58380000;
#10;x=58390000;
#10;x=58400000;
#10;x=58410000;
#10;x=58420000;
#10;x=58430000;
#10;x=58440000;
#10;x=58450000;
#10;x=58460000;
#10;x=58470000;
#10;x=58480000;
#10;x=58490000;
#10;x=58500000;
#10;x=58510000;
#10;x=58520000;
#10;x=58530000;
#10;x=58540000;
#10;x=58550000;
#10;x=58560000;
#10;x=58570000;
#10;x=58580000;
#10;x=58590000;
#10;x=58600000;
#10;x=58610000;
#10;x=58620000;
#10;x=58630000;
#10;x=58640000;
#10;x=58650000;
#10;x=58660000;
#10;x=58670000;
#10;x=58680000;
#10;x=58690000;
#10;x=58700000;
#10;x=58710000;
#10;x=58720000;
#10;x=58730000;
#10;x=58740000;
#10;x=58750000;
#10;x=58760000;
#10;x=58770000;
#10;x=58780000;
#10;x=58790000;
#10;x=58800000;
#10;x=58810000;
#10;x=58820000;
#10;x=58830000;
#10;x=58840000;
#10;x=58850000;
#10;x=58860000;
#10;x=58870000;
#10;x=58880000;
#10;x=58890000;
#10;x=58900000;
#10;x=58910000;
#10;x=58920000;
#10;x=58930000;
#10;x=58940000;
#10;x=58950000;
#10;x=58960000;
#10;x=58970000;
#10;x=58980000;
#10;x=58990000;
#10;x=59000000;
#10;x=59010000;
#10;x=59020000;
#10;x=59030000;
#10;x=59040000;
#10;x=59050000;
#10;x=59060000;
#10;x=59070000;
#10;x=59080000;
#10;x=59090000;
#10;x=59100000;
#10;x=59110000;
#10;x=59120000;
#10;x=59130000;
#10;x=59140000;
#10;x=59150000;
#10;x=59160000;
#10;x=59170000;
#10;x=59180000;
#10;x=59190000;
#10;x=59200000;
#10;x=59210000;
#10;x=59220000;
#10;x=59230000;
#10;x=59240000;
#10;x=59250000;
#10;x=59260000;
#10;x=59270000;
#10;x=59280000;
#10;x=59290000;
#10;x=59300000;
#10;x=59310000;
#10;x=59320000;
#10;x=59330000;
#10;x=59340000;
#10;x=59350000;
#10;x=59360000;
#10;x=59370000;
#10;x=59380000;
#10;x=59390000;
#10;x=59400000;
#10;x=59410000;
#10;x=59420000;
#10;x=59430000;
#10;x=59440000;
#10;x=59450000;
#10;x=59460000;
#10;x=59470000;
#10;x=59480000;
#10;x=59490000;
#10;x=59500000;
#10;x=59510000;
#10;x=59520000;
#10;x=59530000;
#10;x=59540000;
#10;x=59550000;
#10;x=59560000;
#10;x=59570000;
#10;x=59580000;
#10;x=59590000;
#10;x=59600000;
#10;x=59610000;
#10;x=59620000;
#10;x=59630000;
#10;x=59640000;
#10;x=59650000;
#10;x=59660000;
#10;x=59670000;
#10;x=59680000;
#10;x=59690000;
#10;x=59700000;
#10;x=59710000;
#10;x=59720000;
#10;x=59730000;
#10;x=59740000;
#10;x=59750000;
#10;x=59760000;
#10;x=59770000;
#10;x=59780000;
#10;x=59790000;
#10;x=59800000;
#10;x=59810000;
#10;x=59820000;
#10;x=59830000;
#10;x=59840000;
#10;x=59850000;
#10;x=59860000;
#10;x=59870000;
#10;x=59880000;
#10;x=59890000;
#10;x=59900000;
#10;x=59910000;
#10;x=59920000;
#10;x=59930000;
#10;x=59940000;
#10;x=59950000;
#10;x=59960000;
#10;x=59970000;
#10;x=59980000;
#10;x=59990000;
#10;x=60000000;
#10;x=60010000;
#10;x=60020000;
#10;x=60030000;
#10;x=60040000;
#10;x=60050000;
#10;x=60060000;
#10;x=60070000;
#10;x=60080000;
#10;x=60090000;
#10;x=60100000;
#10;x=60110000;
#10;x=60120000;
#10;x=60130000;
#10;x=60140000;
#10;x=60150000;
#10;x=60160000;
#10;x=60170000;
#10;x=60180000;
#10;x=60190000;
#10;x=60200000;
#10;x=60210000;
#10;x=60220000;
#10;x=60230000;
#10;x=60240000;
#10;x=60250000;
#10;x=60260000;
#10;x=60270000;
#10;x=60280000;
#10;x=60290000;
#10;x=60300000;
#10;x=60310000;
#10;x=60320000;
#10;x=60330000;
#10;x=60340000;
#10;x=60350000;
#10;x=60360000;
#10;x=60370000;
#10;x=60380000;
#10;x=60390000;
#10;x=60400000;
#10;x=60410000;
#10;x=60420000;
#10;x=60430000;
#10;x=60440000;
#10;x=60450000;
#10;x=60460000;
#10;x=60470000;
#10;x=60480000;
#10;x=60490000;
#10;x=60500000;
#10;x=60510000;
#10;x=60520000;
#10;x=60530000;
#10;x=60540000;
#10;x=60550000;
#10;x=60560000;
#10;x=60570000;
#10;x=60580000;
#10;x=60590000;
#10;x=60600000;
#10;x=60610000;
#10;x=60620000;
#10;x=60630000;
#10;x=60640000;
#10;x=60650000;
#10;x=60660000;
#10;x=60670000;
#10;x=60680000;
#10;x=60690000;
#10;x=60700000;
#10;x=60710000;
#10;x=60720000;
#10;x=60730000;
#10;x=60740000;
#10;x=60750000;
#10;x=60760000;
#10;x=60770000;
#10;x=60780000;
#10;x=60790000;
#10;x=60800000;
#10;x=60810000;
#10;x=60820000;
#10;x=60830000;
#10;x=60840000;
#10;x=60850000;
#10;x=60860000;
#10;x=60870000;
#10;x=60880000;
#10;x=60890000;
#10;x=60900000;
#10;x=60910000;
#10;x=60920000;
#10;x=60930000;
#10;x=60940000;
#10;x=60950000;
#10;x=60960000;
#10;x=60970000;
#10;x=60980000;
#10;x=60990000;
#10;x=61000000;
#10;x=61010000;
#10;x=61020000;
#10;x=61030000;
#10;x=61040000;
#10;x=61050000;
#10;x=61060000;
#10;x=61070000;
#10;x=61080000;
#10;x=61090000;
#10;x=61100000;
#10;x=61110000;
#10;x=61120000;
#10;x=61130000;
#10;x=61140000;
#10;x=61150000;
#10;x=61160000;
#10;x=61170000;
#10;x=61180000;
#10;x=61190000;
#10;x=61200000;
#10;x=61210000;
#10;x=61220000;
#10;x=61230000;
#10;x=61240000;
#10;x=61250000;
#10;x=61260000;
#10;x=61270000;
#10;x=61280000;
#10;x=61290000;
#10;x=61300000;
#10;x=61310000;
#10;x=61320000;
#10;x=61330000;
#10;x=61340000;
#10;x=61350000;
#10;x=61360000;
#10;x=61370000;
#10;x=61380000;
#10;x=61390000;
#10;x=61400000;
#10;x=61410000;
#10;x=61420000;
#10;x=61430000;
#10;x=61440000;
#10;x=61450000;
#10;x=61460000;
#10;x=61470000;
#10;x=61480000;
#10;x=61490000;
#10;x=61500000;
#10;x=61510000;
#10;x=61520000;
#10;x=61530000;
#10;x=61540000;
#10;x=61550000;
#10;x=61560000;
#10;x=61570000;
#10;x=61580000;
#10;x=61590000;
#10;x=61600000;
#10;x=61610000;
#10;x=61620000;
#10;x=61630000;
#10;x=61640000;
#10;x=61650000;
#10;x=61660000;
#10;x=61670000;
#10;x=61680000;
#10;x=61690000;
#10;x=61700000;
#10;x=61710000;
#10;x=61720000;
#10;x=61730000;
#10;x=61740000;
#10;x=61750000;
#10;x=61760000;
#10;x=61770000;
#10;x=61780000;
#10;x=61790000;
#10;x=61800000;
#10;x=61810000;
#10;x=61820000;
#10;x=61830000;
#10;x=61840000;
#10;x=61850000;
#10;x=61860000;
#10;x=61870000;
#10;x=61880000;
#10;x=61890000;
#10;x=61900000;
#10;x=61910000;
#10;x=61920000;
#10;x=61930000;
#10;x=61940000;
#10;x=61950000;
#10;x=61960000;
#10;x=61970000;
#10;x=61980000;
#10;x=61990000;
#10;x=62000000;
#10;x=62010000;
#10;x=62020000;
#10;x=62030000;
#10;x=62040000;
#10;x=62050000;
#10;x=62060000;
#10;x=62070000;
#10;x=62080000;
#10;x=62090000;
#10;x=62100000;
#10;x=62110000;
#10;x=62120000;
#10;x=62130000;
#10;x=62140000;
#10;x=62150000;
#10;x=62160000;
#10;x=62170000;
#10;x=62180000;
#10;x=62190000;
#10;x=62200000;
#10;x=62210000;
#10;x=62220000;
#10;x=62230000;
#10;x=62240000;
#10;x=62250000;
#10;x=62260000;
#10;x=62270000;
#10;x=62280000;
#10;x=62290000;
#10;x=62300000;
#10;x=62310000;
#10;x=62320000;
#10;x=62330000;
#10;x=62340000;
#10;x=62350000;
#10;x=62360000;
#10;x=62370000;
#10;x=62380000;
#10;x=62390000;
#10;x=62400000;
#10;x=62410000;
#10;x=62420000;
#10;x=62430000;
#10;x=62440000;
#10;x=62450000;
#10;x=62460000;
#10;x=62470000;
#10;x=62480000;
#10;x=62490000;
#10;x=62500000;
#10;x=62510000;
#10;x=62520000;
#10;x=62530000;
#10;x=62540000;
#10;x=62550000;
#10;x=62560000;
#10;x=62570000;
#10;x=62580000;
#10;x=62590000;
#10;x=62600000;
#10;x=62610000;
#10;x=62620000;
#10;x=62630000;
#10;x=62640000;
#10;x=62650000;
#10;x=62660000;
#10;x=62670000;
#10;x=62680000;
#10;x=62690000;
#10;x=62700000;
#10;x=62710000;
#10;x=62720000;
#10;x=62730000;
#10;x=62740000;
#10;x=62750000;
#10;x=62760000;
#10;x=62770000;
#10;x=62780000;
#10;x=62790000;
#10;x=62800000;
#10;x=62810000;
#10;x=62820000;
#10;x=62830000;
#10;x=62840000;
#10;x=62850000;
#10;x=62860000;
#10;x=62870000;
#10;x=62880000;
#10;x=62890000;
#10;x=62900000;
#10;x=62910000;
#10;x=62920000;
#10;x=62930000;
#10;x=62940000;
#10;x=62950000;
#10;x=62960000;
#10;x=62970000;
#10;x=62980000;
#10;x=62990000;
#10;x=63000000;
#10;x=63010000;
#10;x=63020000;
#10;x=63030000;
#10;x=63040000;
#10;x=63050000;
#10;x=63060000;
#10;x=63070000;
#10;x=63080000;
#10;x=63090000;
#10;x=63100000;
#10;x=63110000;
#10;x=63120000;
#10;x=63130000;
#10;x=63140000;
#10;x=63150000;
#10;x=63160000;
#10;x=63170000;
#10;x=63180000;
#10;x=63190000;
#10;x=63200000;
#10;x=63210000;
#10;x=63220000;
#10;x=63230000;
#10;x=63240000;
#10;x=63250000;
#10;x=63260000;
#10;x=63270000;
#10;x=63280000;
#10;x=63290000;
#10;x=63300000;
#10;x=63310000;
#10;x=63320000;
#10;x=63330000;
#10;x=63340000;
#10;x=63350000;
#10;x=63360000;
#10;x=63370000;
#10;x=63380000;
#10;x=63390000;
#10;x=63400000;
#10;x=63410000;
#10;x=63420000;
#10;x=63430000;
#10;x=63440000;
#10;x=63450000;
#10;x=63460000;
#10;x=63470000;
#10;x=63480000;
#10;x=63490000;
#10;x=63500000;
#10;x=63510000;
#10;x=63520000;
#10;x=63530000;
#10;x=63540000;
#10;x=63550000;
#10;x=63560000;
#10;x=63570000;
#10;x=63580000;
#10;x=63590000;
#10;x=63600000;
#10;x=63610000;
#10;x=63620000;
#10;x=63630000;
#10;x=63640000;
#10;x=63650000;
#10;x=63660000;
#10;x=63670000;
#10;x=63680000;
#10;x=63690000;
#10;x=63700000;
#10;x=63710000;
#10;x=63720000;
#10;x=63730000;
#10;x=63740000;
#10;x=63750000;
#10;x=63760000;
#10;x=63770000;
#10;x=63780000;
#10;x=63790000;
#10;x=63800000;
#10;x=63810000;
#10;x=63820000;
#10;x=63830000;
#10;x=63840000;
#10;x=63850000;
#10;x=63860000;
#10;x=63870000;
#10;x=63880000;
#10;x=63890000;
#10;x=63900000;
#10;x=63910000;
#10;x=63920000;
#10;x=63930000;
#10;x=63940000;
#10;x=63950000;
#10;x=63960000;
#10;x=63970000;
#10;x=63980000;
#10;x=63990000;
#10;x=64000000;
#10;x=64010000;
#10;x=64020000;
#10;x=64030000;
#10;x=64040000;
#10;x=64050000;
#10;x=64060000;
#10;x=64070000;
#10;x=64080000;
#10;x=64090000;
#10;x=64100000;
#10;x=64110000;
#10;x=64120000;
#10;x=64130000;
#10;x=64140000;
#10;x=64150000;
#10;x=64160000;
#10;x=64170000;
#10;x=64180000;
#10;x=64190000;
#10;x=64200000;
#10;x=64210000;
#10;x=64220000;
#10;x=64230000;
#10;x=64240000;
#10;x=64250000;
#10;x=64260000;
#10;x=64270000;
#10;x=64280000;
#10;x=64290000;
#10;x=64300000;
#10;x=64310000;
#10;x=64320000;
#10;x=64330000;
#10;x=64340000;
#10;x=64350000;
#10;x=64360000;
#10;x=64370000;
#10;x=64380000;
#10;x=64390000;
#10;x=64400000;
#10;x=64410000;
#10;x=64420000;
#10;x=64430000;
#10;x=64440000;
#10;x=64450000;
#10;x=64460000;
#10;x=64470000;
#10;x=64480000;
#10;x=64490000;
#10;x=64500000;
#10;x=64510000;
#10;x=64520000;
#10;x=64530000;
#10;x=64540000;
#10;x=64550000;
#10;x=64560000;
#10;x=64570000;
#10;x=64580000;
#10;x=64590000;
#10;x=64600000;
#10;x=64610000;
#10;x=64620000;
#10;x=64630000;
#10;x=64640000;
#10;x=64650000;
#10;x=64660000;
#10;x=64670000;
#10;x=64680000;
#10;x=64690000;
#10;x=64700000;
#10;x=64710000;
#10;x=64720000;
#10;x=64730000;
#10;x=64740000;
#10;x=64750000;
#10;x=64760000;
#10;x=64770000;
#10;x=64780000;
#10;x=64790000;
#10;x=64800000;
#10;x=64810000;
#10;x=64820000;
#10;x=64830000;
#10;x=64840000;
#10;x=64850000;
#10;x=64860000;
#10;x=64870000;
#10;x=64880000;
#10;x=64890000;
#10;x=64900000;
#10;x=64910000;
#10;x=64920000;
#10;x=64930000;
#10;x=64940000;
#10;x=64950000;
#10;x=64960000;
#10;x=64970000;
#10;x=64980000;
#10;x=64990000;
#10;x=65000000;
#10;x=65010000;
#10;x=65020000;
#10;x=65030000;
#10;x=65040000;
#10;x=65050000;
#10;x=65060000;
#10;x=65070000;
#10;x=65080000;
#10;x=65090000;
#10;x=65100000;
#10;x=65110000;
#10;x=65120000;
#10;x=65130000;
#10;x=65140000;
#10;x=65150000;
#10;x=65160000;
#10;x=65170000;
#10;x=65180000;
#10;x=65190000;
#10;x=65200000;
#10;x=65210000;
#10;x=65220000;
#10;x=65230000;
#10;x=65240000;
#10;x=65250000;
#10;x=65260000;
#10;x=65270000;
#10;x=65280000;
#10;x=65290000;
#10;x=65300000;
#10;x=65310000;
#10;x=65320000;
#10;x=65330000;
#10;x=65340000;
#10;x=65350000;
#10;x=65360000;
#10;x=65370000;
#10;x=65380000;
#10;x=65390000;
#10;x=65400000;
#10;x=65410000;
#10;x=65420000;
#10;x=65430000;
#10;x=65440000;
#10;x=65450000;
#10;x=65460000;
#10;x=65470000;
#10;x=65480000;
#10;x=65490000;
#10;x=65500000;
#10;x=65510000;
#10;x=65520000;
#10;x=65530000;
#10;x=65540000;
#10;x=65550000;
#10;x=65560000;
#10;x=65570000;
#10;x=65580000;
#10;x=65590000;
#10;x=65600000;
#10;x=65610000;
#10;x=65620000;
#10;x=65630000;
#10;x=65640000;
#10;x=65650000;
#10;x=65660000;
#10;x=65670000;
#10;x=65680000;
#10;x=65690000;
#10;x=65700000;
#10;x=65710000;
#10;x=65720000;
#10;x=65730000;
#10;x=65740000;
#10;x=65750000;
#10;x=65760000;
#10;x=65770000;
#10;x=65780000;
#10;x=65790000;
#10;x=65800000;
#10;x=65810000;
#10;x=65820000;
#10;x=65830000;
#10;x=65840000;
#10;x=65850000;
#10;x=65860000;
#10;x=65870000;
#10;x=65880000;
#10;x=65890000;
#10;x=65900000;
#10;x=65910000;
#10;x=65920000;
#10;x=65930000;
#10;x=65940000;
#10;x=65950000;
#10;x=65960000;
#10;x=65970000;
#10;x=65980000;
#10;x=65990000;
#10;x=66000000;
#10;x=66010000;
#10;x=66020000;
#10;x=66030000;
#10;x=66040000;
#10;x=66050000;
#10;x=66060000;
#10;x=66070000;
#10;x=66080000;
#10;x=66090000;
#10;x=66100000;
#10;x=66110000;
#10;x=66120000;
#10;x=66130000;
#10;x=66140000;
#10;x=66150000;
#10;x=66160000;
#10;x=66170000;
#10;x=66180000;
#10;x=66190000;
#10;x=66200000;
#10;x=66210000;
#10;x=66220000;
#10;x=66230000;
#10;x=66240000;
#10;x=66250000;
#10;x=66260000;
#10;x=66270000;
#10;x=66280000;
#10;x=66290000;
#10;x=66300000;
#10;x=66310000;
#10;x=66320000;
#10;x=66330000;
#10;x=66340000;
#10;x=66350000;
#10;x=66360000;
#10;x=66370000;
#10;x=66380000;
#10;x=66390000;
#10;x=66400000;
#10;x=66410000;
#10;x=66420000;
#10;x=66430000;
#10;x=66440000;
#10;x=66450000;
#10;x=66460000;
#10;x=66470000;
#10;x=66480000;
#10;x=66490000;
#10;x=66500000;
#10;x=66510000;
#10;x=66520000;
#10;x=66530000;
#10;x=66540000;
#10;x=66550000;
#10;x=66560000;
#10;x=66570000;
#10;x=66580000;
#10;x=66590000;
#10;x=66600000;
#10;x=66610000;
#10;x=66620000;
#10;x=66630000;
#10;x=66640000;
#10;x=66650000;
#10;x=66660000;
#10;x=66670000;
#10;x=66680000;
#10;x=66690000;
#10;x=66700000;
#10;x=66710000;
#10;x=66720000;
#10;x=66730000;
#10;x=66740000;
#10;x=66750000;
#10;x=66760000;
#10;x=66770000;
#10;x=66780000;
#10;x=66790000;
#10;x=66800000;
#10;x=66810000;
#10;x=66820000;
#10;x=66830000;
#10;x=66840000;
#10;x=66850000;
#10;x=66860000;
#10;x=66870000;
#10;x=66880000;
#10;x=66890000;
#10;x=66900000;
#10;x=66910000;
#10;x=66920000;
#10;x=66930000;
#10;x=66940000;
#10;x=66950000;
#10;x=66960000;
#10;x=66970000;
#10;x=66980000;
#10;x=66990000;
#10;x=67000000;
#10;x=67010000;
#10;x=67020000;
#10;x=67030000;
#10;x=67040000;
#10;x=67050000;
#10;x=67060000;
#10;x=67070000;
#10;x=67080000;
#10;x=67090000;
#10;x=67100000;
#10;x=67110000;
#10;x=67120000;
#10;x=67130000;
#10;x=67140000;
#10;x=67150000;
#10;x=67160000;
#10;x=67170000;
#10;x=67180000;
#10;x=67190000;
#10;x=67200000;
#10;x=67210000;
#10;x=67220000;
#10;x=67230000;
#10;x=67240000;
#10;x=67250000;
#10;x=67260000;
#10;x=67270000;
#10;x=67280000;
#10;x=67290000;
#10;x=67300000;
#10;x=67310000;
#10;x=67320000;
#10;x=67330000;
#10;x=67340000;
#10;x=67350000;
#10;x=67360000;
#10;x=67370000;
#10;x=67380000;
#10;x=67390000;
#10;x=67400000;
#10;x=67410000;
#10;x=67420000;
#10;x=67430000;
#10;x=67440000;
#10;x=67450000;
#10;x=67460000;
#10;x=67470000;
#10;x=67480000;
#10;x=67490000;
#10;x=67500000;
#10;x=67510000;
#10;x=67520000;
#10;x=67530000;
#10;x=67540000;
#10;x=67550000;
#10;x=67560000;
#10;x=67570000;
#10;x=67580000;
#10;x=67590000;
#10;x=67600000;
#10;x=67610000;
#10;x=67620000;
#10;x=67630000;
#10;x=67640000;
#10;x=67650000;
#10;x=67660000;
#10;x=67670000;
#10;x=67680000;
#10;x=67690000;
#10;x=67700000;
#10;x=67710000;
#10;x=67720000;
#10;x=67730000;
#10;x=67740000;
#10;x=67750000;
#10;x=67760000;
#10;x=67770000;
#10;x=67780000;
#10;x=67790000;
#10;x=67800000;
#10;x=67810000;
#10;x=67820000;
#10;x=67830000;
#10;x=67840000;
#10;x=67850000;
#10;x=67860000;
#10;x=67870000;
#10;x=67880000;
#10;x=67890000;
#10;x=67900000;
#10;x=67910000;
#10;x=67920000;
#10;x=67930000;
#10;x=67940000;
#10;x=67950000;
#10;x=67960000;
#10;x=67970000;
#10;x=67980000;
#10;x=67990000;
#10;x=68000000;
#10;x=68010000;
#10;x=68020000;
#10;x=68030000;
#10;x=68040000;
#10;x=68050000;
#10;x=68060000;
#10;x=68070000;
#10;x=68080000;
#10;x=68090000;
#10;x=68100000;
#10;x=68110000;
#10;x=68120000;
#10;x=68130000;
#10;x=68140000;
#10;x=68150000;
#10;x=68160000;
#10;x=68170000;
#10;x=68180000;
#10;x=68190000;
#10;x=68200000;
#10;x=68210000;
#10;x=68220000;
#10;x=68230000;
#10;x=68240000;
#10;x=68250000;
#10;x=68260000;
#10;x=68270000;
#10;x=68280000;
#10;x=68290000;
#10;x=68300000;
#10;x=68310000;
#10;x=68320000;
#10;x=68330000;
#10;x=68340000;
#10;x=68350000;
#10;x=68360000;
#10;x=68370000;
#10;x=68380000;
#10;x=68390000;
#10;x=68400000;
#10;x=68410000;
#10;x=68420000;
#10;x=68430000;
#10;x=68440000;
#10;x=68450000;
#10;x=68460000;
#10;x=68470000;
#10;x=68480000;
#10;x=68490000;
#10;x=68500000;
#10;x=68510000;
#10;x=68520000;
#10;x=68530000;
#10;x=68540000;
#10;x=68550000;
#10;x=68560000;
#10;x=68570000;
#10;x=68580000;
#10;x=68590000;
#10;x=68600000;
#10;x=68610000;
#10;x=68620000;
#10;x=68630000;
#10;x=68640000;
#10;x=68650000;
#10;x=68660000;
#10;x=68670000;
#10;x=68680000;
#10;x=68690000;
#10;x=68700000;
#10;x=68710000;
#10;x=68720000;
#10;x=68730000;
#10;x=68740000;
#10;x=68750000;
#10;x=68760000;
#10;x=68770000;
#10;x=68780000;
#10;x=68790000;
#10;x=68800000;
#10;x=68810000;
#10;x=68820000;
#10;x=68830000;
#10;x=68840000;
#10;x=68850000;
#10;x=68860000;
#10;x=68870000;
#10;x=68880000;
#10;x=68890000;
#10;x=68900000;
#10;x=68910000;
#10;x=68920000;
#10;x=68930000;
#10;x=68940000;
#10;x=68950000;
#10;x=68960000;
#10;x=68970000;
#10;x=68980000;
#10;x=68990000;
#10;x=69000000;
#10;x=69010000;
#10;x=69020000;
#10;x=69030000;
#10;x=69040000;
#10;x=69050000;
#10;x=69060000;
#10;x=69070000;
#10;x=69080000;
#10;x=69090000;
#10;x=69100000;
#10;x=69110000;
#10;x=69120000;
#10;x=69130000;
#10;x=69140000;
#10;x=69150000;
#10;x=69160000;
#10;x=69170000;
#10;x=69180000;
#10;x=69190000;
#10;x=69200000;
#10;x=69210000;
#10;x=69220000;
#10;x=69230000;
#10;x=69240000;
#10;x=69250000;
#10;x=69260000;
#10;x=69270000;
#10;x=69280000;
#10;x=69290000;
#10;x=69300000;
#10;x=69310000;
#10;x=69320000;
#10;x=69330000;
#10;x=69340000;
#10;x=69350000;
#10;x=69360000;
#10;x=69370000;
#10;x=69380000;
#10;x=69390000;
#10;x=69400000;
#10;x=69410000;
#10;x=69420000;
#10;x=69430000;
#10;x=69440000;
#10;x=69450000;
#10;x=69460000;
#10;x=69470000;
#10;x=69480000;
#10;x=69490000;
#10;x=69500000;
#10;x=69510000;
#10;x=69520000;
#10;x=69530000;
#10;x=69540000;
#10;x=69550000;
#10;x=69560000;
#10;x=69570000;
#10;x=69580000;
#10;x=69590000;
#10;x=69600000;
#10;x=69610000;
#10;x=69620000;
#10;x=69630000;
#10;x=69640000;
#10;x=69650000;
#10;x=69660000;
#10;x=69670000;
#10;x=69680000;
#10;x=69690000;
#10;x=69700000;
#10;x=69710000;
#10;x=69720000;
#10;x=69730000;
#10;x=69740000;
#10;x=69750000;
#10;x=69760000;
#10;x=69770000;
#10;x=69780000;
#10;x=69790000;
#10;x=69800000;
#10;x=69810000;
#10;x=69820000;
#10;x=69830000;
#10;x=69840000;
#10;x=69850000;
#10;x=69860000;
#10;x=69870000;
#10;x=69880000;
#10;x=69890000;
#10;x=69900000;
#10;x=69910000;
#10;x=69920000;
#10;x=69930000;
#10;x=69940000;
#10;x=69950000;
#10;x=69960000;
#10;x=69970000;
#10;x=69980000;
#10;x=69990000;
#10;x=70000000;
#10;x=70010000;
#10;x=70020000;
#10;x=70030000;
#10;x=70040000;
#10;x=70050000;
#10;x=70060000;
#10;x=70070000;
#10;x=70080000;
#10;x=70090000;
#10;x=70100000;
#10;x=70110000;
#10;x=70120000;
#10;x=70130000;
#10;x=70140000;
#10;x=70150000;
#10;x=70160000;
#10;x=70170000;
#10;x=70180000;
#10;x=70190000;
#10;x=70200000;
#10;x=70210000;
#10;x=70220000;
#10;x=70230000;
#10;x=70240000;
#10;x=70250000;
#10;x=70260000;
#10;x=70270000;
#10;x=70280000;
#10;x=70290000;
#10;x=70300000;
#10;x=70310000;
#10;x=70320000;
#10;x=70330000;
#10;x=70340000;
#10;x=70350000;
#10;x=70360000;
#10;x=70370000;
#10;x=70380000;
#10;x=70390000;
#10;x=70400000;
#10;x=70410000;
#10;x=70420000;
#10;x=70430000;
#10;x=70440000;
#10;x=70450000;
#10;x=70460000;
#10;x=70470000;
#10;x=70480000;
#10;x=70490000;
#10;x=70500000;
#10;x=70510000;
#10;x=70520000;
#10;x=70530000;
#10;x=70540000;
#10;x=70550000;
#10;x=70560000;
#10;x=70570000;
#10;x=70580000;
#10;x=70590000;
#10;x=70600000;
#10;x=70610000;
#10;x=70620000;
#10;x=70630000;
#10;x=70640000;
#10;x=70650000;
#10;x=70660000;
#10;x=70670000;
#10;x=70680000;
#10;x=70690000;
#10;x=70700000;
#10;x=70710000;
#10;x=70720000;
#10;x=70730000;
#10;x=70740000;
#10;x=70750000;
#10;x=70760000;
#10;x=70770000;
#10;x=70780000;
#10;x=70790000;
#10;x=70800000;
#10;x=70810000;
#10;x=70820000;
#10;x=70830000;
#10;x=70840000;
#10;x=70850000;
#10;x=70860000;
#10;x=70870000;
#10;x=70880000;
#10;x=70890000;
#10;x=70900000;
#10;x=70910000;
#10;x=70920000;
#10;x=70930000;
#10;x=70940000;
#10;x=70950000;
#10;x=70960000;
#10;x=70970000;
#10;x=70980000;
#10;x=70990000;
#10;x=71000000;
#10;x=71010000;
#10;x=71020000;
#10;x=71030000;
#10;x=71040000;
#10;x=71050000;
#10;x=71060000;
#10;x=71070000;
#10;x=71080000;
#10;x=71090000;
#10;x=71100000;
#10;x=71110000;
#10;x=71120000;
#10;x=71130000;
#10;x=71140000;
#10;x=71150000;
#10;x=71160000;
#10;x=71170000;
#10;x=71180000;
#10;x=71190000;
#10;x=71200000;
#10;x=71210000;
#10;x=71220000;
#10;x=71230000;
#10;x=71240000;
#10;x=71250000;
#10;x=71260000;
#10;x=71270000;
#10;x=71280000;
#10;x=71290000;
#10;x=71300000;
#10;x=71310000;
#10;x=71320000;
#10;x=71330000;
#10;x=71340000;
#10;x=71350000;
#10;x=71360000;
#10;x=71370000;
#10;x=71380000;
#10;x=71390000;
#10;x=71400000;
#10;x=71410000;
#10;x=71420000;
#10;x=71430000;
#10;x=71440000;
#10;x=71450000;
#10;x=71460000;
#10;x=71470000;
#10;x=71480000;
#10;x=71490000;
#10;x=71500000;
#10;x=71510000;
#10;x=71520000;
#10;x=71530000;
#10;x=71540000;
#10;x=71550000;
#10;x=71560000;
#10;x=71570000;
#10;x=71580000;
#10;x=71590000;
#10;x=71600000;
#10;x=71610000;
#10;x=71620000;
#10;x=71630000;
#10;x=71640000;
#10;x=71650000;
#10;x=71660000;
#10;x=71670000;
#10;x=71680000;
#10;x=71690000;
#10;x=71700000;
#10;x=71710000;
#10;x=71720000;
#10;x=71730000;
#10;x=71740000;
#10;x=71750000;
#10;x=71760000;
#10;x=71770000;
#10;x=71780000;
#10;x=71790000;
#10;x=71800000;
#10;x=71810000;
#10;x=71820000;
#10;x=71830000;
#10;x=71840000;
#10;x=71850000;
#10;x=71860000;
#10;x=71870000;
#10;x=71880000;
#10;x=71890000;
#10;x=71900000;
#10;x=71910000;
#10;x=71920000;
#10;x=71930000;
#10;x=71940000;
#10;x=71950000;
#10;x=71960000;
#10;x=71970000;
#10;x=71980000;
#10;x=71990000;
#10;x=72000000;
#10;x=72010000;
#10;x=72020000;
#10;x=72030000;
#10;x=72040000;
#10;x=72050000;
#10;x=72060000;
#10;x=72070000;
#10;x=72080000;
#10;x=72090000;
#10;x=72100000;
#10;x=72110000;
#10;x=72120000;
#10;x=72130000;
#10;x=72140000;
#10;x=72150000;
#10;x=72160000;
#10;x=72170000;
#10;x=72180000;
#10;x=72190000;
#10;x=72200000;
#10;x=72210000;
#10;x=72220000;
#10;x=72230000;
#10;x=72240000;
#10;x=72250000;
#10;x=72260000;
#10;x=72270000;
#10;x=72280000;
#10;x=72290000;
#10;x=72300000;
#10;x=72310000;
#10;x=72320000;
#10;x=72330000;
#10;x=72340000;
#10;x=72350000;
#10;x=72360000;
#10;x=72370000;
#10;x=72380000;
#10;x=72390000;
#10;x=72400000;
#10;x=72410000;
#10;x=72420000;
#10;x=72430000;
#10;x=72440000;
#10;x=72450000;
#10;x=72460000;
#10;x=72470000;
#10;x=72480000;
#10;x=72490000;
#10;x=72500000;
#10;x=72510000;
#10;x=72520000;
#10;x=72530000;
#10;x=72540000;
#10;x=72550000;
#10;x=72560000;
#10;x=72570000;
#10;x=72580000;
#10;x=72590000;
#10;x=72600000;
#10;x=72610000;
#10;x=72620000;
#10;x=72630000;
#10;x=72640000;
#10;x=72650000;
#10;x=72660000;
#10;x=72670000;
#10;x=72680000;
#10;x=72690000;
#10;x=72700000;
#10;x=72710000;
#10;x=72720000;
#10;x=72730000;
#10;x=72740000;
#10;x=72750000;
#10;x=72760000;
#10;x=72770000;
#10;x=72780000;
#10;x=72790000;
#10;x=72800000;
#10;x=72810000;
#10;x=72820000;
#10;x=72830000;
#10;x=72840000;
#10;x=72850000;
#10;x=72860000;
#10;x=72870000;
#10;x=72880000;
#10;x=72890000;
#10;x=72900000;
#10;x=72910000;
#10;x=72920000;
#10;x=72930000;
#10;x=72940000;
#10;x=72950000;
#10;x=72960000;
#10;x=72970000;
#10;x=72980000;
#10;x=72990000;
#10;x=73000000;
#10;x=73010000;
#10;x=73020000;
#10;x=73030000;
#10;x=73040000;
#10;x=73050000;
#10;x=73060000;
#10;x=73070000;
#10;x=73080000;
#10;x=73090000;
#10;x=73100000;
#10;x=73110000;
#10;x=73120000;
#10;x=73130000;
#10;x=73140000;
#10;x=73150000;
#10;x=73160000;
#10;x=73170000;
#10;x=73180000;
#10;x=73190000;
#10;x=73200000;
#10;x=73210000;
#10;x=73220000;
#10;x=73230000;
#10;x=73240000;
#10;x=73250000;
#10;x=73260000;
#10;x=73270000;
#10;x=73280000;
#10;x=73290000;
#10;x=73300000;
#10;x=73310000;
#10;x=73320000;
#10;x=73330000;
#10;x=73340000;
#10;x=73350000;
#10;x=73360000;
#10;x=73370000;
#10;x=73380000;
#10;x=73390000;
#10;x=73400000;
#10;x=73410000;
#10;x=73420000;
#10;x=73430000;
#10;x=73440000;
#10;x=73450000;
#10;x=73460000;
#10;x=73470000;
#10;x=73480000;
#10;x=73490000;
#10;x=73500000;
#10;x=73510000;
#10;x=73520000;
#10;x=73530000;
#10;x=73540000;
#10;x=73550000;
#10;x=73560000;
#10;x=73570000;
#10;x=73580000;
#10;x=73590000;
#10;x=73600000;
#10;x=73610000;
#10;x=73620000;
#10;x=73630000;
#10;x=73640000;
#10;x=73650000;
#10;x=73660000;
#10;x=73670000;
#10;x=73680000;
#10;x=73690000;
#10;x=73700000;
#10;x=73710000;
#10;x=73720000;
#10;x=73730000;
#10;x=73740000;
#10;x=73750000;
#10;x=73760000;
#10;x=73770000;
#10;x=73780000;
#10;x=73790000;
#10;x=73800000;
#10;x=73810000;
#10;x=73820000;
#10;x=73830000;
#10;x=73840000;
#10;x=73850000;
#10;x=73860000;
#10;x=73870000;
#10;x=73880000;
#10;x=73890000;
#10;x=73900000;
#10;x=73910000;
#10;x=73920000;
#10;x=73930000;
#10;x=73940000;
#10;x=73950000;
#10;x=73960000;
#10;x=73970000;
#10;x=73980000;
#10;x=73990000;
#10;x=74000000;
#10;x=74010000;
#10;x=74020000;
#10;x=74030000;
#10;x=74040000;
#10;x=74050000;
#10;x=74060000;
#10;x=74070000;
#10;x=74080000;
#10;x=74090000;
#10;x=74100000;
#10;x=74110000;
#10;x=74120000;
#10;x=74130000;
#10;x=74140000;
#10;x=74150000;
#10;x=74160000;
#10;x=74170000;
#10;x=74180000;
#10;x=74190000;
#10;x=74200000;
#10;x=74210000;
#10;x=74220000;
#10;x=74230000;
#10;x=74240000;
#10;x=74250000;
#10;x=74260000;
#10;x=74270000;
#10;x=74280000;
#10;x=74290000;
#10;x=74300000;
#10;x=74310000;
#10;x=74320000;
#10;x=74330000;
#10;x=74340000;
#10;x=74350000;
#10;x=74360000;
#10;x=74370000;
#10;x=74380000;
#10;x=74390000;
#10;x=74400000;
#10;x=74410000;
#10;x=74420000;
#10;x=74430000;
#10;x=74440000;
#10;x=74450000;
#10;x=74460000;
#10;x=74470000;
#10;x=74480000;
#10;x=74490000;
#10;x=74500000;
#10;x=74510000;
#10;x=74520000;
#10;x=74530000;
#10;x=74540000;
#10;x=74550000;
#10;x=74560000;
#10;x=74570000;
#10;x=74580000;
#10;x=74590000;
#10;x=74600000;
#10;x=74610000;
#10;x=74620000;
#10;x=74630000;
#10;x=74640000;
#10;x=74650000;
#10;x=74660000;
#10;x=74670000;
#10;x=74680000;
#10;x=74690000;
#10;x=74700000;
#10;x=74710000;
#10;x=74720000;
#10;x=74730000;
#10;x=74740000;
#10;x=74750000;
#10;x=74760000;
#10;x=74770000;
#10;x=74780000;
#10;x=74790000;
#10;x=74800000;
#10;x=74810000;
#10;x=74820000;
#10;x=74830000;
#10;x=74840000;
#10;x=74850000;
#10;x=74860000;
#10;x=74870000;
#10;x=74880000;
#10;x=74890000;
#10;x=74900000;
#10;x=74910000;
#10;x=74920000;
#10;x=74930000;
#10;x=74940000;
#10;x=74950000;
#10;x=74960000;
#10;x=74970000;
#10;x=74980000;
#10;x=74990000;
#10;x=75000000;
#10;x=75010000;
#10;x=75020000;
#10;x=75030000;
#10;x=75040000;
#10;x=75050000;
#10;x=75060000;
#10;x=75070000;
#10;x=75080000;
#10;x=75090000;
#10;x=75100000;
#10;x=75110000;
#10;x=75120000;
#10;x=75130000;
#10;x=75140000;
#10;x=75150000;
#10;x=75160000;
#10;x=75170000;
#10;x=75180000;
#10;x=75190000;
#10;x=75200000;
#10;x=75210000;
#10;x=75220000;
#10;x=75230000;
#10;x=75240000;
#10;x=75250000;
#10;x=75260000;
#10;x=75270000;
#10;x=75280000;
#10;x=75290000;
#10;x=75300000;
#10;x=75310000;
#10;x=75320000;
#10;x=75330000;
#10;x=75340000;
#10;x=75350000;
#10;x=75360000;
#10;x=75370000;
#10;x=75380000;
#10;x=75390000;
#10;x=75400000;
#10;x=75410000;
#10;x=75420000;
#10;x=75430000;
#10;x=75440000;
#10;x=75450000;
#10;x=75460000;
#10;x=75470000;
#10;x=75480000;
#10;x=75490000;
#10;x=75500000;
#10;x=75510000;
#10;x=75520000;
#10;x=75530000;
#10;x=75540000;
#10;x=75550000;
#10;x=75560000;
#10;x=75570000;
#10;x=75580000;
#10;x=75590000;
#10;x=75600000;
#10;x=75610000;
#10;x=75620000;
#10;x=75630000;
#10;x=75640000;
#10;x=75650000;
#10;x=75660000;
#10;x=75670000;
#10;x=75680000;
#10;x=75690000;
#10;x=75700000;
#10;x=75710000;
#10;x=75720000;
#10;x=75730000;
#10;x=75740000;
#10;x=75750000;
#10;x=75760000;
#10;x=75770000;
#10;x=75780000;
#10;x=75790000;
#10;x=75800000;
#10;x=75810000;
#10;x=75820000;
#10;x=75830000;
#10;x=75840000;
#10;x=75850000;
#10;x=75860000;
#10;x=75870000;
#10;x=75880000;
#10;x=75890000;
#10;x=75900000;
#10;x=75910000;
#10;x=75920000;
#10;x=75930000;
#10;x=75940000;
#10;x=75950000;
#10;x=75960000;
#10;x=75970000;
#10;x=75980000;
#10;x=75990000;
#10;x=76000000;
#10;x=76010000;
#10;x=76020000;
#10;x=76030000;
#10;x=76040000;
#10;x=76050000;
#10;x=76060000;
#10;x=76070000;
#10;x=76080000;
#10;x=76090000;
#10;x=76100000;
#10;x=76110000;
#10;x=76120000;
#10;x=76130000;
#10;x=76140000;
#10;x=76150000;
#10;x=76160000;
#10;x=76170000;
#10;x=76180000;
#10;x=76190000;
#10;x=76200000;
#10;x=76210000;
#10;x=76220000;
#10;x=76230000;
#10;x=76240000;
#10;x=76250000;
#10;x=76260000;
#10;x=76270000;
#10;x=76280000;
#10;x=76290000;
#10;x=76300000;
#10;x=76310000;
#10;x=76320000;
#10;x=76330000;
#10;x=76340000;
#10;x=76350000;
#10;x=76360000;
#10;x=76370000;
#10;x=76380000;
#10;x=76390000;
#10;x=76400000;
#10;x=76410000;
#10;x=76420000;
#10;x=76430000;
#10;x=76440000;
#10;x=76450000;
#10;x=76460000;
#10;x=76470000;
#10;x=76480000;
#10;x=76490000;
#10;x=76500000;
#10;x=76510000;
#10;x=76520000;
#10;x=76530000;
#10;x=76540000;
#10;x=76550000;
#10;x=76560000;
#10;x=76570000;
#10;x=76580000;
#10;x=76590000;
#10;x=76600000;
#10;x=76610000;
#10;x=76620000;
#10;x=76630000;
#10;x=76640000;
#10;x=76650000;
#10;x=76660000;
#10;x=76670000;
#10;x=76680000;
#10;x=76690000;
#10;x=76700000;
#10;x=76710000;
#10;x=76720000;
#10;x=76730000;
#10;x=76740000;
#10;x=76750000;
#10;x=76760000;
#10;x=76770000;
#10;x=76780000;
#10;x=76790000;
#10;x=76800000;
#10;x=76810000;
#10;x=76820000;
#10;x=76830000;
#10;x=76840000;
#10;x=76850000;
#10;x=76860000;
#10;x=76870000;
#10;x=76880000;
#10;x=76890000;
#10;x=76900000;
#10;x=76910000;
#10;x=76920000;
#10;x=76930000;
#10;x=76940000;
#10;x=76950000;
#10;x=76960000;
#10;x=76970000;
#10;x=76980000;
#10;x=76990000;
#10;x=77000000;
#10;x=77010000;
#10;x=77020000;
#10;x=77030000;
#10;x=77040000;
#10;x=77050000;
#10;x=77060000;
#10;x=77070000;
#10;x=77080000;
#10;x=77090000;
#10;x=77100000;
#10;x=77110000;
#10;x=77120000;
#10;x=77130000;
#10;x=77140000;
#10;x=77150000;
#10;x=77160000;
#10;x=77170000;
#10;x=77180000;
#10;x=77190000;
#10;x=77200000;
#10;x=77210000;
#10;x=77220000;
#10;x=77230000;
#10;x=77240000;
#10;x=77250000;
#10;x=77260000;
#10;x=77270000;
#10;x=77280000;
#10;x=77290000;
#10;x=77300000;
#10;x=77310000;
#10;x=77320000;
#10;x=77330000;
#10;x=77340000;
#10;x=77350000;
#10;x=77360000;
#10;x=77370000;
#10;x=77380000;
#10;x=77390000;
#10;x=77400000;
#10;x=77410000;
#10;x=77420000;
#10;x=77430000;
#10;x=77440000;
#10;x=77450000;
#10;x=77460000;
#10;x=77470000;
#10;x=77480000;
#10;x=77490000;
#10;x=77500000;
#10;x=77510000;
#10;x=77520000;
#10;x=77530000;
#10;x=77540000;
#10;x=77550000;
#10;x=77560000;
#10;x=77570000;
#10;x=77580000;
#10;x=77590000;
#10;x=77600000;
#10;x=77610000;
#10;x=77620000;
#10;x=77630000;
#10;x=77640000;
#10;x=77650000;
#10;x=77660000;
#10;x=77670000;
#10;x=77680000;
#10;x=77690000;
#10;x=77700000;
#10;x=77710000;
#10;x=77720000;
#10;x=77730000;
#10;x=77740000;
#10;x=77750000;
#10;x=77760000;
#10;x=77770000;
#10;x=77780000;
#10;x=77790000;
#10;x=77800000;
#10;x=77810000;
#10;x=77820000;
#10;x=77830000;
#10;x=77840000;
#10;x=77850000;
#10;x=77860000;
#10;x=77870000;
#10;x=77880000;
#10;x=77890000;
#10;x=77900000;
#10;x=77910000;
#10;x=77920000;
#10;x=77930000;
#10;x=77940000;
#10;x=77950000;
#10;x=77960000;
#10;x=77970000;
#10;x=77980000;
#10;x=77990000;
#10;x=78000000;
#10;x=78010000;
#10;x=78020000;
#10;x=78030000;
#10;x=78040000;
#10;x=78050000;
#10;x=78060000;
#10;x=78070000;
#10;x=78080000;
#10;x=78090000;
#10;x=78100000;
#10;x=78110000;
#10;x=78120000;
#10;x=78130000;
#10;x=78140000;
#10;x=78150000;
#10;x=78160000;
#10;x=78170000;
#10;x=78180000;
#10;x=78190000;
#10;x=78200000;
#10;x=78210000;
#10;x=78220000;
#10;x=78230000;
#10;x=78240000;
#10;x=78250000;
#10;x=78260000;
#10;x=78270000;
#10;x=78280000;
#10;x=78290000;
#10;x=78300000;
#10;x=78310000;
#10;x=78320000;
#10;x=78330000;
#10;x=78340000;
#10;x=78350000;
#10;x=78360000;
#10;x=78370000;
#10;x=78380000;
#10;x=78390000;
#10;x=78400000;
#10;x=78410000;
#10;x=78420000;
#10;x=78430000;
#10;x=78440000;
#10;x=78450000;
#10;x=78460000;
#10;x=78470000;
#10;x=78480000;
#10;x=78490000;
#10;x=78500000;
#10;x=78510000;
#10;x=78520000;
#10;x=78530000;
#10;x=78540000;
#10;x=78550000;
#10;x=78560000;
#10;x=78570000;
#10;x=78580000;
#10;x=78590000;
#10;x=78600000;
#10;x=78610000;
#10;x=78620000;
#10;x=78630000;
#10;x=78640000;
#10;x=78650000;
#10;x=78660000;
#10;x=78670000;
#10;x=78680000;
#10;x=78690000;
#10;x=78700000;
#10;x=78710000;
#10;x=78720000;
#10;x=78730000;
#10;x=78740000;
#10;x=78750000;
#10;x=78760000;
#10;x=78770000;
#10;x=78780000;
#10;x=78790000;
#10;x=78800000;
#10;x=78810000;
#10;x=78820000;
#10;x=78830000;
#10;x=78840000;
#10;x=78850000;
#10;x=78860000;
#10;x=78870000;
#10;x=78880000;
#10;x=78890000;
#10;x=78900000;
#10;x=78910000;
#10;x=78920000;
#10;x=78930000;
#10;x=78940000;
#10;x=78950000;
#10;x=78960000;
#10;x=78970000;
#10;x=78980000;
#10;x=78990000;
#10;x=79000000;
#10;x=79010000;
#10;x=79020000;
#10;x=79030000;
#10;x=79040000;
#10;x=79050000;
#10;x=79060000;
#10;x=79070000;
#10;x=79080000;
#10;x=79090000;
#10;x=79100000;
#10;x=79110000;
#10;x=79120000;
#10;x=79130000;
#10;x=79140000;
#10;x=79150000;
#10;x=79160000;
#10;x=79170000;
#10;x=79180000;
#10;x=79190000;
#10;x=79200000;
#10;x=79210000;
#10;x=79220000;
#10;x=79230000;
#10;x=79240000;
#10;x=79250000;
#10;x=79260000;
#10;x=79270000;
#10;x=79280000;
#10;x=79290000;
#10;x=79300000;
#10;x=79310000;
#10;x=79320000;
#10;x=79330000;
#10;x=79340000;
#10;x=79350000;
#10;x=79360000;
#10;x=79370000;
#10;x=79380000;
#10;x=79390000;
#10;x=79400000;
#10;x=79410000;
#10;x=79420000;
#10;x=79430000;
#10;x=79440000;
#10;x=79450000;
#10;x=79460000;
#10;x=79470000;
#10;x=79480000;
#10;x=79490000;
#10;x=79500000;
#10;x=79510000;
#10;x=79520000;
#10;x=79530000;
#10;x=79540000;
#10;x=79550000;
#10;x=79560000;
#10;x=79570000;
#10;x=79580000;
#10;x=79590000;
#10;x=79600000;
#10;x=79610000;
#10;x=79620000;
#10;x=79630000;
#10;x=79640000;
#10;x=79650000;
#10;x=79660000;
#10;x=79670000;
#10;x=79680000;
#10;x=79690000;
#10;x=79700000;
#10;x=79710000;
#10;x=79720000;
#10;x=79730000;
#10;x=79740000;
#10;x=79750000;
#10;x=79760000;
#10;x=79770000;
#10;x=79780000;
#10;x=79790000;
#10;x=79800000;
#10;x=79810000;
#10;x=79820000;
#10;x=79830000;
#10;x=79840000;
#10;x=79850000;
#10;x=79860000;
#10;x=79870000;
#10;x=79880000;
#10;x=79890000;
#10;x=79900000;
#10;x=79910000;
#10;x=79920000;
#10;x=79930000;
#10;x=79940000;
#10;x=79950000;
#10;x=79960000;
#10;x=79970000;
#10;x=79980000;
#10;x=79990000;
#10;x=80000000;
#10;x=80010000;
#10;x=80020000;
#10;x=80030000;
#10;x=80040000;
#10;x=80050000;
#10;x=80060000;
#10;x=80070000;
#10;x=80080000;
#10;x=80090000;
#10;x=80100000;
#10;x=80110000;
#10;x=80120000;
#10;x=80130000;
#10;x=80140000;
#10;x=80150000;
#10;x=80160000;
#10;x=80170000;
#10;x=80180000;
#10;x=80190000;
#10;x=80200000;
#10;x=80210000;
#10;x=80220000;
#10;x=80230000;
#10;x=80240000;
#10;x=80250000;
#10;x=80260000;
#10;x=80270000;
#10;x=80280000;
#10;x=80290000;
#10;x=80300000;
#10;x=80310000;
#10;x=80320000;
#10;x=80330000;
#10;x=80340000;
#10;x=80350000;
#10;x=80360000;
#10;x=80370000;
#10;x=80380000;
#10;x=80390000;
#10;x=80400000;
#10;x=80410000;
#10;x=80420000;
#10;x=80430000;
#10;x=80440000;
#10;x=80450000;
#10;x=80460000;
#10;x=80470000;
#10;x=80480000;
#10;x=80490000;
#10;x=80500000;
#10;x=80510000;
#10;x=80520000;
#10;x=80530000;
#10;x=80540000;
#10;x=80550000;
#10;x=80560000;
#10;x=80570000;
#10;x=80580000;
#10;x=80590000;
#10;x=80600000;
#10;x=80610000;
#10;x=80620000;
#10;x=80630000;
#10;x=80640000;
#10;x=80650000;
#10;x=80660000;
#10;x=80670000;
#10;x=80680000;
#10;x=80690000;
#10;x=80700000;
#10;x=80710000;
#10;x=80720000;
#10;x=80730000;
#10;x=80740000;
#10;x=80750000;
#10;x=80760000;
#10;x=80770000;
#10;x=80780000;
#10;x=80790000;
#10;x=80800000;
#10;x=80810000;
#10;x=80820000;
#10;x=80830000;
#10;x=80840000;
#10;x=80850000;
#10;x=80860000;
#10;x=80870000;
#10;x=80880000;
#10;x=80890000;
#10;x=80900000;
#10;x=80910000;
#10;x=80920000;
#10;x=80930000;
#10;x=80940000;
#10;x=80950000;
#10;x=80960000;
#10;x=80970000;
#10;x=80980000;
#10;x=80990000;
#10;x=81000000;
#10;x=81010000;
#10;x=81020000;
#10;x=81030000;
#10;x=81040000;
#10;x=81050000;
#10;x=81060000;
#10;x=81070000;
#10;x=81080000;
#10;x=81090000;
#10;x=81100000;
#10;x=81110000;
#10;x=81120000;
#10;x=81130000;
#10;x=81140000;
#10;x=81150000;
#10;x=81160000;
#10;x=81170000;
#10;x=81180000;
#10;x=81190000;
#10;x=81200000;
#10;x=81210000;
#10;x=81220000;
#10;x=81230000;
#10;x=81240000;
#10;x=81250000;
#10;x=81260000;
#10;x=81270000;
#10;x=81280000;
#10;x=81290000;
#10;x=81300000;
#10;x=81310000;
#10;x=81320000;
#10;x=81330000;
#10;x=81340000;
#10;x=81350000;
#10;x=81360000;
#10;x=81370000;
#10;x=81380000;
#10;x=81390000;
#10;x=81400000;
#10;x=81410000;
#10;x=81420000;
#10;x=81430000;
#10;x=81440000;
#10;x=81450000;
#10;x=81460000;
#10;x=81470000;
#10;x=81480000;
#10;x=81490000;
#10;x=81500000;
#10;x=81510000;
#10;x=81520000;
#10;x=81530000;
#10;x=81540000;
#10;x=81550000;
#10;x=81560000;
#10;x=81570000;
#10;x=81580000;
#10;x=81590000;
#10;x=81600000;
#10;x=81610000;
#10;x=81620000;
#10;x=81630000;
#10;x=81640000;
#10;x=81650000;
#10;x=81660000;
#10;x=81670000;
#10;x=81680000;
#10;x=81690000;
#10;x=81700000;
#10;x=81710000;
#10;x=81720000;
#10;x=81730000;
#10;x=81740000;
#10;x=81750000;
#10;x=81760000;
#10;x=81770000;
#10;x=81780000;
#10;x=81790000;
#10;x=81800000;
#10;x=81810000;
#10;x=81820000;
#10;x=81830000;
#10;x=81840000;
#10;x=81850000;
#10;x=81860000;
#10;x=81870000;
#10;x=81880000;
#10;x=81890000;
#10;x=81900000;
#10;x=81910000;
#10;x=81920000;
#10;x=81930000;
#10;x=81940000;
#10;x=81950000;
#10;x=81960000;
#10;x=81970000;
#10;x=81980000;
#10;x=81990000;
#10;x=82000000;
#10;x=82010000;
#10;x=82020000;
#10;x=82030000;
#10;x=82040000;
#10;x=82050000;
#10;x=82060000;
#10;x=82070000;
#10;x=82080000;
#10;x=82090000;
#10;x=82100000;
#10;x=82110000;
#10;x=82120000;
#10;x=82130000;
#10;x=82140000;
#10;x=82150000;
#10;x=82160000;
#10;x=82170000;
#10;x=82180000;
#10;x=82190000;
#10;x=82200000;
#10;x=82210000;
#10;x=82220000;
#10;x=82230000;
#10;x=82240000;
#10;x=82250000;
#10;x=82260000;
#10;x=82270000;
#10;x=82280000;
#10;x=82290000;
#10;x=82300000;
#10;x=82310000;
#10;x=82320000;
#10;x=82330000;
#10;x=82340000;
#10;x=82350000;
#10;x=82360000;
#10;x=82370000;
#10;x=82380000;
#10;x=82390000;
#10;x=82400000;
#10;x=82410000;
#10;x=82420000;
#10;x=82430000;
#10;x=82440000;
#10;x=82450000;
#10;x=82460000;
#10;x=82470000;
#10;x=82480000;
#10;x=82490000;
#10;x=82500000;
#10;x=82510000;
#10;x=82520000;
#10;x=82530000;
#10;x=82540000;
#10;x=82550000;
#10;x=82560000;
#10;x=82570000;
#10;x=82580000;
#10;x=82590000;
#10;x=82600000;
#10;x=82610000;
#10;x=82620000;
#10;x=82630000;
#10;x=82640000;
#10;x=82650000;
#10;x=82660000;
#10;x=82670000;
#10;x=82680000;
#10;x=82690000;
#10;x=82700000;
#10;x=82710000;
#10;x=82720000;
#10;x=82730000;
#10;x=82740000;
#10;x=82750000;
#10;x=82760000;
#10;x=82770000;
#10;x=82780000;
#10;x=82790000;
#10;x=82800000;
#10;x=82810000;
#10;x=82820000;
#10;x=82830000;
#10;x=82840000;
#10;x=82850000;
#10;x=82860000;
#10;x=82870000;
#10;x=82880000;
#10;x=82890000;
#10;x=82900000;
#10;x=82910000;
#10;x=82920000;
#10;x=82930000;
#10;x=82940000;
#10;x=82950000;
#10;x=82960000;
#10;x=82970000;
#10;x=82980000;
#10;x=82990000;
#10;x=83000000;
#10;x=83010000;
#10;x=83020000;
#10;x=83030000;
#10;x=83040000;
#10;x=83050000;
#10;x=83060000;
#10;x=83070000;
#10;x=83080000;
#10;x=83090000;
#10;x=83100000;
#10;x=83110000;
#10;x=83120000;
#10;x=83130000;
#10;x=83140000;
#10;x=83150000;
#10;x=83160000;
#10;x=83170000;
#10;x=83180000;
#10;x=83190000;
#10;x=83200000;
#10;x=83210000;
#10;x=83220000;
#10;x=83230000;
#10;x=83240000;
#10;x=83250000;
#10;x=83260000;
#10;x=83270000;
#10;x=83280000;
#10;x=83290000;
#10;x=83300000;
#10;x=83310000;
#10;x=83320000;
#10;x=83330000;
#10;x=83340000;
#10;x=83350000;
#10;x=83360000;
#10;x=83370000;
#10;x=83380000;
#10;x=83390000;
#10;x=83400000;
#10;x=83410000;
#10;x=83420000;
#10;x=83430000;
#10;x=83440000;
#10;x=83450000;
#10;x=83460000;
#10;x=83470000;
#10;x=83480000;
#10;x=83490000;
#10;x=83500000;
#10;x=83510000;
#10;x=83520000;
#10;x=83530000;
#10;x=83540000;
#10;x=83550000;
#10;x=83560000;
#10;x=83570000;
#10;x=83580000;
#10;x=83590000;
#10;x=83600000;
#10;x=83610000;
#10;x=83620000;
#10;x=83630000;
#10;x=83640000;
#10;x=83650000;
#10;x=83660000;
#10;x=83670000;
#10;x=83680000;
#10;x=83690000;
#10;x=83700000;
#10;x=83710000;
#10;x=83720000;
#10;x=83730000;
#10;x=83740000;
#10;x=83750000;
#10;x=83760000;
#10;x=83770000;
#10;x=83780000;
#10;x=83790000;
#10;x=83800000;
#10;x=83810000;
#10;x=83820000;
#10;x=83830000;
#10;x=83840000;
#10;x=83850000;
#10;x=83860000;
#10;x=83870000;
#10;x=83880000;
#10;x=83890000;
#10;x=83900000;
#10;x=83910000;
#10;x=83920000;
#10;x=83930000;
#10;x=83940000;
#10;x=83950000;
#10;x=83960000;
#10;x=83970000;
#10;x=83980000;
#10;x=83990000;
#10;x=84000000;
#10;x=84010000;
#10;x=84020000;
#10;x=84030000;
#10;x=84040000;
#10;x=84050000;
#10;x=84060000;
#10;x=84070000;
#10;x=84080000;
#10;x=84090000;
#10;x=84100000;
#10;x=84110000;
#10;x=84120000;
#10;x=84130000;
#10;x=84140000;
#10;x=84150000;
#10;x=84160000;
#10;x=84170000;
#10;x=84180000;
#10;x=84190000;
#10;x=84200000;
#10;x=84210000;
#10;x=84220000;
#10;x=84230000;
#10;x=84240000;
#10;x=84250000;
#10;x=84260000;
#10;x=84270000;
#10;x=84280000;
#10;x=84290000;
#10;x=84300000;
#10;x=84310000;
#10;x=84320000;
#10;x=84330000;
#10;x=84340000;
#10;x=84350000;
#10;x=84360000;
#10;x=84370000;
#10;x=84380000;
#10;x=84390000;
#10;x=84400000;
#10;x=84410000;
#10;x=84420000;
#10;x=84430000;
#10;x=84440000;
#10;x=84450000;
#10;x=84460000;
#10;x=84470000;
#10;x=84480000;
#10;x=84490000;
#10;x=84500000;
#10;x=84510000;
#10;x=84520000;
#10;x=84530000;
#10;x=84540000;
#10;x=84550000;
#10;x=84560000;
#10;x=84570000;
#10;x=84580000;
#10;x=84590000;
#10;x=84600000;
#10;x=84610000;
#10;x=84620000;
#10;x=84630000;
#10;x=84640000;
#10;x=84650000;
#10;x=84660000;
#10;x=84670000;
#10;x=84680000;
#10;x=84690000;
#10;x=84700000;
#10;x=84710000;
#10;x=84720000;
#10;x=84730000;
#10;x=84740000;
#10;x=84750000;
#10;x=84760000;
#10;x=84770000;
#10;x=84780000;
#10;x=84790000;
#10;x=84800000;
#10;x=84810000;
#10;x=84820000;
#10;x=84830000;
#10;x=84840000;
#10;x=84850000;
#10;x=84860000;
#10;x=84870000;
#10;x=84880000;
#10;x=84890000;
#10;x=84900000;
#10;x=84910000;
#10;x=84920000;
#10;x=84930000;
#10;x=84940000;
#10;x=84950000;
#10;x=84960000;
#10;x=84970000;
#10;x=84980000;
#10;x=84990000;
#10;x=85000000;
#10;x=85010000;
#10;x=85020000;
#10;x=85030000;
#10;x=85040000;
#10;x=85050000;
#10;x=85060000;
#10;x=85070000;
#10;x=85080000;
#10;x=85090000;
#10;x=85100000;
#10;x=85110000;
#10;x=85120000;
#10;x=85130000;
#10;x=85140000;
#10;x=85150000;
#10;x=85160000;
#10;x=85170000;
#10;x=85180000;
#10;x=85190000;
#10;x=85200000;
#10;x=85210000;
#10;x=85220000;
#10;x=85230000;
#10;x=85240000;
#10;x=85250000;
#10;x=85260000;
#10;x=85270000;
#10;x=85280000;
#10;x=85290000;
#10;x=85300000;
#10;x=85310000;
#10;x=85320000;
#10;x=85330000;
#10;x=85340000;
#10;x=85350000;
#10;x=85360000;
#10;x=85370000;
#10;x=85380000;
#10;x=85390000;
#10;x=85400000;
#10;x=85410000;
#10;x=85420000;
#10;x=85430000;
#10;x=85440000;
#10;x=85450000;
#10;x=85460000;
#10;x=85470000;
#10;x=85480000;
#10;x=85490000;
#10;x=85500000;
#10;x=85510000;
#10;x=85520000;
#10;x=85530000;
#10;x=85540000;
#10;x=85550000;
#10;x=85560000;
#10;x=85570000;
#10;x=85580000;
#10;x=85590000;
#10;x=85600000;
#10;x=85610000;
#10;x=85620000;
#10;x=85630000;
#10;x=85640000;
#10;x=85650000;
#10;x=85660000;
#10;x=85670000;
#10;x=85680000;
#10;x=85690000;
#10;x=85700000;
#10;x=85710000;
#10;x=85720000;
#10;x=85730000;
#10;x=85740000;
#10;x=85750000;
#10;x=85760000;
#10;x=85770000;
#10;x=85780000;
#10;x=85790000;
#10;x=85800000;
#10;x=85810000;
#10;x=85820000;
#10;x=85830000;
#10;x=85840000;
#10;x=85850000;
#10;x=85860000;
#10;x=85870000;
#10;x=85880000;
#10;x=85890000;
#10;x=85900000;
#10;x=85910000;
#10;x=85920000;
#10;x=85930000;
#10;x=85940000;
#10;x=85950000;
#10;x=85960000;
#10;x=85970000;
#10;x=85980000;
#10;x=85990000;
#10;x=86000000;
#10;x=86010000;
#10;x=86020000;
#10;x=86030000;
#10;x=86040000;
#10;x=86050000;
#10;x=86060000;
#10;x=86070000;
#10;x=86080000;
#10;x=86090000;
#10;x=86100000;
#10;x=86110000;
#10;x=86120000;
#10;x=86130000;
#10;x=86140000;
#10;x=86150000;
#10;x=86160000;
#10;x=86170000;
#10;x=86180000;
#10;x=86190000;
#10;x=86200000;
#10;x=86210000;
#10;x=86220000;
#10;x=86230000;
#10;x=86240000;
#10;x=86250000;
#10;x=86260000;
#10;x=86270000;
#10;x=86280000;
#10;x=86290000;
#10;x=86300000;
#10;x=86310000;
#10;x=86320000;
#10;x=86330000;
#10;x=86340000;
#10;x=86350000;
#10;x=86360000;
#10;x=86370000;
#10;x=86380000;
#10;x=86390000;
#10;x=86400000;
#10;x=86410000;
#10;x=86420000;
#10;x=86430000;
#10;x=86440000;
#10;x=86450000;
#10;x=86460000;
#10;x=86470000;
#10;x=86480000;
#10;x=86490000;
#10;x=86500000;
#10;x=86510000;
#10;x=86520000;
#10;x=86530000;
#10;x=86540000;
#10;x=86550000;
#10;x=86560000;
#10;x=86570000;
#10;x=86580000;
#10;x=86590000;
#10;x=86600000;
#10;x=86610000;
#10;x=86620000;
#10;x=86630000;
#10;x=86640000;
#10;x=86650000;
#10;x=86660000;
#10;x=86670000;
#10;x=86680000;
#10;x=86690000;
#10;x=86700000;
#10;x=86710000;
#10;x=86720000;
#10;x=86730000;
#10;x=86740000;
#10;x=86750000;
#10;x=86760000;
#10;x=86770000;
#10;x=86780000;
#10;x=86790000;
#10;x=86800000;
#10;x=86810000;
#10;x=86820000;
#10;x=86830000;
#10;x=86840000;
#10;x=86850000;
#10;x=86860000;
#10;x=86870000;
#10;x=86880000;
#10;x=86890000;
#10;x=86900000;
#10;x=86910000;
#10;x=86920000;
#10;x=86930000;
#10;x=86940000;
#10;x=86950000;
#10;x=86960000;
#10;x=86970000;
#10;x=86980000;
#10;x=86990000;
#10;x=87000000;
#10;x=87010000;
#10;x=87020000;
#10;x=87030000;
#10;x=87040000;
#10;x=87050000;
#10;x=87060000;
#10;x=87070000;
#10;x=87080000;
#10;x=87090000;
#10;x=87100000;
#10;x=87110000;
#10;x=87120000;
#10;x=87130000;
#10;x=87140000;
#10;x=87150000;
#10;x=87160000;
#10;x=87170000;
#10;x=87180000;
#10;x=87190000;
#10;x=87200000;
#10;x=87210000;
#10;x=87220000;
#10;x=87230000;
#10;x=87240000;
#10;x=87250000;
#10;x=87260000;
#10;x=87270000;
#10;x=87280000;
#10;x=87290000;
#10;x=87300000;
#10;x=87310000;
#10;x=87320000;
#10;x=87330000;
#10;x=87340000;
#10;x=87350000;
#10;x=87360000;
#10;x=87370000;
#10;x=87380000;
#10;x=87390000;
#10;x=87400000;
#10;x=87410000;
#10;x=87420000;
#10;x=87430000;
#10;x=87440000;
#10;x=87450000;
#10;x=87460000;
#10;x=87470000;
#10;x=87480000;
#10;x=87490000;
#10;x=87500000;
#10;x=87510000;
#10;x=87520000;
#10;x=87530000;
#10;x=87540000;
#10;x=87550000;
#10;x=87560000;
#10;x=87570000;
#10;x=87580000;
#10;x=87590000;
#10;x=87600000;
#10;x=87610000;
#10;x=87620000;
#10;x=87630000;
#10;x=87640000;
#10;x=87650000;
#10;x=87660000;
#10;x=87670000;
#10;x=87680000;
#10;x=87690000;
#10;x=87700000;
#10;x=87710000;
#10;x=87720000;
#10;x=87730000;
#10;x=87740000;
#10;x=87750000;
#10;x=87760000;
#10;x=87770000;
#10;x=87780000;
#10;x=87790000;
#10;x=87800000;
#10;x=87810000;
#10;x=87820000;
#10;x=87830000;
#10;x=87840000;
#10;x=87850000;
#10;x=87860000;
#10;x=87870000;
#10;x=87880000;
#10;x=87890000;
#10;x=87900000;
#10;x=87910000;
#10;x=87920000;
#10;x=87930000;
#10;x=87940000;
#10;x=87950000;
#10;x=87960000;
#10;x=87970000;
#10;x=87980000;
#10;x=87990000;
#10;x=88000000;
#10;x=88010000;
#10;x=88020000;
#10;x=88030000;
#10;x=88040000;
#10;x=88050000;
#10;x=88060000;
#10;x=88070000;
#10;x=88080000;
#10;x=88090000;
#10;x=88100000;
#10;x=88110000;
#10;x=88120000;
#10;x=88130000;
#10;x=88140000;
#10;x=88150000;
#10;x=88160000;
#10;x=88170000;
#10;x=88180000;
#10;x=88190000;
#10;x=88200000;
#10;x=88210000;
#10;x=88220000;
#10;x=88230000;
#10;x=88240000;
#10;x=88250000;
#10;x=88260000;
#10;x=88270000;
#10;x=88280000;
#10;x=88290000;
#10;x=88300000;
#10;x=88310000;
#10;x=88320000;
#10;x=88330000;
#10;x=88340000;
#10;x=88350000;
#10;x=88360000;
#10;x=88370000;
#10;x=88380000;
#10;x=88390000;
#10;x=88400000;
#10;x=88410000;
#10;x=88420000;
#10;x=88430000;
#10;x=88440000;
#10;x=88450000;
#10;x=88460000;
#10;x=88470000;
#10;x=88480000;
#10;x=88490000;
#10;x=88500000;
#10;x=88510000;
#10;x=88520000;
#10;x=88530000;
#10;x=88540000;
#10;x=88550000;
#10;x=88560000;
#10;x=88570000;
#10;x=88580000;
#10;x=88590000;
#10;x=88600000;
#10;x=88610000;
#10;x=88620000;
#10;x=88630000;
#10;x=88640000;
#10;x=88650000;
#10;x=88660000;
#10;x=88670000;
#10;x=88680000;
#10;x=88690000;
#10;x=88700000;
#10;x=88710000;
#10;x=88720000;
#10;x=88730000;
#10;x=88740000;
#10;x=88750000;
#10;x=88760000;
#10;x=88770000;
#10;x=88780000;
#10;x=88790000;
#10;x=88800000;
#10;x=88810000;
#10;x=88820000;
#10;x=88830000;
#10;x=88840000;
#10;x=88850000;
#10;x=88860000;
#10;x=88870000;
#10;x=88880000;
#10;x=88890000;
#10;x=88900000;
#10;x=88910000;
#10;x=88920000;
#10;x=88930000;
#10;x=88940000;
#10;x=88950000;
#10;x=88960000;
#10;x=88970000;
#10;x=88980000;
#10;x=88990000;
#10;x=89000000;
#10;x=89010000;
#10;x=89020000;
#10;x=89030000;
#10;x=89040000;
#10;x=89050000;
#10;x=89060000;
#10;x=89070000;
#10;x=89080000;
#10;x=89090000;
#10;x=89100000;
#10;x=89110000;
#10;x=89120000;
#10;x=89130000;
#10;x=89140000;
#10;x=89150000;
#10;x=89160000;
#10;x=89170000;
#10;x=89180000;
#10;x=89190000;
#10;x=89200000;
#10;x=89210000;
#10;x=89220000;
#10;x=89230000;
#10;x=89240000;
#10;x=89250000;
#10;x=89260000;
#10;x=89270000;
#10;x=89280000;
#10;x=89290000;
#10;x=89300000;
#10;x=89310000;
#10;x=89320000;
#10;x=89330000;
#10;x=89340000;
#10;x=89350000;
#10;x=89360000;
#10;x=89370000;
#10;x=89380000;
#10;x=89390000;
#10;x=89400000;
#10;x=89410000;
#10;x=89420000;
#10;x=89430000;
#10;x=89440000;
#10;x=89450000;
#10;x=89460000;
#10;x=89470000;
#10;x=89480000;
#10;x=89490000;
#10;x=89500000;
#10;x=89510000;
#10;x=89520000;
#10;x=89530000;
#10;x=89540000;
#10;x=89550000;
#10;x=89560000;
#10;x=89570000;
#10;x=89580000;
#10;x=89590000;
#10;x=89600000;
#10;x=89610000;
#10;x=89620000;
#10;x=89630000;
#10;x=89640000;
#10;x=89650000;
#10;x=89660000;
#10;x=89670000;
#10;x=89680000;
#10;x=89690000;
#10;x=89700000;
#10;x=89710000;
#10;x=89720000;
#10;x=89730000;
#10;x=89740000;
#10;x=89750000;
#10;x=89760000;
#10;x=89770000;
#10;x=89780000;
#10;x=89790000;
#10;x=89800000;
#10;x=89810000;
#10;x=89820000;
#10;x=89830000;
#10;x=89840000;
#10;x=89850000;
#10;x=89860000;
#10;x=89870000;
#10;x=89880000;
#10;x=89890000;
#10;x=89900000;
#10;x=89910000;
#10;x=89920000;
#10;x=89930000;
#10;x=89940000;
#10;x=89950000;
#10;x=89960000;
#10;x=89970000;
#10;x=89980000;
#10;x=89990000;
#10;x=90000000;
#10;x=90010000;
#10;x=90020000;
#10;x=90030000;
#10;x=90040000;
#10;x=90050000;
#10;x=90060000;
#10;x=90070000;
#10;x=90080000;
#10;x=90090000;
#10;x=90100000;
#10;x=90110000;
#10;x=90120000;
#10;x=90130000;
#10;x=90140000;
#10;x=90150000;
#10;x=90160000;
#10;x=90170000;
#10;x=90180000;
#10;x=90190000;
#10;x=90200000;
#10;x=90210000;
#10;x=90220000;
#10;x=90230000;
#10;x=90240000;
#10;x=90250000;
#10;x=90260000;
#10;x=90270000;
#10;x=90280000;
#10;x=90290000;
#10;x=90300000;
#10;x=90310000;
#10;x=90320000;
#10;x=90330000;
#10;x=90340000;
#10;x=90350000;
#10;x=90360000;
#10;x=90370000;
#10;x=90380000;
#10;x=90390000;
#10;x=90400000;
#10;x=90410000;
#10;x=90420000;
#10;x=90430000;
#10;x=90440000;
#10;x=90450000;
#10;x=90460000;
#10;x=90470000;
#10;x=90480000;
#10;x=90490000;
#10;x=90500000;
#10;x=90510000;
#10;x=90520000;
#10;x=90530000;
#10;x=90540000;
#10;x=90550000;
#10;x=90560000;
#10;x=90570000;
#10;x=90580000;
#10;x=90590000;
#10;x=90600000;
#10;x=90610000;
#10;x=90620000;
#10;x=90630000;
#10;x=90640000;
#10;x=90650000;
#10;x=90660000;
#10;x=90670000;
#10;x=90680000;
#10;x=90690000;
#10;x=90700000;
#10;x=90710000;
#10;x=90720000;
#10;x=90730000;
#10;x=90740000;
#10;x=90750000;
#10;x=90760000;
#10;x=90770000;
#10;x=90780000;
#10;x=90790000;
#10;x=90800000;
#10;x=90810000;
#10;x=90820000;
#10;x=90830000;
#10;x=90840000;
#10;x=90850000;
#10;x=90860000;
#10;x=90870000;
#10;x=90880000;
#10;x=90890000;
#10;x=90900000;
#10;x=90910000;
#10;x=90920000;
#10;x=90930000;
#10;x=90940000;
#10;x=90950000;
#10;x=90960000;
#10;x=90970000;
#10;x=90980000;
#10;x=90990000;
#10;x=91000000;
#10;x=91010000;
#10;x=91020000;
#10;x=91030000;
#10;x=91040000;
#10;x=91050000;
#10;x=91060000;
#10;x=91070000;
#10;x=91080000;
#10;x=91090000;
#10;x=91100000;
#10;x=91110000;
#10;x=91120000;
#10;x=91130000;
#10;x=91140000;
#10;x=91150000;
#10;x=91160000;
#10;x=91170000;
#10;x=91180000;
#10;x=91190000;
#10;x=91200000;
#10;x=91210000;
#10;x=91220000;
#10;x=91230000;
#10;x=91240000;
#10;x=91250000;
#10;x=91260000;
#10;x=91270000;
#10;x=91280000;
#10;x=91290000;
#10;x=91300000;
#10;x=91310000;
#10;x=91320000;
#10;x=91330000;
#10;x=91340000;
#10;x=91350000;
#10;x=91360000;
#10;x=91370000;
#10;x=91380000;
#10;x=91390000;
#10;x=91400000;
#10;x=91410000;
#10;x=91420000;
#10;x=91430000;
#10;x=91440000;
#10;x=91450000;
#10;x=91460000;
#10;x=91470000;
#10;x=91480000;
#10;x=91490000;
#10;x=91500000;
#10;x=91510000;
#10;x=91520000;
#10;x=91530000;
#10;x=91540000;
#10;x=91550000;
#10;x=91560000;
#10;x=91570000;
#10;x=91580000;
#10;x=91590000;
#10;x=91600000;
#10;x=91610000;
#10;x=91620000;
#10;x=91630000;
#10;x=91640000;
#10;x=91650000;
#10;x=91660000;
#10;x=91670000;
#10;x=91680000;
#10;x=91690000;
#10;x=91700000;
#10;x=91710000;
#10;x=91720000;
#10;x=91730000;
#10;x=91740000;
#10;x=91750000;
#10;x=91760000;
#10;x=91770000;
#10;x=91780000;
#10;x=91790000;
#10;x=91800000;
#10;x=91810000;
#10;x=91820000;
#10;x=91830000;
#10;x=91840000;
#10;x=91850000;
#10;x=91860000;
#10;x=91870000;
#10;x=91880000;
#10;x=91890000;
#10;x=91900000;
#10;x=91910000;
#10;x=91920000;
#10;x=91930000;
#10;x=91940000;
#10;x=91950000;
#10;x=91960000;
#10;x=91970000;
#10;x=91980000;
#10;x=91990000;
#10;x=92000000;
#10;x=92010000;
#10;x=92020000;
#10;x=92030000;
#10;x=92040000;
#10;x=92050000;
#10;x=92060000;
#10;x=92070000;
#10;x=92080000;
#10;x=92090000;
#10;x=92100000;
#10;x=92110000;
#10;x=92120000;
#10;x=92130000;
#10;x=92140000;
#10;x=92150000;
#10;x=92160000;
#10;x=92170000;
#10;x=92180000;
#10;x=92190000;
#10;x=92200000;
#10;x=92210000;
#10;x=92220000;
#10;x=92230000;
#10;x=92240000;
#10;x=92250000;
#10;x=92260000;
#10;x=92270000;
#10;x=92280000;
#10;x=92290000;
#10;x=92300000;
#10;x=92310000;
#10;x=92320000;
#10;x=92330000;
#10;x=92340000;
#10;x=92350000;
#10;x=92360000;
#10;x=92370000;
#10;x=92380000;
#10;x=92390000;
#10;x=92400000;
#10;x=92410000;
#10;x=92420000;
#10;x=92430000;
#10;x=92440000;
#10;x=92450000;
#10;x=92460000;
#10;x=92470000;
#10;x=92480000;
#10;x=92490000;
#10;x=92500000;
#10;x=92510000;
#10;x=92520000;
#10;x=92530000;
#10;x=92540000;
#10;x=92550000;
#10;x=92560000;
#10;x=92570000;
#10;x=92580000;
#10;x=92590000;
#10;x=92600000;
#10;x=92610000;
#10;x=92620000;
#10;x=92630000;
#10;x=92640000;
#10;x=92650000;
#10;x=92660000;
#10;x=92670000;
#10;x=92680000;
#10;x=92690000;
#10;x=92700000;
#10;x=92710000;
#10;x=92720000;
#10;x=92730000;
#10;x=92740000;
#10;x=92750000;
#10;x=92760000;
#10;x=92770000;
#10;x=92780000;
#10;x=92790000;
#10;x=92800000;
#10;x=92810000;
#10;x=92820000;
#10;x=92830000;
#10;x=92840000;
#10;x=92850000;
#10;x=92860000;
#10;x=92870000;
#10;x=92880000;
#10;x=92890000;
#10;x=92900000;
#10;x=92910000;
#10;x=92920000;
#10;x=92930000;
#10;x=92940000;
#10;x=92950000;
#10;x=92960000;
#10;x=92970000;
#10;x=92980000;
#10;x=92990000;
#10;x=93000000;
#10;x=93010000;
#10;x=93020000;
#10;x=93030000;
#10;x=93040000;
#10;x=93050000;
#10;x=93060000;
#10;x=93070000;
#10;x=93080000;
#10;x=93090000;
#10;x=93100000;
#10;x=93110000;
#10;x=93120000;
#10;x=93130000;
#10;x=93140000;
#10;x=93150000;
#10;x=93160000;
#10;x=93170000;
#10;x=93180000;
#10;x=93190000;
#10;x=93200000;
#10;x=93210000;
#10;x=93220000;
#10;x=93230000;
#10;x=93240000;
#10;x=93250000;
#10;x=93260000;
#10;x=93270000;
#10;x=93280000;
#10;x=93290000;
#10;x=93300000;
#10;x=93310000;
#10;x=93320000;
#10;x=93330000;
#10;x=93340000;
#10;x=93350000;
#10;x=93360000;
#10;x=93370000;
#10;x=93380000;
#10;x=93390000;
#10;x=93400000;
#10;x=93410000;
#10;x=93420000;
#10;x=93430000;
#10;x=93440000;
#10;x=93450000;
#10;x=93460000;
#10;x=93470000;
#10;x=93480000;
#10;x=93490000;
#10;x=93500000;
#10;x=93510000;
#10;x=93520000;
#10;x=93530000;
#10;x=93540000;
#10;x=93550000;
#10;x=93560000;
#10;x=93570000;
#10;x=93580000;
#10;x=93590000;
#10;x=93600000;
#10;x=93610000;
#10;x=93620000;
#10;x=93630000;
#10;x=93640000;
#10;x=93650000;
#10;x=93660000;
#10;x=93670000;
#10;x=93680000;
#10;x=93690000;
#10;x=93700000;
#10;x=93710000;
#10;x=93720000;
#10;x=93730000;
#10;x=93740000;
#10;x=93750000;
#10;x=93760000;
#10;x=93770000;
#10;x=93780000;
#10;x=93790000;
#10;x=93800000;
#10;x=93810000;
#10;x=93820000;
#10;x=93830000;
#10;x=93840000;
#10;x=93850000;
#10;x=93860000;
#10;x=93870000;
#10;x=93880000;
#10;x=93890000;
#10;x=93900000;
#10;x=93910000;
#10;x=93920000;
#10;x=93930000;
#10;x=93940000;
#10;x=93950000;
#10;x=93960000;
#10;x=93970000;
#10;x=93980000;
#10;x=93990000;
#10;x=94000000;
#10;x=94010000;
#10;x=94020000;
#10;x=94030000;
#10;x=94040000;
#10;x=94050000;
#10;x=94060000;
#10;x=94070000;
#10;x=94080000;
#10;x=94090000;
#10;x=94100000;
#10;x=94110000;
#10;x=94120000;
#10;x=94130000;
#10;x=94140000;
#10;x=94150000;
#10;x=94160000;
#10;x=94170000;
#10;x=94180000;
#10;x=94190000;
#10;x=94200000;
#10;x=94210000;
#10;x=94220000;
#10;x=94230000;
#10;x=94240000;
#10;x=94250000;
#10;x=94260000;
#10;x=94270000;
#10;x=94280000;
#10;x=94290000;
#10;x=94300000;
#10;x=94310000;
#10;x=94320000;
#10;x=94330000;
#10;x=94340000;
#10;x=94350000;
#10;x=94360000;
#10;x=94370000;
#10;x=94380000;
#10;x=94390000;
#10;x=94400000;
#10;x=94410000;
#10;x=94420000;
#10;x=94430000;
#10;x=94440000;
#10;x=94450000;
#10;x=94460000;
#10;x=94470000;
#10;x=94480000;
#10;x=94490000;
#10;x=94500000;
#10;x=94510000;
#10;x=94520000;
#10;x=94530000;
#10;x=94540000;
#10;x=94550000;
#10;x=94560000;
#10;x=94570000;
#10;x=94580000;
#10;x=94590000;
#10;x=94600000;
#10;x=94610000;
#10;x=94620000;
#10;x=94630000;
#10;x=94640000;
#10;x=94650000;
#10;x=94660000;
#10;x=94670000;
#10;x=94680000;
#10;x=94690000;
#10;x=94700000;
#10;x=94710000;
#10;x=94720000;
#10;x=94730000;
#10;x=94740000;
#10;x=94750000;
#10;x=94760000;
#10;x=94770000;
#10;x=94780000;
#10;x=94790000;
#10;x=94800000;
#10;x=94810000;
#10;x=94820000;
#10;x=94830000;
#10;x=94840000;
#10;x=94850000;
#10;x=94860000;
#10;x=94870000;
#10;x=94880000;
#10;x=94890000;
#10;x=94900000;
#10;x=94910000;
#10;x=94920000;
#10;x=94930000;
#10;x=94940000;
#10;x=94950000;
#10;x=94960000;
#10;x=94970000;
#10;x=94980000;
#10;x=94990000;
#10;x=95000000;
#10;x=95010000;
#10;x=95020000;
#10;x=95030000;
#10;x=95040000;
#10;x=95050000;
#10;x=95060000;
#10;x=95070000;
#10;x=95080000;
#10;x=95090000;
#10;x=95100000;
#10;x=95110000;
#10;x=95120000;
#10;x=95130000;
#10;x=95140000;
#10;x=95150000;
#10;x=95160000;
#10;x=95170000;
#10;x=95180000;
#10;x=95190000;
#10;x=95200000;
#10;x=95210000;
#10;x=95220000;
#10;x=95230000;
#10;x=95240000;
#10;x=95250000;
#10;x=95260000;
#10;x=95270000;
#10;x=95280000;
#10;x=95290000;
#10;x=95300000;
#10;x=95310000;
#10;x=95320000;
#10;x=95330000;
#10;x=95340000;
#10;x=95350000;
#10;x=95360000;
#10;x=95370000;
#10;x=95380000;
#10;x=95390000;
#10;x=95400000;
#10;x=95410000;
#10;x=95420000;
#10;x=95430000;
#10;x=95440000;
#10;x=95450000;
#10;x=95460000;
#10;x=95470000;
#10;x=95480000;
#10;x=95490000;
#10;x=95500000;
#10;x=95510000;
#10;x=95520000;
#10;x=95530000;
#10;x=95540000;
#10;x=95550000;
#10;x=95560000;
#10;x=95570000;
#10;x=95580000;
#10;x=95590000;
#10;x=95600000;
#10;x=95610000;
#10;x=95620000;
#10;x=95630000;
#10;x=95640000;
#10;x=95650000;
#10;x=95660000;
#10;x=95670000;
#10;x=95680000;
#10;x=95690000;
#10;x=95700000;
#10;x=95710000;
#10;x=95720000;
#10;x=95730000;
#10;x=95740000;
#10;x=95750000;
#10;x=95760000;
#10;x=95770000;
#10;x=95780000;
#10;x=95790000;
#10;x=95800000;
#10;x=95810000;
#10;x=95820000;
#10;x=95830000;
#10;x=95840000;
#10;x=95850000;
#10;x=95860000;
#10;x=95870000;
#10;x=95880000;
#10;x=95890000;
#10;x=95900000;
#10;x=95910000;
#10;x=95920000;
#10;x=95930000;
#10;x=95940000;
#10;x=95950000;
#10;x=95960000;
#10;x=95970000;
#10;x=95980000;
#10;x=95990000;
#10;x=96000000;
#10;x=96010000;
#10;x=96020000;
#10;x=96030000;
#10;x=96040000;
#10;x=96050000;
#10;x=96060000;
#10;x=96070000;
#10;x=96080000;
#10;x=96090000;
#10;x=96100000;
#10;x=96110000;
#10;x=96120000;
#10;x=96130000;
#10;x=96140000;
#10;x=96150000;
#10;x=96160000;
#10;x=96170000;
#10;x=96180000;
#10;x=96190000;
#10;x=96200000;
#10;x=96210000;
#10;x=96220000;
#10;x=96230000;
#10;x=96240000;
#10;x=96250000;
#10;x=96260000;
#10;x=96270000;
#10;x=96280000;
#10;x=96290000;
#10;x=96300000;
#10;x=96310000;
#10;x=96320000;
#10;x=96330000;
#10;x=96340000;
#10;x=96350000;
#10;x=96360000;
#10;x=96370000;
#10;x=96380000;
#10;x=96390000;
#10;x=96400000;
#10;x=96410000;
#10;x=96420000;
#10;x=96430000;
#10;x=96440000;
#10;x=96450000;
#10;x=96460000;
#10;x=96470000;
#10;x=96480000;
#10;x=96490000;
#10;x=96500000;
#10;x=96510000;
#10;x=96520000;
#10;x=96530000;
#10;x=96540000;
#10;x=96550000;
#10;x=96560000;
#10;x=96570000;
#10;x=96580000;
#10;x=96590000;
#10;x=96600000;
#10;x=96610000;
#10;x=96620000;
#10;x=96630000;
#10;x=96640000;
#10;x=96650000;
#10;x=96660000;
#10;x=96670000;
#10;x=96680000;
#10;x=96690000;
#10;x=96700000;
#10;x=96710000;
#10;x=96720000;
#10;x=96730000;
#10;x=96740000;
#10;x=96750000;
#10;x=96760000;
#10;x=96770000;
#10;x=96780000;
#10;x=96790000;
#10;x=96800000;
#10;x=96810000;
#10;x=96820000;
#10;x=96830000;
#10;x=96840000;
#10;x=96850000;
#10;x=96860000;
#10;x=96870000;
#10;x=96880000;
#10;x=96890000;
#10;x=96900000;
#10;x=96910000;
#10;x=96920000;
#10;x=96930000;
#10;x=96940000;
#10;x=96950000;
#10;x=96960000;
#10;x=96970000;
#10;x=96980000;
#10;x=96990000;
#10;x=97000000;
#10;x=97010000;
#10;x=97020000;
#10;x=97030000;
#10;x=97040000;
#10;x=97050000;
#10;x=97060000;
#10;x=97070000;
#10;x=97080000;
#10;x=97090000;
#10;x=97100000;
#10;x=97110000;
#10;x=97120000;
#10;x=97130000;
#10;x=97140000;
#10;x=97150000;
#10;x=97160000;
#10;x=97170000;
#10;x=97180000;
#10;x=97190000;
#10;x=97200000;
#10;x=97210000;
#10;x=97220000;
#10;x=97230000;
#10;x=97240000;
#10;x=97250000;
#10;x=97260000;
#10;x=97270000;
#10;x=97280000;
#10;x=97290000;
#10;x=97300000;
#10;x=97310000;
#10;x=97320000;
#10;x=97330000;
#10;x=97340000;
#10;x=97350000;
#10;x=97360000;
#10;x=97370000;
#10;x=97380000;
#10;x=97390000;
#10;x=97400000;
#10;x=97410000;
#10;x=97420000;
#10;x=97430000;
#10;x=97440000;
#10;x=97450000;
#10;x=97460000;
#10;x=97470000;
#10;x=97480000;
#10;x=97490000;
#10;x=97500000;
#10;x=97510000;
#10;x=97520000;
#10;x=97530000;
#10;x=97540000;
#10;x=97550000;
#10;x=97560000;
#10;x=97570000;
#10;x=97580000;
#10;x=97590000;
#10;x=97600000;
#10;x=97610000;
#10;x=97620000;
#10;x=97630000;
#10;x=97640000;
#10;x=97650000;
#10;x=97660000;
#10;x=97670000;
#10;x=97680000;
#10;x=97690000;
#10;x=97700000;
#10;x=97710000;
#10;x=97720000;
#10;x=97730000;
#10;x=97740000;
#10;x=97750000;
#10;x=97760000;
#10;x=97770000;
#10;x=97780000;
#10;x=97790000;
#10;x=97800000;
#10;x=97810000;
#10;x=97820000;
#10;x=97830000;
#10;x=97840000;
#10;x=97850000;
#10;x=97860000;
#10;x=97870000;
#10;x=97880000;
#10;x=97890000;
#10;x=97900000;
#10;x=97910000;
#10;x=97920000;
#10;x=97930000;
#10;x=97940000;
#10;x=97950000;
#10;x=97960000;
#10;x=97970000;
#10;x=97980000;
#10;x=97990000;
#10;x=98000000;
#10;x=98010000;
#10;x=98020000;
#10;x=98030000;
#10;x=98040000;
#10;x=98050000;
#10;x=98060000;
#10;x=98070000;
#10;x=98080000;
#10;x=98090000;
#10;x=98100000;
#10;x=98110000;
#10;x=98120000;
#10;x=98130000;
#10;x=98140000;
#10;x=98150000;
#10;x=98160000;
#10;x=98170000;
#10;x=98180000;
#10;x=98190000;
#10;x=98200000;
#10;x=98210000;
#10;x=98220000;
#10;x=98230000;
#10;x=98240000;
#10;x=98250000;
#10;x=98260000;
#10;x=98270000;
#10;x=98280000;
#10;x=98290000;
#10;x=98300000;
#10;x=98310000;
#10;x=98320000;
#10;x=98330000;
#10;x=98340000;
#10;x=98350000;
#10;x=98360000;
#10;x=98370000;
#10;x=98380000;
#10;x=98390000;
#10;x=98400000;
#10;x=98410000;
#10;x=98420000;
#10;x=98430000;
#10;x=98440000;
#10;x=98450000;
#10;x=98460000;
#10;x=98470000;
#10;x=98480000;
#10;x=98490000;
#10;x=98500000;
#10;x=98510000;
#10;x=98520000;
#10;x=98530000;
#10;x=98540000;
#10;x=98550000;
#10;x=98560000;
#10;x=98570000;
#10;x=98580000;
#10;x=98590000;
#10;x=98600000;
#10;x=98610000;
#10;x=98620000;
#10;x=98630000;
#10;x=98640000;
#10;x=98650000;
#10;x=98660000;
#10;x=98670000;
#10;x=98680000;
#10;x=98690000;
#10;x=98700000;
#10;x=98710000;
#10;x=98720000;
#10;x=98730000;
#10;x=98740000;
#10;x=98750000;
#10;x=98760000;
#10;x=98770000;
#10;x=98780000;
#10;x=98790000;
#10;x=98800000;
#10;x=98810000;
#10;x=98820000;
#10;x=98830000;
#10;x=98840000;
#10;x=98850000;
#10;x=98860000;
#10;x=98870000;
#10;x=98880000;
#10;x=98890000;
#10;x=98900000;
#10;x=98910000;
#10;x=98920000;
#10;x=98930000;
#10;x=98940000;
#10;x=98950000;
#10;x=98960000;
#10;x=98970000;
#10;x=98980000;
#10;x=98990000;
#10;x=99000000;
#10;x=99010000;
#10;x=99020000;
#10;x=99030000;
#10;x=99040000;
#10;x=99050000;
#10;x=99060000;
#10;x=99070000;
#10;x=99080000;
#10;x=99090000;
#10;x=99100000;
#10;x=99110000;
#10;x=99120000;
#10;x=99130000;
#10;x=99140000;
#10;x=99150000;
#10;x=99160000;
#10;x=99170000;
#10;x=99180000;
#10;x=99190000;
#10;x=99200000;
#10;x=99210000;
#10;x=99220000;
#10;x=99230000;
#10;x=99240000;
#10;x=99250000;
#10;x=99260000;
#10;x=99270000;
#10;x=99280000;
#10;x=99290000;
#10;x=99300000;
#10;x=99310000;
#10;x=99320000;
#10;x=99330000;
#10;x=99340000;
#10;x=99350000;
#10;x=99360000;
#10;x=99370000;
#10;x=99380000;
#10;x=99390000;
#10;x=99400000;
#10;x=99410000;
#10;x=99420000;
#10;x=99430000;
#10;x=99440000;
#10;x=99450000;
#10;x=99460000;
#10;x=99470000;
#10;x=99480000;
#10;x=99490000;
#10;x=99500000;
#10;x=99510000;
#10;x=99520000;
#10;x=99530000;
#10;x=99540000;
#10;x=99550000;
#10;x=99560000;
#10;x=99570000;
#10;x=99580000;
#10;x=99590000;
#10;x=99600000;
#10;x=99610000;
#10;x=99620000;
#10;x=99630000;
#10;x=99640000;
#10;x=99650000;
#10;x=99660000;
#10;x=99670000;
#10;x=99680000;
#10;x=99690000;
#10;x=99700000;
#10;x=99710000;
#10;x=99720000;
#10;x=99730000;
#10;x=99740000;
#10;x=99750000;
#10;x=99760000;
#10;x=99770000;
#10;x=99780000;
#10;x=99790000;
#10;x=99800000;
#10;x=99810000;
#10;x=99820000;
#10;x=99830000;
#10;x=99840000;
#10;x=99850000;
#10;x=99860000;
#10;x=99870000;
#10;x=99880000;
#10;x=99890000;
#10;x=99900000;
#10;x=99910000;
#10;x=99920000;
#10;x=99930000;
#10;x=99940000;
#10;x=99950000;
#10;x=99960000;
#10;x=99970000;
#10;x=99980000;
#10;x=99990000;
#10;x=100000000;
#10;x=100010000;
#10;x=100020000;
#10;x=100030000;
#10;x=100040000;
#10;x=100050000;
#10;x=100060000;
#10;x=100070000;
#10;x=100080000;
#10;x=100090000;
#10;x=100100000;
#10;x=100110000;
#10;x=100120000;
#10;x=100130000;
#10;x=100140000;
#10;x=100150000;
#10;x=100160000;
#10;x=100170000;
#10;x=100180000;
#10;x=100190000;
#10;x=100200000;
#10;x=100210000;
#10;x=100220000;
#10;x=100230000;
#10;x=100240000;
#10;x=100250000;
#10;x=100260000;
#10;x=100270000;
#10;x=100280000;
#10;x=100290000;
#10;x=100300000;
#10;x=100310000;
#10;x=100320000;
#10;x=100330000;
#10;x=100340000;
#10;x=100350000;
#10;x=100360000;
#10;x=100370000;
#10;x=100380000;
#10;x=100390000;
#10;x=100400000;
#10;x=100410000;
#10;x=100420000;
#10;x=100430000;
#10;x=100440000;
#10;x=100450000;
#10;x=100460000;
#10;x=100470000;
#10;x=100480000;
#10;x=100490000;
#10;x=100500000;
#10;x=100510000;
#10;x=100520000;
#10;x=100530000;
#10;x=100540000;
#10;x=100550000;
#10;x=100560000;
#10;x=100570000;
#10;x=100580000;
#10;x=100590000;
#10;x=100600000;
#10;x=100610000;
#10;x=100620000;
#10;x=100630000;
#10;x=100640000;
#10;x=100650000;
#10;x=100660000;
#10;x=100670000;
#10;x=100680000;
#10;x=100690000;
#10;x=100700000;
#10;x=100710000;
#10;x=100720000;
#10;x=100730000;
#10;x=100740000;
#10;x=100750000;
#10;x=100760000;
#10;x=100770000;
#10;x=100780000;
#10;x=100790000;
#10;x=100800000;
#10;x=100810000;
#10;x=100820000;
#10;x=100830000;
#10;x=100840000;
#10;x=100850000;
#10;x=100860000;
#10;x=100870000;
#10;x=100880000;
#10;x=100890000;
#10;x=100900000;
#10;x=100910000;
#10;x=100920000;
#10;x=100930000;
#10;x=100940000;
#10;x=100950000;
#10;x=100960000;
#10;x=100970000;
#10;x=100980000;
#10;x=100990000;
#10;x=101000000;
#10;x=101010000;
#10;x=101020000;
#10;x=101030000;
#10;x=101040000;
#10;x=101050000;
#10;x=101060000;
#10;x=101070000;
#10;x=101080000;
#10;x=101090000;
#10;x=101100000;
#10;x=101110000;
#10;x=101120000;
#10;x=101130000;
#10;x=101140000;
#10;x=101150000;
#10;x=101160000;
#10;x=101170000;
#10;x=101180000;
#10;x=101190000;
#10;x=101200000;
#10;x=101210000;
#10;x=101220000;
#10;x=101230000;
#10;x=101240000;
#10;x=101250000;
#10;x=101260000;
#10;x=101270000;
#10;x=101280000;
#10;x=101290000;
#10;x=101300000;
#10;x=101310000;
#10;x=101320000;
#10;x=101330000;
#10;x=101340000;
#10;x=101350000;
#10;x=101360000;
#10;x=101370000;
#10;x=101380000;
#10;x=101390000;
#10;x=101400000;
#10;x=101410000;
#10;x=101420000;
#10;x=101430000;
#10;x=101440000;
#10;x=101450000;
#10;x=101460000;
#10;x=101470000;
#10;x=101480000;
#10;x=101490000;
#10;x=101500000;
#10;x=101510000;
#10;x=101520000;
#10;x=101530000;
#10;x=101540000;
#10;x=101550000;
#10;x=101560000;
#10;x=101570000;
#10;x=101580000;
#10;x=101590000;
#10;x=101600000;
#10;x=101610000;
#10;x=101620000;
#10;x=101630000;
#10;x=101640000;
#10;x=101650000;
#10;x=101660000;
#10;x=101670000;
#10;x=101680000;
#10;x=101690000;
#10;x=101700000;
#10;x=101710000;
#10;x=101720000;
#10;x=101730000;
#10;x=101740000;
#10;x=101750000;
#10;x=101760000;
#10;x=101770000;
#10;x=101780000;
#10;x=101790000;
#10;x=101800000;
#10;x=101810000;
#10;x=101820000;
#10;x=101830000;
#10;x=101840000;
#10;x=101850000;
#10;x=101860000;
#10;x=101870000;
#10;x=101880000;
#10;x=101890000;
#10;x=101900000;
#10;x=101910000;
#10;x=101920000;
#10;x=101930000;
#10;x=101940000;
#10;x=101950000;
#10;x=101960000;
#10;x=101970000;
#10;x=101980000;
#10;x=101990000;
#10;x=102000000;
#10;x=102010000;
#10;x=102020000;
#10;x=102030000;
#10;x=102040000;
#10;x=102050000;
#10;x=102060000;
#10;x=102070000;
#10;x=102080000;
#10;x=102090000;
#10;x=102100000;
#10;x=102110000;
#10;x=102120000;
#10;x=102130000;
#10;x=102140000;
#10;x=102150000;
#10;x=102160000;
#10;x=102170000;
#10;x=102180000;
#10;x=102190000;
#10;x=102200000;
#10;x=102210000;
#10;x=102220000;
#10;x=102230000;
#10;x=102240000;
#10;x=102250000;
#10;x=102260000;
#10;x=102270000;
#10;x=102280000;
#10;x=102290000;
#10;x=102300000;
#10;x=102310000;
#10;x=102320000;
#10;x=102330000;
#10;x=102340000;
#10;x=102350000;
#10;x=102360000;
#10;x=102370000;
#10;x=102380000;
#10;x=102390000;
#10;x=102400000;
#10;x=102410000;
#10;x=102420000;
#10;x=102430000;
#10;x=102440000;
#10;x=102450000;
#10;x=102460000;
#10;x=102470000;
#10;x=102480000;
#10;x=102490000;
#10;x=102500000;
#10;x=102510000;
#10;x=102520000;
#10;x=102530000;
#10;x=102540000;
#10;x=102550000;
#10;x=102560000;
#10;x=102570000;
#10;x=102580000;
#10;x=102590000;
#10;x=102600000;
#10;x=102610000;
#10;x=102620000;
#10;x=102630000;
#10;x=102640000;
#10;x=102650000;
#10;x=102660000;
#10;x=102670000;
#10;x=102680000;
#10;x=102690000;
#10;x=102700000;
#10;x=102710000;
#10;x=102720000;
#10;x=102730000;
#10;x=102740000;
#10;x=102750000;
#10;x=102760000;
#10;x=102770000;
#10;x=102780000;
#10;x=102790000;
#10;x=102800000;
#10;x=102810000;
#10;x=102820000;
#10;x=102830000;
#10;x=102840000;
#10;x=102850000;
#10;x=102860000;
#10;x=102870000;
#10;x=102880000;
#10;x=102890000;
#10;x=102900000;
#10;x=102910000;
#10;x=102920000;
#10;x=102930000;
#10;x=102940000;
#10;x=102950000;
#10;x=102960000;
#10;x=102970000;
#10;x=102980000;
#10;x=102990000;
#10;x=103000000;
#10;x=103010000;
#10;x=103020000;
#10;x=103030000;
#10;x=103040000;
#10;x=103050000;
#10;x=103060000;
#10;x=103070000;
#10;x=103080000;
#10;x=103090000;
#10;x=103100000;
#10;x=103110000;
#10;x=103120000;
#10;x=103130000;
#10;x=103140000;
#10;x=103150000;
#10;x=103160000;
#10;x=103170000;
#10;x=103180000;
#10;x=103190000;
#10;x=103200000;
#10;x=103210000;
#10;x=103220000;
#10;x=103230000;
#10;x=103240000;
#10;x=103250000;
#10;x=103260000;
#10;x=103270000;
#10;x=103280000;
#10;x=103290000;
#10;x=103300000;
#10;x=103310000;
#10;x=103320000;
#10;x=103330000;
#10;x=103340000;
#10;x=103350000;
#10;x=103360000;
#10;x=103370000;
#10;x=103380000;
#10;x=103390000;
#10;x=103400000;
#10;x=103410000;
#10;x=103420000;
#10;x=103430000;
#10;x=103440000;
#10;x=103450000;
#10;x=103460000;
#10;x=103470000;
#10;x=103480000;
#10;x=103490000;
#10;x=103500000;
#10;x=103510000;
#10;x=103520000;
#10;x=103530000;
#10;x=103540000;
#10;x=103550000;
#10;x=103560000;
#10;x=103570000;
#10;x=103580000;
#10;x=103590000;
#10;x=103600000;
#10;x=103610000;
#10;x=103620000;
#10;x=103630000;
#10;x=103640000;
#10;x=103650000;
#10;x=103660000;
#10;x=103670000;
#10;x=103680000;
#10;x=103690000;
#10;x=103700000;
#10;x=103710000;
#10;x=103720000;
#10;x=103730000;
#10;x=103740000;
#10;x=103750000;
#10;x=103760000;
#10;x=103770000;
#10;x=103780000;
#10;x=103790000;
#10;x=103800000;
#10;x=103810000;
#10;x=103820000;
#10;x=103830000;
#10;x=103840000;
#10;x=103850000;
#10;x=103860000;
#10;x=103870000;
#10;x=103880000;
#10;x=103890000;
#10;x=103900000;
#10;x=103910000;
#10;x=103920000;
#10;x=103930000;
#10;x=103940000;
#10;x=103950000;
#10;x=103960000;
#10;x=103970000;
#10;x=103980000;
#10;x=103990000;
#10;x=104000000;
#10;x=104010000;
#10;x=104020000;
#10;x=104030000;
#10;x=104040000;
#10;x=104050000;
#10;x=104060000;
#10;x=104070000;
#10;x=104080000;
#10;x=104090000;
#10;x=104100000;
#10;x=104110000;
#10;x=104120000;
#10;x=104130000;
#10;x=104140000;
#10;x=104150000;
#10;x=104160000;
#10;x=104170000;
#10;x=104180000;
#10;x=104190000;
#10;x=104200000;
#10;x=104210000;
#10;x=104220000;
#10;x=104230000;
#10;x=104240000;
#10;x=104250000;
#10;x=104260000;
#10;x=104270000;
#10;x=104280000;
#10;x=104290000;
#10;x=104300000;
#10;x=104310000;
#10;x=104320000;
#10;x=104330000;
#10;x=104340000;
#10;x=104350000;
#10;x=104360000;
#10;x=104370000;
#10;x=104380000;
#10;x=104390000;
#10;x=104400000;
#10;x=104410000;
#10;x=104420000;
#10;x=104430000;
#10;x=104440000;
#10;x=104450000;
#10;x=104460000;
#10;x=104470000;
#10;x=104480000;
#10;x=104490000;
#10;x=104500000;
#10;x=104510000;
#10;x=104520000;
#10;x=104530000;
#10;x=104540000;
#10;x=104550000;
#10;x=104560000;
#10;x=104570000;
#10;x=104580000;
#10;x=104590000;
#10;x=104600000;
#10;x=104610000;
#10;x=104620000;
#10;x=104630000;
#10;x=104640000;
#10;x=104650000;
#10;x=104660000;
#10;x=104670000;
#10;x=104680000;
#10;x=104690000;
#10;x=104700000;
#10;x=104710000;
#10;x=104720000;
#10;x=104730000;
#10;x=104740000;
#10;x=104750000;
#10;x=104760000;
#10;x=104770000;
#10;x=104780000;
#10;x=104790000;
#10;x=104800000;
#10;x=104810000;
#10;x=104820000;
#10;x=104830000;
#10;x=104840000;
#10;x=104850000;
#10;x=104860000;
#10;x=104870000;
#10;x=104880000;
#10;x=104890000;
#10;x=104900000;
#10;x=104910000;
#10;x=104920000;
#10;x=104930000;
#10;x=104940000;
#10;x=104950000;
#10;x=104960000;
#10;x=104970000;
#10;x=104980000;
#10;x=104990000;
#10;x=105000000;
#10;x=105010000;
#10;x=105020000;
#10;x=105030000;
#10;x=105040000;
#10;x=105050000;
#10;x=105060000;
#10;x=105070000;
#10;x=105080000;
#10;x=105090000;
#10;x=105100000;
#10;x=105110000;
#10;x=105120000;
#10;x=105130000;
#10;x=105140000;
#10;x=105150000;
#10;x=105160000;
#10;x=105170000;
#10;x=105180000;
#10;x=105190000;
#10;x=105200000;
#10;x=105210000;
#10;x=105220000;
#10;x=105230000;
#10;x=105240000;
#10;x=105250000;
#10;x=105260000;
#10;x=105270000;
#10;x=105280000;
#10;x=105290000;
#10;x=105300000;
#10;x=105310000;
#10;x=105320000;
#10;x=105330000;
#10;x=105340000;
#10;x=105350000;
#10;x=105360000;
#10;x=105370000;
#10;x=105380000;
#10;x=105390000;
#10;x=105400000;
#10;x=105410000;
#10;x=105420000;
#10;x=105430000;
#10;x=105440000;
#10;x=105450000;
#10;x=105460000;
#10;x=105470000;
#10;x=105480000;
#10;x=105490000;
#10;x=105500000;
#10;x=105510000;
#10;x=105520000;
#10;x=105530000;
#10;x=105540000;
#10;x=105550000;
#10;x=105560000;
#10;x=105570000;
#10;x=105580000;
#10;x=105590000;
#10;x=105600000;
#10;x=105610000;
#10;x=105620000;
#10;x=105630000;
#10;x=105640000;
#10;x=105650000;
#10;x=105660000;
#10;x=105670000;
#10;x=105680000;
#10;x=105690000;
#10;x=105700000;
#10;x=105710000;
#10;x=105720000;
#10;x=105730000;
#10;x=105740000;
#10;x=105750000;
#10;x=105760000;
#10;x=105770000;
#10;x=105780000;
#10;x=105790000;
#10;x=105800000;
#10;x=105810000;
#10;x=105820000;
#10;x=105830000;
#10;x=105840000;
#10;x=105850000;
#10;x=105860000;
#10;x=105870000;
#10;x=105880000;
#10;x=105890000;
#10;x=105900000;
#10;x=105910000;
#10;x=105920000;
#10;x=105930000;
#10;x=105940000;
#10;x=105950000;
#10;x=105960000;
#10;x=105970000;
#10;x=105980000;
#10;x=105990000;
#10;x=106000000;
#10;x=106010000;
#10;x=106020000;
#10;x=106030000;
#10;x=106040000;
#10;x=106050000;
#10;x=106060000;
#10;x=106070000;
#10;x=106080000;
#10;x=106090000;
#10;x=106100000;
#10;x=106110000;
#10;x=106120000;
#10;x=106130000;
#10;x=106140000;
#10;x=106150000;
#10;x=106160000;
#10;x=106170000;
#10;x=106180000;
#10;x=106190000;
#10;x=106200000;
#10;x=106210000;
#10;x=106220000;
#10;x=106230000;
#10;x=106240000;
#10;x=106250000;
#10;x=106260000;
#10;x=106270000;
#10;x=106280000;
#10;x=106290000;
#10;x=106300000;
#10;x=106310000;
#10;x=106320000;
#10;x=106330000;
#10;x=106340000;
#10;x=106350000;
#10;x=106360000;
#10;x=106370000;
#10;x=106380000;
#10;x=106390000;
#10;x=106400000;
#10;x=106410000;
#10;x=106420000;
#10;x=106430000;
#10;x=106440000;
#10;x=106450000;
#10;x=106460000;
#10;x=106470000;
#10;x=106480000;
#10;x=106490000;
#10;x=106500000;
#10;x=106510000;
#10;x=106520000;
#10;x=106530000;
#10;x=106540000;
#10;x=106550000;
#10;x=106560000;
#10;x=106570000;
#10;x=106580000;
#10;x=106590000;
#10;x=106600000;
#10;x=106610000;
#10;x=106620000;
#10;x=106630000;
#10;x=106640000;
#10;x=106650000;
#10;x=106660000;
#10;x=106670000;
#10;x=106680000;
#10;x=106690000;
#10;x=106700000;
#10;x=106710000;
#10;x=106720000;
#10;x=106730000;
#10;x=106740000;
#10;x=106750000;
#10;x=106760000;
#10;x=106770000;
#10;x=106780000;
#10;x=106790000;
#10;x=106800000;
#10;x=106810000;
#10;x=106820000;
#10;x=106830000;
#10;x=106840000;
#10;x=106850000;
#10;x=106860000;
#10;x=106870000;
#10;x=106880000;
#10;x=106890000;
#10;x=106900000;
#10;x=106910000;
#10;x=106920000;
#10;x=106930000;
#10;x=106940000;
#10;x=106950000;
#10;x=106960000;
#10;x=106970000;
#10;x=106980000;
#10;x=106990000;
#10;x=107000000;
#10;x=107010000;
#10;x=107020000;
#10;x=107030000;
#10;x=107040000;
#10;x=107050000;
#10;x=107060000;
#10;x=107070000;
#10;x=107080000;
#10;x=107090000;
#10;x=107100000;
#10;x=107110000;
#10;x=107120000;
#10;x=107130000;
#10;x=107140000;
#10;x=107150000;
#10;x=107160000;
#10;x=107170000;
#10;x=107180000;
#10;x=107190000;
#10;x=107200000;
#10;x=107210000;
#10;x=107220000;
#10;x=107230000;
#10;x=107240000;
#10;x=107250000;
#10;x=107260000;
#10;x=107270000;
#10;x=107280000;
#10;x=107290000;
#10;x=107300000;
#10;x=107310000;
#10;x=107320000;
#10;x=107330000;
#10;x=107340000;
#10;x=107350000;
#10;x=107360000;
#10;x=107370000;
#10;x=107380000;
#10;x=107390000;
#10;x=107400000;
#10;x=107410000;
#10;x=107420000;
#10;x=107430000;
#10;x=107440000;
#10;x=107450000;
#10;x=107460000;
#10;x=107470000;
#10;x=107480000;
#10;x=107490000;
#10;x=107500000;
#10;x=107510000;
#10;x=107520000;
#10;x=107530000;
#10;x=107540000;
#10;x=107550000;
#10;x=107560000;
#10;x=107570000;
#10;x=107580000;
#10;x=107590000;
#10;x=107600000;
#10;x=107610000;
#10;x=107620000;
#10;x=107630000;
#10;x=107640000;
#10;x=107650000;
#10;x=107660000;
#10;x=107670000;
#10;x=107680000;
#10;x=107690000;
#10;x=107700000;
#10;x=107710000;
#10;x=107720000;
#10;x=107730000;
#10;x=107740000;
#10;x=107750000;
#10;x=107760000;
#10;x=107770000;
#10;x=107780000;
#10;x=107790000;
#10;x=107800000;
#10;x=107810000;
#10;x=107820000;
#10;x=107830000;
#10;x=107840000;
#10;x=107850000;
#10;x=107860000;
#10;x=107870000;
#10;x=107880000;
#10;x=107890000;
#10;x=107900000;
#10;x=107910000;
#10;x=107920000;
#10;x=107930000;
#10;x=107940000;
#10;x=107950000;
#10;x=107960000;
#10;x=107970000;
#10;x=107980000;
#10;x=107990000;
#10;x=108000000;
#10;x=108010000;
#10;x=108020000;
#10;x=108030000;
#10;x=108040000;
#10;x=108050000;
#10;x=108060000;
#10;x=108070000;
#10;x=108080000;
#10;x=108090000;
#10;x=108100000;
#10;x=108110000;
#10;x=108120000;
#10;x=108130000;
#10;x=108140000;
#10;x=108150000;
#10;x=108160000;
#10;x=108170000;
#10;x=108180000;
#10;x=108190000;
#10;x=108200000;
#10;x=108210000;
#10;x=108220000;
#10;x=108230000;
#10;x=108240000;
#10;x=108250000;
#10;x=108260000;
#10;x=108270000;
#10;x=108280000;
#10;x=108290000;
#10;x=108300000;
#10;x=108310000;
#10;x=108320000;
#10;x=108330000;
#10;x=108340000;
#10;x=108350000;
#10;x=108360000;
#10;x=108370000;
#10;x=108380000;
#10;x=108390000;
#10;x=108400000;
#10;x=108410000;
#10;x=108420000;
#10;x=108430000;
#10;x=108440000;
#10;x=108450000;
#10;x=108460000;
#10;x=108470000;
#10;x=108480000;
#10;x=108490000;
#10;x=108500000;
#10;x=108510000;
#10;x=108520000;
#10;x=108530000;
#10;x=108540000;
#10;x=108550000;
#10;x=108560000;
#10;x=108570000;
#10;x=108580000;
#10;x=108590000;
#10;x=108600000;
#10;x=108610000;
#10;x=108620000;
#10;x=108630000;
#10;x=108640000;
#10;x=108650000;
#10;x=108660000;
#10;x=108670000;
#10;x=108680000;
#10;x=108690000;
#10;x=108700000;
#10;x=108710000;
#10;x=108720000;
#10;x=108730000;
#10;x=108740000;
#10;x=108750000;
#10;x=108760000;
#10;x=108770000;
#10;x=108780000;
#10;x=108790000;
#10;x=108800000;
#10;x=108810000;
#10;x=108820000;
#10;x=108830000;
#10;x=108840000;
#10;x=108850000;
#10;x=108860000;
#10;x=108870000;
#10;x=108880000;
#10;x=108890000;
#10;x=108900000;
#10;x=108910000;
#10;x=108920000;
#10;x=108930000;
#10;x=108940000;
#10;x=108950000;
#10;x=108960000;
#10;x=108970000;
#10;x=108980000;
#10;x=108990000;
#10;x=109000000;
#10;x=109010000;
#10;x=109020000;
#10;x=109030000;
#10;x=109040000;
#10;x=109050000;
#10;x=109060000;
#10;x=109070000;
#10;x=109080000;
#10;x=109090000;
#10;x=109100000;
#10;x=109110000;
#10;x=109120000;
#10;x=109130000;
#10;x=109140000;
#10;x=109150000;
#10;x=109160000;
#10;x=109170000;
#10;x=109180000;
#10;x=109190000;
#10;x=109200000;
#10;x=109210000;
#10;x=109220000;
#10;x=109230000;
#10;x=109240000;
#10;x=109250000;
#10;x=109260000;
#10;x=109270000;
#10;x=109280000;
#10;x=109290000;
#10;x=109300000;
#10;x=109310000;
#10;x=109320000;
#10;x=109330000;
#10;x=109340000;
#10;x=109350000;
#10;x=109360000;
#10;x=109370000;
#10;x=109380000;
#10;x=109390000;
#10;x=109400000;
#10;x=109410000;
#10;x=109420000;
#10;x=109430000;
#10;x=109440000;
#10;x=109450000;
#10;x=109460000;
#10;x=109470000;
#10;x=109480000;
#10;x=109490000;
#10;x=109500000;
#10;x=109510000;
#10;x=109520000;
#10;x=109530000;
#10;x=109540000;
#10;x=109550000;
#10;x=109560000;
#10;x=109570000;
#10;x=109580000;
#10;x=109590000;
#10;x=109600000;
#10;x=109610000;
#10;x=109620000;
#10;x=109630000;
#10;x=109640000;
#10;x=109650000;
#10;x=109660000;
#10;x=109670000;
#10;x=109680000;
#10;x=109690000;
#10;x=109700000;
#10;x=109710000;
#10;x=109720000;
#10;x=109730000;
#10;x=109740000;
#10;x=109750000;
#10;x=109760000;
#10;x=109770000;
#10;x=109780000;
#10;x=109790000;
#10;x=109800000;
#10;x=109810000;
#10;x=109820000;
#10;x=109830000;
#10;x=109840000;
#10;x=109850000;
#10;x=109860000;
#10;x=109870000;
#10;x=109880000;
#10;x=109890000;
#10;x=109900000;
#10;x=109910000;
#10;x=109920000;
#10;x=109930000;
#10;x=109940000;
#10;x=109950000;
#10;x=109960000;
#10;x=109970000;
#10;x=109980000;
#10;x=109990000;
#10;x=110000000;
#10;x=110010000;
#10;x=110020000;
#10;x=110030000;
#10;x=110040000;
#10;x=110050000;
#10;x=110060000;
#10;x=110070000;
#10;x=110080000;
#10;x=110090000;
#10;x=110100000;
#10;x=110110000;
#10;x=110120000;
#10;x=110130000;
#10;x=110140000;
#10;x=110150000;
#10;x=110160000;
#10;x=110170000;
#10;x=110180000;
#10;x=110190000;
#10;x=110200000;
#10;x=110210000;
#10;x=110220000;
#10;x=110230000;
#10;x=110240000;
#10;x=110250000;
#10;x=110260000;
#10;x=110270000;
#10;x=110280000;
#10;x=110290000;
#10;x=110300000;
#10;x=110310000;
#10;x=110320000;
#10;x=110330000;
#10;x=110340000;
#10;x=110350000;
#10;x=110360000;
#10;x=110370000;
#10;x=110380000;
#10;x=110390000;
#10;x=110400000;
#10;x=110410000;
#10;x=110420000;
#10;x=110430000;
#10;x=110440000;
#10;x=110450000;
#10;x=110460000;
#10;x=110470000;
#10;x=110480000;
#10;x=110490000;
#10;x=110500000;
#10;x=110510000;
#10;x=110520000;
#10;x=110530000;
#10;x=110540000;
#10;x=110550000;
#10;x=110560000;
#10;x=110570000;
#10;x=110580000;
#10;x=110590000;
#10;x=110600000;
#10;x=110610000;
#10;x=110620000;
#10;x=110630000;
#10;x=110640000;
#10;x=110650000;
#10;x=110660000;
#10;x=110670000;
#10;x=110680000;
#10;x=110690000;
#10;x=110700000;
#10;x=110710000;
#10;x=110720000;
#10;x=110730000;
#10;x=110740000;
#10;x=110750000;
#10;x=110760000;
#10;x=110770000;
#10;x=110780000;
#10;x=110790000;
#10;x=110800000;
#10;x=110810000;
#10;x=110820000;
#10;x=110830000;
#10;x=110840000;
#10;x=110850000;
#10;x=110860000;
#10;x=110870000;
#10;x=110880000;
#10;x=110890000;
#10;x=110900000;
#10;x=110910000;
#10;x=110920000;
#10;x=110930000;
#10;x=110940000;
#10;x=110950000;
#10;x=110960000;
#10;x=110970000;
#10;x=110980000;
#10;x=110990000;
#10;x=111000000;
#10;x=111010000;
#10;x=111020000;
#10;x=111030000;
#10;x=111040000;
#10;x=111050000;
#10;x=111060000;
#10;x=111070000;
#10;x=111080000;
#10;x=111090000;
#10;x=111100000;
#10;x=111110000;
#10;x=111120000;
#10;x=111130000;
#10;x=111140000;
#10;x=111150000;
#10;x=111160000;
#10;x=111170000;
#10;x=111180000;
#10;x=111190000;
#10;x=111200000;
#10;x=111210000;
#10;x=111220000;
#10;x=111230000;
#10;x=111240000;
#10;x=111250000;
#10;x=111260000;
#10;x=111270000;
#10;x=111280000;
#10;x=111290000;
#10;x=111300000;
#10;x=111310000;
#10;x=111320000;
#10;x=111330000;
#10;x=111340000;
#10;x=111350000;
#10;x=111360000;
#10;x=111370000;
#10;x=111380000;
#10;x=111390000;
#10;x=111400000;
#10;x=111410000;
#10;x=111420000;
#10;x=111430000;
#10;x=111440000;
#10;x=111450000;
#10;x=111460000;
#10;x=111470000;
#10;x=111480000;
#10;x=111490000;
#10;x=111500000;
#10;x=111510000;
#10;x=111520000;
#10;x=111530000;
#10;x=111540000;
#10;x=111550000;
#10;x=111560000;
#10;x=111570000;
#10;x=111580000;
#10;x=111590000;
#10;x=111600000;
#10;x=111610000;
#10;x=111620000;
#10;x=111630000;
#10;x=111640000;
#10;x=111650000;
#10;x=111660000;
#10;x=111670000;
#10;x=111680000;
#10;x=111690000;
#10;x=111700000;
#10;x=111710000;
#10;x=111720000;
#10;x=111730000;
#10;x=111740000;
#10;x=111750000;
#10;x=111760000;
#10;x=111770000;
#10;x=111780000;
#10;x=111790000;
#10;x=111800000;
#10;x=111810000;
#10;x=111820000;
#10;x=111830000;
#10;x=111840000;
#10;x=111850000;
#10;x=111860000;
#10;x=111870000;
#10;x=111880000;
#10;x=111890000;
#10;x=111900000;
#10;x=111910000;
#10;x=111920000;
#10;x=111930000;
#10;x=111940000;
#10;x=111950000;
#10;x=111960000;
#10;x=111970000;
#10;x=111980000;
#10;x=111990000;
#10;x=112000000;
#10;x=112010000;
#10;x=112020000;
#10;x=112030000;
#10;x=112040000;
#10;x=112050000;
#10;x=112060000;
#10;x=112070000;
#10;x=112080000;
#10;x=112090000;
#10;x=112100000;
#10;x=112110000;
#10;x=112120000;
#10;x=112130000;
#10;x=112140000;
#10;x=112150000;
#10;x=112160000;
#10;x=112170000;
#10;x=112180000;
#10;x=112190000;
#10;x=112200000;
#10;x=112210000;
#10;x=112220000;
#10;x=112230000;
#10;x=112240000;
#10;x=112250000;
#10;x=112260000;
#10;x=112270000;
#10;x=112280000;
#10;x=112290000;
#10;x=112300000;
#10;x=112310000;
#10;x=112320000;
#10;x=112330000;
#10;x=112340000;
#10;x=112350000;
#10;x=112360000;
#10;x=112370000;
#10;x=112380000;
#10;x=112390000;
#10;x=112400000;
#10;x=112410000;
#10;x=112420000;
#10;x=112430000;
#10;x=112440000;
#10;x=112450000;
#10;x=112460000;
#10;x=112470000;
#10;x=112480000;
#10;x=112490000;
#10;x=112500000;
#10;x=112510000;
#10;x=112520000;
#10;x=112530000;
#10;x=112540000;
#10;x=112550000;
#10;x=112560000;
#10;x=112570000;
#10;x=112580000;
#10;x=112590000;
#10;x=112600000;
#10;x=112610000;
#10;x=112620000;
#10;x=112630000;
#10;x=112640000;
#10;x=112650000;
#10;x=112660000;
#10;x=112670000;
#10;x=112680000;
#10;x=112690000;
#10;x=112700000;
#10;x=112710000;
#10;x=112720000;
#10;x=112730000;
#10;x=112740000;
#10;x=112750000;
#10;x=112760000;
#10;x=112770000;
#10;x=112780000;
#10;x=112790000;
#10;x=112800000;
#10;x=112810000;
#10;x=112820000;
#10;x=112830000;
#10;x=112840000;
#10;x=112850000;
#10;x=112860000;
#10;x=112870000;
#10;x=112880000;
#10;x=112890000;
#10;x=112900000;
#10;x=112910000;
#10;x=112920000;
#10;x=112930000;
#10;x=112940000;
#10;x=112950000;
#10;x=112960000;
#10;x=112970000;
#10;x=112980000;
#10;x=112990000;
#10;x=113000000;
#10;x=113010000;
#10;x=113020000;
#10;x=113030000;
#10;x=113040000;
#10;x=113050000;
#10;x=113060000;
#10;x=113070000;
#10;x=113080000;
#10;x=113090000;
#10;x=113100000;
#10;x=113110000;
#10;x=113120000;
#10;x=113130000;
#10;x=113140000;
#10;x=113150000;
#10;x=113160000;
#10;x=113170000;
#10;x=113180000;
#10;x=113190000;
#10;x=113200000;
#10;x=113210000;
#10;x=113220000;
#10;x=113230000;
#10;x=113240000;
#10;x=113250000;
#10;x=113260000;
#10;x=113270000;
#10;x=113280000;
#10;x=113290000;
#10;x=113300000;
#10;x=113310000;
#10;x=113320000;
#10;x=113330000;
#10;x=113340000;
#10;x=113350000;
#10;x=113360000;
#10;x=113370000;
#10;x=113380000;
#10;x=113390000;
#10;x=113400000;
#10;x=113410000;
#10;x=113420000;
#10;x=113430000;
#10;x=113440000;
#10;x=113450000;
#10;x=113460000;
#10;x=113470000;
#10;x=113480000;
#10;x=113490000;
#10;x=113500000;
#10;x=113510000;
#10;x=113520000;
#10;x=113530000;
#10;x=113540000;
#10;x=113550000;
#10;x=113560000;
#10;x=113570000;
#10;x=113580000;
#10;x=113590000;
#10;x=113600000;
#10;x=113610000;
#10;x=113620000;
#10;x=113630000;
#10;x=113640000;
#10;x=113650000;
#10;x=113660000;
#10;x=113670000;
#10;x=113680000;
#10;x=113690000;
#10;x=113700000;
#10;x=113710000;
#10;x=113720000;
#10;x=113730000;
#10;x=113740000;
#10;x=113750000;
#10;x=113760000;
#10;x=113770000;
#10;x=113780000;
#10;x=113790000;
#10;x=113800000;
#10;x=113810000;
#10;x=113820000;
#10;x=113830000;
#10;x=113840000;
#10;x=113850000;
#10;x=113860000;
#10;x=113870000;
#10;x=113880000;
#10;x=113890000;
#10;x=113900000;
#10;x=113910000;
#10;x=113920000;
#10;x=113930000;
#10;x=113940000;
#10;x=113950000;
#10;x=113960000;
#10;x=113970000;
#10;x=113980000;
#10;x=113990000;
#10;x=114000000;
#10;x=114010000;
#10;x=114020000;
#10;x=114030000;
#10;x=114040000;
#10;x=114050000;
#10;x=114060000;
#10;x=114070000;
#10;x=114080000;
#10;x=114090000;
#10;x=114100000;
#10;x=114110000;
#10;x=114120000;
#10;x=114130000;
#10;x=114140000;
#10;x=114150000;
#10;x=114160000;
#10;x=114170000;
#10;x=114180000;
#10;x=114190000;
#10;x=114200000;
#10;x=114210000;
#10;x=114220000;
#10;x=114230000;
#10;x=114240000;
#10;x=114250000;
#10;x=114260000;
#10;x=114270000;
#10;x=114280000;
#10;x=114290000;
#10;x=114300000;
#10;x=114310000;
#10;x=114320000;
#10;x=114330000;
#10;x=114340000;
#10;x=114350000;
#10;x=114360000;
#10;x=114370000;
#10;x=114380000;
#10;x=114390000;
#10;x=114400000;
#10;x=114410000;
#10;x=114420000;
#10;x=114430000;
#10;x=114440000;
#10;x=114450000;
#10;x=114460000;
#10;x=114470000;
#10;x=114480000;
#10;x=114490000;
#10;x=114500000;
#10;x=114510000;
#10;x=114520000;
#10;x=114530000;
#10;x=114540000;
#10;x=114550000;
#10;x=114560000;
#10;x=114570000;
#10;x=114580000;
#10;x=114590000;
#10;x=114600000;
#10;x=114610000;
#10;x=114620000;
#10;x=114630000;
#10;x=114640000;
#10;x=114650000;
#10;x=114660000;
#10;x=114670000;
#10;x=114680000;
#10;x=114690000;
#10;x=114700000;
#10;x=114710000;
#10;x=114720000;
#10;x=114730000;
#10;x=114740000;
#10;x=114750000;
#10;x=114760000;
#10;x=114770000;
#10;x=114780000;
#10;x=114790000;
#10;x=114800000;
#10;x=114810000;
#10;x=114820000;
#10;x=114830000;
#10;x=114840000;
#10;x=114850000;
#10;x=114860000;
#10;x=114870000;
#10;x=114880000;
#10;x=114890000;
#10;x=114900000;
#10;x=114910000;
#10;x=114920000;
#10;x=114930000;
#10;x=114940000;
#10;x=114950000;
#10;x=114960000;
#10;x=114970000;
#10;x=114980000;
#10;x=114990000;
#10;x=115000000;
#10;x=115010000;
#10;x=115020000;
#10;x=115030000;
#10;x=115040000;
#10;x=115050000;
#10;x=115060000;
#10;x=115070000;
#10;x=115080000;
#10;x=115090000;
#10;x=115100000;
#10;x=115110000;
#10;x=115120000;
#10;x=115130000;
#10;x=115140000;
#10;x=115150000;
#10;x=115160000;
#10;x=115170000;
#10;x=115180000;
#10;x=115190000;
#10;x=115200000;
#10;x=115210000;
#10;x=115220000;
#10;x=115230000;
#10;x=115240000;
#10;x=115250000;
#10;x=115260000;
#10;x=115270000;
#10;x=115280000;
#10;x=115290000;
#10;x=115300000;
#10;x=115310000;
#10;x=115320000;
#10;x=115330000;
#10;x=115340000;
#10;x=115350000;
#10;x=115360000;
#10;x=115370000;
#10;x=115380000;
#10;x=115390000;
#10;x=115400000;
#10;x=115410000;
#10;x=115420000;
#10;x=115430000;
#10;x=115440000;
#10;x=115450000;
#10;x=115460000;
#10;x=115470000;
#10;x=115480000;
#10;x=115490000;
#10;x=115500000;
#10;x=115510000;
#10;x=115520000;
#10;x=115530000;
#10;x=115540000;
#10;x=115550000;
#10;x=115560000;
#10;x=115570000;
#10;x=115580000;
#10;x=115590000;
#10;x=115600000;
#10;x=115610000;
#10;x=115620000;
#10;x=115630000;
#10;x=115640000;
#10;x=115650000;
#10;x=115660000;
#10;x=115670000;
#10;x=115680000;
#10;x=115690000;
#10;x=115700000;
#10;x=115710000;
#10;x=115720000;
#10;x=115730000;
#10;x=115740000;
#10;x=115750000;
#10;x=115760000;
#10;x=115770000;
#10;x=115780000;
#10;x=115790000;
#10;x=115800000;
#10;x=115810000;
#10;x=115820000;
#10;x=115830000;
#10;x=115840000;
#10;x=115850000;
#10;x=115860000;
#10;x=115870000;
#10;x=115880000;
#10;x=115890000;
#10;x=115900000;
#10;x=115910000;
#10;x=115920000;
#10;x=115930000;
#10;x=115940000;
#10;x=115950000;
#10;x=115960000;
#10;x=115970000;
#10;x=115980000;
#10;x=115990000;
#10;x=116000000;
#10;x=116010000;
#10;x=116020000;
#10;x=116030000;
#10;x=116040000;
#10;x=116050000;
#10;x=116060000;
#10;x=116070000;
#10;x=116080000;
#10;x=116090000;
#10;x=116100000;
#10;x=116110000;
#10;x=116120000;
#10;x=116130000;
#10;x=116140000;
#10;x=116150000;
#10;x=116160000;
#10;x=116170000;
#10;x=116180000;
#10;x=116190000;
#10;x=116200000;
#10;x=116210000;
#10;x=116220000;
#10;x=116230000;
#10;x=116240000;
#10;x=116250000;
#10;x=116260000;
#10;x=116270000;
#10;x=116280000;
#10;x=116290000;
#10;x=116300000;
#10;x=116310000;
#10;x=116320000;
#10;x=116330000;
#10;x=116340000;
#10;x=116350000;
#10;x=116360000;
#10;x=116370000;
#10;x=116380000;
#10;x=116390000;
#10;x=116400000;
#10;x=116410000;
#10;x=116420000;
#10;x=116430000;
#10;x=116440000;
#10;x=116450000;
#10;x=116460000;
#10;x=116470000;
#10;x=116480000;
#10;x=116490000;
#10;x=116500000;
#10;x=116510000;
#10;x=116520000;
#10;x=116530000;
#10;x=116540000;
#10;x=116550000;
#10;x=116560000;
#10;x=116570000;
#10;x=116580000;
#10;x=116590000;
#10;x=116600000;
#10;x=116610000;
#10;x=116620000;
#10;x=116630000;
#10;x=116640000;
#10;x=116650000;
#10;x=116660000;
#10;x=116670000;
#10;x=116680000;
#10;x=116690000;
#10;x=116700000;
#10;x=116710000;
#10;x=116720000;
#10;x=116730000;
#10;x=116740000;
#10;x=116750000;
#10;x=116760000;
#10;x=116770000;
#10;x=116780000;
#10;x=116790000;
#10;x=116800000;
#10;x=116810000;
#10;x=116820000;
#10;x=116830000;
#10;x=116840000;
#10;x=116850000;
#10;x=116860000;
#10;x=116870000;
#10;x=116880000;
#10;x=116890000;
#10;x=116900000;
#10;x=116910000;
#10;x=116920000;
#10;x=116930000;
#10;x=116940000;
#10;x=116950000;
#10;x=116960000;
#10;x=116970000;
#10;x=116980000;
#10;x=116990000;
#10;x=117000000;
#10;x=117010000;
#10;x=117020000;
#10;x=117030000;
#10;x=117040000;
#10;x=117050000;
#10;x=117060000;
#10;x=117070000;
#10;x=117080000;
#10;x=117090000;
#10;x=117100000;
#10;x=117110000;
#10;x=117120000;
#10;x=117130000;
#10;x=117140000;
#10;x=117150000;
#10;x=117160000;
#10;x=117170000;
#10;x=117180000;
#10;x=117190000;
#10;x=117200000;
#10;x=117210000;
#10;x=117220000;
#10;x=117230000;
#10;x=117240000;
#10;x=117250000;
#10;x=117260000;
#10;x=117270000;
#10;x=117280000;
#10;x=117290000;
#10;x=117300000;
#10;x=117310000;
#10;x=117320000;
#10;x=117330000;
#10;x=117340000;
#10;x=117350000;
#10;x=117360000;
#10;x=117370000;
#10;x=117380000;
#10;x=117390000;
#10;x=117400000;
#10;x=117410000;
#10;x=117420000;
#10;x=117430000;
#10;x=117440000;
#10;x=117450000;
#10;x=117460000;
#10;x=117470000;
#10;x=117480000;
#10;x=117490000;
#10;x=117500000;
#10;x=117510000;
#10;x=117520000;
#10;x=117530000;
#10;x=117540000;
#10;x=117550000;
#10;x=117560000;
#10;x=117570000;
#10;x=117580000;
#10;x=117590000;
#10;x=117600000;
#10;x=117610000;
#10;x=117620000;
#10;x=117630000;
#10;x=117640000;
#10;x=117650000;
#10;x=117660000;
#10;x=117670000;
#10;x=117680000;
#10;x=117690000;
#10;x=117700000;
#10;x=117710000;
#10;x=117720000;
#10;x=117730000;
#10;x=117740000;
#10;x=117750000;
#10;x=117760000;
#10;x=117770000;
#10;x=117780000;
#10;x=117790000;
#10;x=117800000;
#10;x=117810000;
#10;x=117820000;
#10;x=117830000;
#10;x=117840000;
#10;x=117850000;
#10;x=117860000;
#10;x=117870000;
#10;x=117880000;
#10;x=117890000;
#10;x=117900000;
#10;x=117910000;
#10;x=117920000;
#10;x=117930000;
#10;x=117940000;
#10;x=117950000;
#10;x=117960000;
#10;x=117970000;
#10;x=117980000;
#10;x=117990000;
#10;x=118000000;
#10;x=118010000;
#10;x=118020000;
#10;x=118030000;
#10;x=118040000;
#10;x=118050000;
#10;x=118060000;
#10;x=118070000;
#10;x=118080000;
#10;x=118090000;
#10;x=118100000;
#10;x=118110000;
#10;x=118120000;
#10;x=118130000;
#10;x=118140000;
#10;x=118150000;
#10;x=118160000;
#10;x=118170000;
#10;x=118180000;
#10;x=118190000;
#10;x=118200000;
#10;x=118210000;
#10;x=118220000;
#10;x=118230000;
#10;x=118240000;
#10;x=118250000;
#10;x=118260000;
#10;x=118270000;
#10;x=118280000;
#10;x=118290000;
#10;x=118300000;
#10;x=118310000;
#10;x=118320000;
#10;x=118330000;
#10;x=118340000;
#10;x=118350000;
#10;x=118360000;
#10;x=118370000;
#10;x=118380000;
#10;x=118390000;
#10;x=118400000;
#10;x=118410000;
#10;x=118420000;
#10;x=118430000;
#10;x=118440000;
#10;x=118450000;
#10;x=118460000;
#10;x=118470000;
#10;x=118480000;
#10;x=118490000;
#10;x=118500000;
#10;x=118510000;
#10;x=118520000;
#10;x=118530000;
#10;x=118540000;
#10;x=118550000;
#10;x=118560000;
#10;x=118570000;
#10;x=118580000;
#10;x=118590000;
#10;x=118600000;
#10;x=118610000;
#10;x=118620000;
#10;x=118630000;
#10;x=118640000;
#10;x=118650000;
#10;x=118660000;
#10;x=118670000;
#10;x=118680000;
#10;x=118690000;
#10;x=118700000;
#10;x=118710000;
#10;x=118720000;
#10;x=118730000;
#10;x=118740000;
#10;x=118750000;
#10;x=118760000;
#10;x=118770000;
#10;x=118780000;
#10;x=118790000;
#10;x=118800000;
#10;x=118810000;
#10;x=118820000;
#10;x=118830000;
#10;x=118840000;
#10;x=118850000;
#10;x=118860000;
#10;x=118870000;
#10;x=118880000;
#10;x=118890000;
#10;x=118900000;
#10;x=118910000;
#10;x=118920000;
#10;x=118930000;
#10;x=118940000;
#10;x=118950000;
#10;x=118960000;
#10;x=118970000;
#10;x=118980000;
#10;x=118990000;
#10;x=119000000;
#10;x=119010000;
#10;x=119020000;
#10;x=119030000;
#10;x=119040000;
#10;x=119050000;
#10;x=119060000;
#10;x=119070000;
#10;x=119080000;
#10;x=119090000;
#10;x=119100000;
#10;x=119110000;
#10;x=119120000;
#10;x=119130000;
#10;x=119140000;
#10;x=119150000;
#10;x=119160000;
#10;x=119170000;
#10;x=119180000;
#10;x=119190000;
#10;x=119200000;
#10;x=119210000;
#10;x=119220000;
#10;x=119230000;
#10;x=119240000;
#10;x=119250000;
#10;x=119260000;
#10;x=119270000;
#10;x=119280000;
#10;x=119290000;
#10;x=119300000;
#10;x=119310000;
#10;x=119320000;
#10;x=119330000;
#10;x=119340000;
#10;x=119350000;
#10;x=119360000;
#10;x=119370000;
#10;x=119380000;
#10;x=119390000;
#10;x=119400000;
#10;x=119410000;
#10;x=119420000;
#10;x=119430000;
#10;x=119440000;
#10;x=119450000;
#10;x=119460000;
#10;x=119470000;
#10;x=119480000;
#10;x=119490000;
#10;x=119500000;
#10;x=119510000;
#10;x=119520000;
#10;x=119530000;
#10;x=119540000;
#10;x=119550000;
#10;x=119560000;
#10;x=119570000;
#10;x=119580000;
#10;x=119590000;
#10;x=119600000;
#10;x=119610000;
#10;x=119620000;
#10;x=119630000;
#10;x=119640000;
#10;x=119650000;
#10;x=119660000;
#10;x=119670000;
#10;x=119680000;
#10;x=119690000;
#10;x=119700000;
#10;x=119710000;
#10;x=119720000;
#10;x=119730000;
#10;x=119740000;
#10;x=119750000;
#10;x=119760000;
#10;x=119770000;
#10;x=119780000;
#10;x=119790000;
#10;x=119800000;
#10;x=119810000;
#10;x=119820000;
#10;x=119830000;
#10;x=119840000;
#10;x=119850000;
#10;x=119860000;
#10;x=119870000;
#10;x=119880000;
#10;x=119890000;
#10;x=119900000;
#10;x=119910000;
#10;x=119920000;
#10;x=119930000;
#10;x=119940000;
#10;x=119950000;
#10;x=119960000;
#10;x=119970000;
#10;x=119980000;
#10;x=119990000;
#10;x=120000000;
#10;x=120010000;
#10;x=120020000;
#10;x=120030000;
#10;x=120040000;
#10;x=120050000;
#10;x=120060000;
#10;x=120070000;
#10;x=120080000;
#10;x=120090000;
#10;x=120100000;
#10;x=120110000;
#10;x=120120000;
#10;x=120130000;
#10;x=120140000;
#10;x=120150000;
#10;x=120160000;
#10;x=120170000;
#10;x=120180000;
#10;x=120190000;
#10;x=120200000;
#10;x=120210000;
#10;x=120220000;
#10;x=120230000;
#10;x=120240000;
#10;x=120250000;
#10;x=120260000;
#10;x=120270000;
#10;x=120280000;
#10;x=120290000;
#10;x=120300000;
#10;x=120310000;
#10;x=120320000;
#10;x=120330000;
#10;x=120340000;
#10;x=120350000;
#10;x=120360000;
#10;x=120370000;
#10;x=120380000;
#10;x=120390000;
#10;x=120400000;
#10;x=120410000;
#10;x=120420000;
#10;x=120430000;
#10;x=120440000;
#10;x=120450000;
#10;x=120460000;
#10;x=120470000;
#10;x=120480000;
#10;x=120490000;
#10;x=120500000;
#10;x=120510000;
#10;x=120520000;
#10;x=120530000;
#10;x=120540000;
#10;x=120550000;
#10;x=120560000;
#10;x=120570000;
#10;x=120580000;
#10;x=120590000;
#10;x=120600000;
#10;x=120610000;
#10;x=120620000;
#10;x=120630000;
#10;x=120640000;
#10;x=120650000;
#10;x=120660000;
#10;x=120670000;
#10;x=120680000;
#10;x=120690000;
#10;x=120700000;
#10;x=120710000;
#10;x=120720000;
#10;x=120730000;
#10;x=120740000;
#10;x=120750000;
#10;x=120760000;
#10;x=120770000;
#10;x=120780000;
#10;x=120790000;
#10;x=120800000;
#10;x=120810000;
#10;x=120820000;
#10;x=120830000;
#10;x=120840000;
#10;x=120850000;
#10;x=120860000;
#10;x=120870000;
#10;x=120880000;
#10;x=120890000;
#10;x=120900000;
#10;x=120910000;
#10;x=120920000;
#10;x=120930000;
#10;x=120940000;
#10;x=120950000;
#10;x=120960000;
#10;x=120970000;
#10;x=120980000;
#10;x=120990000;
#10;x=121000000;
#10;x=121010000;
#10;x=121020000;
#10;x=121030000;
#10;x=121040000;
#10;x=121050000;
#10;x=121060000;
#10;x=121070000;
#10;x=121080000;
#10;x=121090000;
#10;x=121100000;
#10;x=121110000;
#10;x=121120000;
#10;x=121130000;
#10;x=121140000;
#10;x=121150000;
#10;x=121160000;
#10;x=121170000;
#10;x=121180000;
#10;x=121190000;
#10;x=121200000;
#10;x=121210000;
#10;x=121220000;
#10;x=121230000;
#10;x=121240000;
#10;x=121250000;
#10;x=121260000;
#10;x=121270000;
#10;x=121280000;
#10;x=121290000;
#10;x=121300000;
#10;x=121310000;
#10;x=121320000;
#10;x=121330000;
#10;x=121340000;
#10;x=121350000;
#10;x=121360000;
#10;x=121370000;
#10;x=121380000;
#10;x=121390000;
#10;x=121400000;
#10;x=121410000;
#10;x=121420000;
#10;x=121430000;
#10;x=121440000;
#10;x=121450000;
#10;x=121460000;
#10;x=121470000;
#10;x=121480000;
#10;x=121490000;
#10;x=121500000;
#10;x=121510000;
#10;x=121520000;
#10;x=121530000;
#10;x=121540000;
#10;x=121550000;
#10;x=121560000;
#10;x=121570000;
#10;x=121580000;
#10;x=121590000;
#10;x=121600000;
#10;x=121610000;
#10;x=121620000;
#10;x=121630000;
#10;x=121640000;
#10;x=121650000;
#10;x=121660000;
#10;x=121670000;
#10;x=121680000;
#10;x=121690000;
#10;x=121700000;
#10;x=121710000;
#10;x=121720000;
#10;x=121730000;
#10;x=121740000;
#10;x=121750000;
#10;x=121760000;
#10;x=121770000;
#10;x=121780000;
#10;x=121790000;
#10;x=121800000;
#10;x=121810000;
#10;x=121820000;
#10;x=121830000;
#10;x=121840000;
#10;x=121850000;
#10;x=121860000;
#10;x=121870000;
#10;x=121880000;
#10;x=121890000;
#10;x=121900000;
#10;x=121910000;
#10;x=121920000;
#10;x=121930000;
#10;x=121940000;
#10;x=121950000;
#10;x=121960000;
#10;x=121970000;
#10;x=121980000;
#10;x=121990000;
#10;x=122000000;
#10;x=122010000;
#10;x=122020000;
#10;x=122030000;
#10;x=122040000;
#10;x=122050000;
#10;x=122060000;
#10;x=122070000;
#10;x=122080000;
#10;x=122090000;
#10;x=122100000;
#10;x=122110000;
#10;x=122120000;
#10;x=122130000;
#10;x=122140000;
#10;x=122150000;
#10;x=122160000;
#10;x=122170000;
#10;x=122180000;
#10;x=122190000;
#10;x=122200000;
#10;x=122210000;
#10;x=122220000;
#10;x=122230000;
#10;x=122240000;
#10;x=122250000;
#10;x=122260000;
#10;x=122270000;
#10;x=122280000;
#10;x=122290000;
#10;x=122300000;
#10;x=122310000;
#10;x=122320000;
#10;x=122330000;
#10;x=122340000;
#10;x=122350000;
#10;x=122360000;
#10;x=122370000;
#10;x=122380000;
#10;x=122390000;
#10;x=122400000;
#10;x=122410000;
#10;x=122420000;
#10;x=122430000;
#10;x=122440000;
#10;x=122450000;
#10;x=122460000;
#10;x=122470000;
#10;x=122480000;
#10;x=122490000;
#10;x=122500000;
#10;x=122510000;
#10;x=122520000;
#10;x=122530000;
#10;x=122540000;
#10;x=122550000;
#10;x=122560000;
#10;x=122570000;
#10;x=122580000;
#10;x=122590000;
#10;x=122600000;
#10;x=122610000;
#10;x=122620000;
#10;x=122630000;
#10;x=122640000;
#10;x=122650000;
#10;x=122660000;
#10;x=122670000;
#10;x=122680000;
#10;x=122690000;
#10;x=122700000;
#10;x=122710000;
#10;x=122720000;
#10;x=122730000;
#10;x=122740000;
#10;x=122750000;
#10;x=122760000;
#10;x=122770000;
#10;x=122780000;
#10;x=122790000;
#10;x=122800000;
#10;x=122810000;
#10;x=122820000;
#10;x=122830000;
#10;x=122840000;
#10;x=122850000;
#10;x=122860000;
#10;x=122870000;
#10;x=122880000;
#10;x=122890000;
#10;x=122900000;
#10;x=122910000;
#10;x=122920000;
#10;x=122930000;
#10;x=122940000;
#10;x=122950000;
#10;x=122960000;
#10;x=122970000;
#10;x=122980000;
#10;x=122990000;
#10;x=123000000;
#10;x=123010000;
#10;x=123020000;
#10;x=123030000;
#10;x=123040000;
#10;x=123050000;
#10;x=123060000;
#10;x=123070000;
#10;x=123080000;
#10;x=123090000;
#10;x=123100000;
#10;x=123110000;
#10;x=123120000;
#10;x=123130000;
#10;x=123140000;
#10;x=123150000;
#10;x=123160000;
#10;x=123170000;
#10;x=123180000;
#10;x=123190000;
#10;x=123200000;
#10;x=123210000;
#10;x=123220000;
#10;x=123230000;
#10;x=123240000;
#10;x=123250000;
#10;x=123260000;
#10;x=123270000;
#10;x=123280000;
#10;x=123290000;
#10;x=123300000;
#10;x=123310000;
#10;x=123320000;
#10;x=123330000;
#10;x=123340000;
#10;x=123350000;
#10;x=123360000;
#10;x=123370000;
#10;x=123380000;
#10;x=123390000;
#10;x=123400000;
#10;x=123410000;
#10;x=123420000;
#10;x=123430000;
#10;x=123440000;
#10;x=123450000;
#10;x=123460000;
#10;x=123470000;
#10;x=123480000;
#10;x=123490000;
#10;x=123500000;
#10;x=123510000;
#10;x=123520000;
#10;x=123530000;
#10;x=123540000;
#10;x=123550000;
#10;x=123560000;
#10;x=123570000;
#10;x=123580000;
#10;x=123590000;
#10;x=123600000;
#10;x=123610000;
#10;x=123620000;
#10;x=123630000;
#10;x=123640000;
#10;x=123650000;
#10;x=123660000;
#10;x=123670000;
#10;x=123680000;
#10;x=123690000;
#10;x=123700000;
#10;x=123710000;
#10;x=123720000;
#10;x=123730000;
#10;x=123740000;
#10;x=123750000;
#10;x=123760000;
#10;x=123770000;
#10;x=123780000;
#10;x=123790000;
#10;x=123800000;
#10;x=123810000;
#10;x=123820000;
#10;x=123830000;
#10;x=123840000;
#10;x=123850000;
#10;x=123860000;
#10;x=123870000;
#10;x=123880000;
#10;x=123890000;
#10;x=123900000;
#10;x=123910000;
#10;x=123920000;
#10;x=123930000;
#10;x=123940000;
#10;x=123950000;
#10;x=123960000;
#10;x=123970000;
#10;x=123980000;
#10;x=123990000;
#10;x=124000000;
#10;x=124010000;
#10;x=124020000;
#10;x=124030000;
#10;x=124040000;
#10;x=124050000;
#10;x=124060000;
#10;x=124070000;
#10;x=124080000;
#10;x=124090000;
#10;x=124100000;
#10;x=124110000;
#10;x=124120000;
#10;x=124130000;
#10;x=124140000;
#10;x=124150000;
#10;x=124160000;
#10;x=124170000;
#10;x=124180000;
#10;x=124190000;
#10;x=124200000;
#10;x=124210000;
#10;x=124220000;
#10;x=124230000;
#10;x=124240000;
#10;x=124250000;
#10;x=124260000;
#10;x=124270000;
#10;x=124280000;
#10;x=124290000;
#10;x=124300000;
#10;x=124310000;
#10;x=124320000;
#10;x=124330000;
#10;x=124340000;
#10;x=124350000;
#10;x=124360000;
#10;x=124370000;
#10;x=124380000;
#10;x=124390000;
#10;x=124400000;
#10;x=124410000;
#10;x=124420000;
#10;x=124430000;
#10;x=124440000;
#10;x=124450000;
#10;x=124460000;
#10;x=124470000;
#10;x=124480000;
#10;x=124490000;
#10;x=124500000;
#10;x=124510000;
#10;x=124520000;
#10;x=124530000;
#10;x=124540000;
#10;x=124550000;
#10;x=124560000;
#10;x=124570000;
#10;x=124580000;
#10;x=124590000;
#10;x=124600000;
#10;x=124610000;
#10;x=124620000;
#10;x=124630000;
#10;x=124640000;
#10;x=124650000;
#10;x=124660000;
#10;x=124670000;
#10;x=124680000;
#10;x=124690000;
#10;x=124700000;
#10;x=124710000;
#10;x=124720000;
#10;x=124730000;
#10;x=124740000;
#10;x=124750000;
#10;x=124760000;
#10;x=124770000;
#10;x=124780000;
#10;x=124790000;
#10;x=124800000;
#10;x=124810000;
#10;x=124820000;
#10;x=124830000;
#10;x=124840000;
#10;x=124850000;
#10;x=124860000;
#10;x=124870000;
#10;x=124880000;
#10;x=124890000;
#10;x=124900000;
#10;x=124910000;
#10;x=124920000;
#10;x=124930000;
#10;x=124940000;
#10;x=124950000;
#10;x=124960000;
#10;x=124970000;
#10;x=124980000;
#10;x=124990000;
#10;x=125000000;
#10;x=125010000;
#10;x=125020000;
#10;x=125030000;
#10;x=125040000;
#10;x=125050000;
#10;x=125060000;
#10;x=125070000;
#10;x=125080000;
#10;x=125090000;
#10;x=125100000;
#10;x=125110000;
#10;x=125120000;
#10;x=125130000;
#10;x=125140000;
#10;x=125150000;
#10;x=125160000;
#10;x=125170000;
#10;x=125180000;
#10;x=125190000;
#10;x=125200000;
#10;x=125210000;
#10;x=125220000;
#10;x=125230000;
#10;x=125240000;
#10;x=125250000;
#10;x=125260000;
#10;x=125270000;
#10;x=125280000;
#10;x=125290000;
#10;x=125300000;
#10;x=125310000;
#10;x=125320000;
#10;x=125330000;
#10;x=125340000;
#10;x=125350000;
#10;x=125360000;
#10;x=125370000;
#10;x=125380000;
#10;x=125390000;
#10;x=125400000;
#10;x=125410000;
#10;x=125420000;
#10;x=125430000;
#10;x=125440000;
#10;x=125450000;
#10;x=125460000;
#10;x=125470000;
#10;x=125480000;
#10;x=125490000;
#10;x=125500000;
#10;x=125510000;
#10;x=125520000;
#10;x=125530000;
#10;x=125540000;
#10;x=125550000;
#10;x=125560000;
#10;x=125570000;
#10;x=125580000;
#10;x=125590000;
#10;x=125600000;
#10;x=125610000;
#10;x=125620000;
#10;x=125630000;
#10;x=125640000;
#10;x=125650000;
#10;x=125660000;
#10;x=125670000;
#10;x=125680000;
#10;x=125690000;
#10;x=125700000;
#10;x=125710000;
#10;x=125720000;
#10;x=125730000;
#10;x=125740000;
#10;x=125750000;
#10;x=125760000;
#10;x=125770000;
#10;x=125780000;
#10;x=125790000;
#10;x=125800000;
#10;x=125810000;
#10;x=125820000;
#10;x=125830000;
#10;x=125840000;
#10;x=125850000;
#10;x=125860000;
#10;x=125870000;
#10;x=125880000;
#10;x=125890000;
#10;x=125900000;
#10;x=125910000;
#10;x=125920000;
#10;x=125930000;
#10;x=125940000;
#10;x=125950000;
#10;x=125960000;
#10;x=125970000;
#10;x=125980000;
#10;x=125990000;
#10;x=126000000;
#10;x=126010000;
#10;x=126020000;
#10;x=126030000;
#10;x=126040000;
#10;x=126050000;
#10;x=126060000;
#10;x=126070000;
#10;x=126080000;
#10;x=126090000;
#10;x=126100000;
#10;x=126110000;
#10;x=126120000;
#10;x=126130000;
#10;x=126140000;
#10;x=126150000;
#10;x=126160000;
#10;x=126170000;
#10;x=126180000;
#10;x=126190000;
#10;x=126200000;
#10;x=126210000;
#10;x=126220000;
#10;x=126230000;
#10;x=126240000;
#10;x=126250000;
#10;x=126260000;
#10;x=126270000;
#10;x=126280000;
#10;x=126290000;
#10;x=126300000;
#10;x=126310000;
#10;x=126320000;
#10;x=126330000;
#10;x=126340000;
#10;x=126350000;
#10;x=126360000;
#10;x=126370000;
#10;x=126380000;
#10;x=126390000;
#10;x=126400000;
#10;x=126410000;
#10;x=126420000;
#10;x=126430000;
#10;x=126440000;
#10;x=126450000;
#10;x=126460000;
#10;x=126470000;
#10;x=126480000;
#10;x=126490000;
#10;x=126500000;
#10;x=126510000;
#10;x=126520000;
#10;x=126530000;
#10;x=126540000;
#10;x=126550000;
#10;x=126560000;
#10;x=126570000;
#10;x=126580000;
#10;x=126590000;
#10;x=126600000;
#10;x=126610000;
#10;x=126620000;
#10;x=126630000;
#10;x=126640000;
#10;x=126650000;
#10;x=126660000;
#10;x=126670000;
#10;x=126680000;
#10;x=126690000;
#10;x=126700000;
#10;x=126710000;
#10;x=126720000;
#10;x=126730000;
#10;x=126740000;
#10;x=126750000;
#10;x=126760000;
#10;x=126770000;
#10;x=126780000;
#10;x=126790000;
#10;x=126800000;
#10;x=126810000;
#10;x=126820000;
#10;x=126830000;
#10;x=126840000;
#10;x=126850000;
#10;x=126860000;
#10;x=126870000;
#10;x=126880000;
#10;x=126890000;
#10;x=126900000;
#10;x=126910000;
#10;x=126920000;
#10;x=126930000;
#10;x=126940000;
#10;x=126950000;
#10;x=126960000;
#10;x=126970000;
#10;x=126980000;
#10;x=126990000;
#10;x=127000000;
#10;x=127010000;
#10;x=127020000;
#10;x=127030000;
#10;x=127040000;
#10;x=127050000;
#10;x=127060000;
#10;x=127070000;
#10;x=127080000;
#10;x=127090000;
#10;x=127100000;
#10;x=127110000;
#10;x=127120000;
#10;x=127130000;
#10;x=127140000;
#10;x=127150000;
#10;x=127160000;
#10;x=127170000;
#10;x=127180000;
#10;x=127190000;
#10;x=127200000;
#10;x=127210000;
#10;x=127220000;
#10;x=127230000;
#10;x=127240000;
#10;x=127250000;
#10;x=127260000;
#10;x=127270000;
#10;x=127280000;
#10;x=127290000;
#10;x=127300000;
#10;x=127310000;
#10;x=127320000;
#10;x=127330000;
#10;x=127340000;
#10;x=127350000;
#10;x=127360000;
#10;x=127370000;
#10;x=127380000;
#10;x=127390000;
#10;x=127400000;
#10;x=127410000;
#10;x=127420000;
#10;x=127430000;
#10;x=127440000;
#10;x=127450000;
#10;x=127460000;
#10;x=127470000;
#10;x=127480000;
#10;x=127490000;
#10;x=127500000;
#10;x=127510000;
#10;x=127520000;
#10;x=127530000;
#10;x=127540000;
#10;x=127550000;
#10;x=127560000;
#10;x=127570000;
#10;x=127580000;
#10;x=127590000;
#10;x=127600000;
#10;x=127610000;
#10;x=127620000;
#10;x=127630000;
#10;x=127640000;
#10;x=127650000;
#10;x=127660000;
#10;x=127670000;
#10;x=127680000;
#10;x=127690000;
#10;x=127700000;
#10;x=127710000;
#10;x=127720000;
#10;x=127730000;
#10;x=127740000;
#10;x=127750000;
#10;x=127760000;
#10;x=127770000;
#10;x=127780000;
#10;x=127790000;
#10;x=127800000;
#10;x=127810000;
#10;x=127820000;
#10;x=127830000;
#10;x=127840000;
#10;x=127850000;
#10;x=127860000;
#10;x=127870000;
#10;x=127880000;
#10;x=127890000;
#10;x=127900000;
#10;x=127910000;
#10;x=127920000;
#10;x=127930000;
#10;x=127940000;
#10;x=127950000;
#10;x=127960000;
#10;x=127970000;
#10;x=127980000;
#10;x=127990000;
#10;x=128000000;
#10;x=128010000;
#10;x=128020000;
#10;x=128030000;
#10;x=128040000;
#10;x=128050000;
#10;x=128060000;
#10;x=128070000;
#10;x=128080000;
#10;x=128090000;
#10;x=128100000;
#10;x=128110000;
#10;x=128120000;
#10;x=128130000;
#10;x=128140000;
#10;x=128150000;
#10;x=128160000;
#10;x=128170000;
#10;x=128180000;
#10;x=128190000;
#10;x=128200000;
#10;x=128210000;
#10;x=128220000;
#10;x=128230000;
#10;x=128240000;
#10;x=128250000;
#10;x=128260000;
#10;x=128270000;
#10;x=128280000;
#10;x=128290000;
#10;x=128300000;
#10;x=128310000;
#10;x=128320000;
#10;x=128330000;
#10;x=128340000;
#10;x=128350000;
#10;x=128360000;
#10;x=128370000;
#10;x=128380000;
#10;x=128390000;
#10;x=128400000;
#10;x=128410000;
#10;x=128420000;
#10;x=128430000;
#10;x=128440000;
#10;x=128450000;
#10;x=128460000;
#10;x=128470000;
#10;x=128480000;
#10;x=128490000;
#10;x=128500000;
#10;x=128510000;
#10;x=128520000;
#10;x=128530000;
#10;x=128540000;
#10;x=128550000;
#10;x=128560000;
#10;x=128570000;
#10;x=128580000;
#10;x=128590000;
#10;x=128600000;
#10;x=128610000;
#10;x=128620000;
#10;x=128630000;
#10;x=128640000;
#10;x=128650000;
#10;x=128660000;
#10;x=128670000;
#10;x=128680000;
#10;x=128690000;
#10;x=128700000;
#10;x=128710000;
#10;x=128720000;
#10;x=128730000;
#10;x=128740000;
#10;x=128750000;
#10;x=128760000;
#10;x=128770000;
#10;x=128780000;
#10;x=128790000;
#10;x=128800000;
#10;x=128810000;
#10;x=128820000;
#10;x=128830000;
#10;x=128840000;
#10;x=128850000;
#10;x=128860000;
#10;x=128870000;
#10;x=128880000;
#10;x=128890000;
#10;x=128900000;
#10;x=128910000;
#10;x=128920000;
#10;x=128930000;
#10;x=128940000;
#10;x=128950000;
#10;x=128960000;
#10;x=128970000;
#10;x=128980000;
#10;x=128990000;
#10;x=129000000;
#10;x=129010000;
#10;x=129020000;
#10;x=129030000;
#10;x=129040000;
#10;x=129050000;
#10;x=129060000;
#10;x=129070000;
#10;x=129080000;
#10;x=129090000;
#10;x=129100000;
#10;x=129110000;
#10;x=129120000;
#10;x=129130000;
#10;x=129140000;
#10;x=129150000;
#10;x=129160000;
#10;x=129170000;
#10;x=129180000;
#10;x=129190000;
#10;x=129200000;
#10;x=129210000;
#10;x=129220000;
#10;x=129230000;
#10;x=129240000;
#10;x=129250000;
#10;x=129260000;
#10;x=129270000;
#10;x=129280000;
#10;x=129290000;
#10;x=129300000;
#10;x=129310000;
#10;x=129320000;
#10;x=129330000;
#10;x=129340000;
#10;x=129350000;
#10;x=129360000;
#10;x=129370000;
#10;x=129380000;
#10;x=129390000;
#10;x=129400000;
#10;x=129410000;
#10;x=129420000;
#10;x=129430000;
#10;x=129440000;
#10;x=129450000;
#10;x=129460000;
#10;x=129470000;
#10;x=129480000;
#10;x=129490000;
#10;x=129500000;
#10;x=129510000;
#10;x=129520000;
#10;x=129530000;
#10;x=129540000;
#10;x=129550000;
#10;x=129560000;
#10;x=129570000;
#10;x=129580000;
#10;x=129590000;
#10;x=129600000;
#10;x=129610000;
#10;x=129620000;
#10;x=129630000;
#10;x=129640000;
#10;x=129650000;
#10;x=129660000;
#10;x=129670000;
#10;x=129680000;
#10;x=129690000;
#10;x=129700000;
#10;x=129710000;
#10;x=129720000;
#10;x=129730000;
#10;x=129740000;
#10;x=129750000;
#10;x=129760000;
#10;x=129770000;
#10;x=129780000;
#10;x=129790000;
#10;x=129800000;
#10;x=129810000;
#10;x=129820000;
#10;x=129830000;
#10;x=129840000;
#10;x=129850000;
#10;x=129860000;
#10;x=129870000;
#10;x=129880000;
#10;x=129890000;
#10;x=129900000;
#10;x=129910000;
#10;x=129920000;
#10;x=129930000;
#10;x=129940000;
#10;x=129950000;
#10;x=129960000;
#10;x=129970000;
#10;x=129980000;
#10;x=129990000;
#10;x=130000000;
#10;x=130010000;
#10;x=130020000;
#10;x=130030000;
#10;x=130040000;
#10;x=130050000;
#10;x=130060000;
#10;x=130070000;
#10;x=130080000;
#10;x=130090000;
#10;x=130100000;
#10;x=130110000;
#10;x=130120000;
#10;x=130130000;
#10;x=130140000;
#10;x=130150000;
#10;x=130160000;
#10;x=130170000;
#10;x=130180000;
#10;x=130190000;
#10;x=130200000;
#10;x=130210000;
#10;x=130220000;
#10;x=130230000;
#10;x=130240000;
#10;x=130250000;
#10;x=130260000;
#10;x=130270000;
#10;x=130280000;
#10;x=130290000;
#10;x=130300000;
#10;x=130310000;
#10;x=130320000;
#10;x=130330000;
#10;x=130340000;
#10;x=130350000;
#10;x=130360000;
#10;x=130370000;
#10;x=130380000;
#10;x=130390000;
#10;x=130400000;
#10;x=130410000;
#10;x=130420000;
#10;x=130430000;
#10;x=130440000;
#10;x=130450000;
#10;x=130460000;
#10;x=130470000;
#10;x=130480000;
#10;x=130490000;
#10;x=130500000;
#10;x=130510000;
#10;x=130520000;
#10;x=130530000;
#10;x=130540000;
#10;x=130550000;
#10;x=130560000;
#10;x=130570000;
#10;x=130580000;
#10;x=130590000;
#10;x=130600000;
#10;x=130610000;
#10;x=130620000;
#10;x=130630000;
#10;x=130640000;
#10;x=130650000;
#10;x=130660000;
#10;x=130670000;
#10;x=130680000;
#10;x=130690000;
#10;x=130700000;
#10;x=130710000;
#10;x=130720000;
#10;x=130730000;
#10;x=130740000;
#10;x=130750000;
#10;x=130760000;
#10;x=130770000;
#10;x=130780000;
#10;x=130790000;
#10;x=130800000;
#10;x=130810000;
#10;x=130820000;
#10;x=130830000;
#10;x=130840000;
#10;x=130850000;
#10;x=130860000;
#10;x=130870000;
#10;x=130880000;
#10;x=130890000;
#10;x=130900000;
#10;x=130910000;
#10;x=130920000;
#10;x=130930000;
#10;x=130940000;
#10;x=130950000;
#10;x=130960000;
#10;x=130970000;
#10;x=130980000;
#10;x=130990000;
#10;x=131000000;
#10;x=131010000;
#10;x=131020000;
#10;x=131030000;
#10;x=131040000;
#10;x=131050000;
#10;x=131060000;
#10;x=131070000;
#10;x=131080000;
#10;x=131090000;
#10;x=131100000;
#10;x=131110000;
#10;x=131120000;
#10;x=131130000;
#10;x=131140000;
#10;x=131150000;
#10;x=131160000;
#10;x=131170000;
#10;x=131180000;
#10;x=131190000;
#10;x=131200000;
#10;x=131210000;
#10;x=131220000;
#10;x=131230000;
#10;x=131240000;
#10;x=131250000;
#10;x=131260000;
#10;x=131270000;
#10;x=131280000;
#10;x=131290000;
#10;x=131300000;
#10;x=131310000;
#10;x=131320000;
#10;x=131330000;
#10;x=131340000;
#10;x=131350000;
#10;x=131360000;
#10;x=131370000;
#10;x=131380000;
#10;x=131390000;
#10;x=131400000;
#10;x=131410000;
#10;x=131420000;
#10;x=131430000;
#10;x=131440000;
#10;x=131450000;
#10;x=131460000;
#10;x=131470000;
#10;x=131480000;
#10;x=131490000;
#10;x=131500000;
#10;x=131510000;
#10;x=131520000;
#10;x=131530000;
#10;x=131540000;
#10;x=131550000;
#10;x=131560000;
#10;x=131570000;
#10;x=131580000;
#10;x=131590000;
#10;x=131600000;
#10;x=131610000;
#10;x=131620000;
#10;x=131630000;
#10;x=131640000;
#10;x=131650000;
#10;x=131660000;
#10;x=131670000;
#10;x=131680000;
#10;x=131690000;
#10;x=131700000;
#10;x=131710000;
#10;x=131720000;
#10;x=131730000;
#10;x=131740000;
#10;x=131750000;
#10;x=131760000;
#10;x=131770000;
#10;x=131780000;
#10;x=131790000;
#10;x=131800000;
#10;x=131810000;
#10;x=131820000;
#10;x=131830000;
#10;x=131840000;
#10;x=131850000;
#10;x=131860000;
#10;x=131870000;
#10;x=131880000;
#10;x=131890000;
#10;x=131900000;
#10;x=131910000;
#10;x=131920000;
#10;x=131930000;
#10;x=131940000;
#10;x=131950000;
#10;x=131960000;
#10;x=131970000;
#10;x=131980000;
#10;x=131990000;
#10;x=132000000;
#10;x=132010000;
#10;x=132020000;
#10;x=132030000;
#10;x=132040000;
#10;x=132050000;
#10;x=132060000;
#10;x=132070000;
#10;x=132080000;
#10;x=132090000;
#10;x=132100000;
#10;x=132110000;
#10;x=132120000;
#10;x=132130000;
#10;x=132140000;
#10;x=132150000;
#10;x=132160000;
#10;x=132170000;
#10;x=132180000;
#10;x=132190000;
#10;x=132200000;
#10;x=132210000;
#10;x=132220000;
#10;x=132230000;
#10;x=132240000;
#10;x=132250000;
#10;x=132260000;
#10;x=132270000;
#10;x=132280000;
#10;x=132290000;
#10;x=132300000;
#10;x=132310000;
#10;x=132320000;
#10;x=132330000;
#10;x=132340000;
#10;x=132350000;
#10;x=132360000;
#10;x=132370000;
#10;x=132380000;
#10;x=132390000;
#10;x=132400000;
#10;x=132410000;
#10;x=132420000;
#10;x=132430000;
#10;x=132440000;
#10;x=132450000;
#10;x=132460000;
#10;x=132470000;
#10;x=132480000;
#10;x=132490000;
#10;x=132500000;
#10;x=132510000;
#10;x=132520000;
#10;x=132530000;
#10;x=132540000;
#10;x=132550000;
#10;x=132560000;
#10;x=132570000;
#10;x=132580000;
#10;x=132590000;
#10;x=132600000;
#10;x=132610000;
#10;x=132620000;
#10;x=132630000;
#10;x=132640000;
#10;x=132650000;
#10;x=132660000;
#10;x=132670000;
#10;x=132680000;
#10;x=132690000;
#10;x=132700000;
#10;x=132710000;
#10;x=132720000;
#10;x=132730000;
#10;x=132740000;
#10;x=132750000;
#10;x=132760000;
#10;x=132770000;
#10;x=132780000;
#10;x=132790000;
#10;x=132800000;
#10;x=132810000;
#10;x=132820000;
#10;x=132830000;
#10;x=132840000;
#10;x=132850000;
#10;x=132860000;
#10;x=132870000;
#10;x=132880000;
#10;x=132890000;
#10;x=132900000;
#10;x=132910000;
#10;x=132920000;
#10;x=132930000;
#10;x=132940000;
#10;x=132950000;
#10;x=132960000;
#10;x=132970000;
#10;x=132980000;
#10;x=132990000;
#10;x=133000000;
#10;x=133010000;
#10;x=133020000;
#10;x=133030000;
#10;x=133040000;
#10;x=133050000;
#10;x=133060000;
#10;x=133070000;
#10;x=133080000;
#10;x=133090000;
#10;x=133100000;
#10;x=133110000;
#10;x=133120000;
#10;x=133130000;
#10;x=133140000;
#10;x=133150000;
#10;x=133160000;
#10;x=133170000;
#10;x=133180000;
#10;x=133190000;
#10;x=133200000;
#10;x=133210000;
#10;x=133220000;
#10;x=133230000;
#10;x=133240000;
#10;x=133250000;
#10;x=133260000;
#10;x=133270000;
#10;x=133280000;
#10;x=133290000;
#10;x=133300000;
#10;x=133310000;
#10;x=133320000;
#10;x=133330000;
#10;x=133340000;
#10;x=133350000;
#10;x=133360000;
#10;x=133370000;
#10;x=133380000;
#10;x=133390000;
#10;x=133400000;
#10;x=133410000;
#10;x=133420000;
#10;x=133430000;
#10;x=133440000;
#10;x=133450000;
#10;x=133460000;
#10;x=133470000;
#10;x=133480000;
#10;x=133490000;
#10;x=133500000;
#10;x=133510000;
#10;x=133520000;
#10;x=133530000;
#10;x=133540000;
#10;x=133550000;
#10;x=133560000;
#10;x=133570000;
#10;x=133580000;
#10;x=133590000;
#10;x=133600000;
#10;x=133610000;
#10;x=133620000;
#10;x=133630000;
#10;x=133640000;
#10;x=133650000;
#10;x=133660000;
#10;x=133670000;
#10;x=133680000;
#10;x=133690000;
#10;x=133700000;
#10;x=133710000;
#10;x=133720000;
#10;x=133730000;
#10;x=133740000;
#10;x=133750000;
#10;x=133760000;
#10;x=133770000;
#10;x=133780000;
#10;x=133790000;
#10;x=133800000;
#10;x=133810000;
#10;x=133820000;
#10;x=133830000;
#10;x=133840000;
#10;x=133850000;
#10;x=133860000;
#10;x=133870000;
#10;x=133880000;
#10;x=133890000;
#10;x=133900000;
#10;x=133910000;
#10;x=133920000;
#10;x=133930000;
#10;x=133940000;
#10;x=133950000;
#10;x=133960000;
#10;x=133970000;
#10;x=133980000;
#10;x=133990000;
#10;x=134000000;
#10;x=134010000;
#10;x=134020000;
#10;x=134030000;
#10;x=134040000;
#10;x=134050000;
#10;x=134060000;
#10;x=134070000;
#10;x=134080000;
#10;x=134090000;
#10;x=134100000;
#10;x=134110000;
#10;x=134120000;
#10;x=134130000;
#10;x=134140000;
#10;x=134150000;
#10;x=134160000;
#10;x=134170000;
#10;x=134180000;
#10;x=134190000;
#10;x=134200000;
#10;x=134210000;
#10;x=134220000;
#10;x=134230000;
#10;x=134240000;
#10;x=134250000;
#10;x=134260000;
#10;x=134270000;
#10;x=134280000;
#10;x=134290000;
#10;x=134300000;
#10;x=134310000;
#10;x=134320000;
#10;x=134330000;
#10;x=134340000;
#10;x=134350000;
#10;x=134360000;
#10;x=134370000;
#10;x=134380000;
#10;x=134390000;
#10;x=134400000;
#10;x=134410000;
#10;x=134420000;
#10;x=134430000;
#10;x=134440000;
#10;x=134450000;
#10;x=134460000;
#10;x=134470000;
#10;x=134480000;
#10;x=134490000;
#10;x=134500000;
#10;x=134510000;
#10;x=134520000;
#10;x=134530000;
#10;x=134540000;
#10;x=134550000;
#10;x=134560000;
#10;x=134570000;
#10;x=134580000;
#10;x=134590000;
#10;x=134600000;
#10;x=134610000;
#10;x=134620000;
#10;x=134630000;
#10;x=134640000;
#10;x=134650000;
#10;x=134660000;
#10;x=134670000;
#10;x=134680000;
#10;x=134690000;
#10;x=134700000;
#10;x=134710000;
#10;x=134720000;
#10;x=134730000;
#10;x=134740000;
#10;x=134750000;
#10;x=134760000;
#10;x=134770000;
#10;x=134780000;
#10;x=134790000;
#10;x=134800000;
#10;x=134810000;
#10;x=134820000;
#10;x=134830000;
#10;x=134840000;
#10;x=134850000;
#10;x=134860000;
#10;x=134870000;
#10;x=134880000;
#10;x=134890000;
#10;x=134900000;
#10;x=134910000;
#10;x=134920000;
#10;x=134930000;
#10;x=134940000;
#10;x=134950000;
#10;x=134960000;
#10;x=134970000;
#10;x=134980000;
#10;x=134990000;
#10;x=135000000;
#10;x=135010000;
#10;x=135020000;
#10;x=135030000;
#10;x=135040000;
#10;x=135050000;
#10;x=135060000;
#10;x=135070000;
#10;x=135080000;
#10;x=135090000;
#10;x=135100000;
#10;x=135110000;
#10;x=135120000;
#10;x=135130000;
#10;x=135140000;
#10;x=135150000;
#10;x=135160000;
#10;x=135170000;
#10;x=135180000;
#10;x=135190000;
#10;x=135200000;
#10;x=135210000;
#10;x=135220000;
#10;x=135230000;
#10;x=135240000;
#10;x=135250000;
#10;x=135260000;
#10;x=135270000;
#10;x=135280000;
#10;x=135290000;
#10;x=135300000;
#10;x=135310000;
#10;x=135320000;
#10;x=135330000;
#10;x=135340000;
#10;x=135350000;
#10;x=135360000;
#10;x=135370000;
#10;x=135380000;
#10;x=135390000;
#10;x=135400000;
#10;x=135410000;
#10;x=135420000;
#10;x=135430000;
#10;x=135440000;
#10;x=135450000;
#10;x=135460000;
#10;x=135470000;
#10;x=135480000;
#10;x=135490000;
#10;x=135500000;
#10;x=135510000;
#10;x=135520000;
#10;x=135530000;
#10;x=135540000;
#10;x=135550000;
#10;x=135560000;
#10;x=135570000;
#10;x=135580000;
#10;x=135590000;
#10;x=135600000;
#10;x=135610000;
#10;x=135620000;
#10;x=135630000;
#10;x=135640000;
#10;x=135650000;
#10;x=135660000;
#10;x=135670000;
#10;x=135680000;
#10;x=135690000;
#10;x=135700000;
#10;x=135710000;
#10;x=135720000;
#10;x=135730000;
#10;x=135740000;
#10;x=135750000;
#10;x=135760000;
#10;x=135770000;
#10;x=135780000;
#10;x=135790000;
#10;x=135800000;
#10;x=135810000;
#10;x=135820000;
#10;x=135830000;
#10;x=135840000;
#10;x=135850000;
#10;x=135860000;
#10;x=135870000;
#10;x=135880000;
#10;x=135890000;
#10;x=135900000;
#10;x=135910000;
#10;x=135920000;
#10;x=135930000;
#10;x=135940000;
#10;x=135950000;
#10;x=135960000;
#10;x=135970000;
#10;x=135980000;
#10;x=135990000;
#10;x=136000000;
#10;x=136010000;
#10;x=136020000;
#10;x=136030000;
#10;x=136040000;
#10;x=136050000;
#10;x=136060000;
#10;x=136070000;
#10;x=136080000;
#10;x=136090000;
#10;x=136100000;
#10;x=136110000;
#10;x=136120000;
#10;x=136130000;
#10;x=136140000;
#10;x=136150000;
#10;x=136160000;
#10;x=136170000;
#10;x=136180000;
#10;x=136190000;
#10;x=136200000;
#10;x=136210000;
#10;x=136220000;
#10;x=136230000;
#10;x=136240000;
#10;x=136250000;
#10;x=136260000;
#10;x=136270000;
#10;x=136280000;
#10;x=136290000;
#10;x=136300000;
#10;x=136310000;
#10;x=136320000;
#10;x=136330000;
#10;x=136340000;
#10;x=136350000;
#10;x=136360000;
#10;x=136370000;
#10;x=136380000;
#10;x=136390000;
#10;x=136400000;
#10;x=136410000;
#10;x=136420000;
#10;x=136430000;
#10;x=136440000;
#10;x=136450000;
#10;x=136460000;
#10;x=136470000;
#10;x=136480000;
#10;x=136490000;
#10;x=136500000;
#10;x=136510000;
#10;x=136520000;
#10;x=136530000;
#10;x=136540000;
#10;x=136550000;
#10;x=136560000;
#10;x=136570000;
#10;x=136580000;
#10;x=136590000;
#10;x=136600000;
#10;x=136610000;
#10;x=136620000;
#10;x=136630000;
#10;x=136640000;
#10;x=136650000;
#10;x=136660000;
#10;x=136670000;
#10;x=136680000;
#10;x=136690000;
#10;x=136700000;
#10;x=136710000;
#10;x=136720000;
#10;x=136730000;
#10;x=136740000;
#10;x=136750000;
#10;x=136760000;
#10;x=136770000;
#10;x=136780000;
#10;x=136790000;
#10;x=136800000;
#10;x=136810000;
#10;x=136820000;
#10;x=136830000;
#10;x=136840000;
#10;x=136850000;
#10;x=136860000;
#10;x=136870000;
#10;x=136880000;
#10;x=136890000;
#10;x=136900000;
#10;x=136910000;
#10;x=136920000;
#10;x=136930000;
#10;x=136940000;
#10;x=136950000;
#10;x=136960000;
#10;x=136970000;
#10;x=136980000;
#10;x=136990000;
#10;x=137000000;
#10;x=137010000;
#10;x=137020000;
#10;x=137030000;
#10;x=137040000;
#10;x=137050000;
#10;x=137060000;
#10;x=137070000;
#10;x=137080000;
#10;x=137090000;
#10;x=137100000;
#10;x=137110000;
#10;x=137120000;
#10;x=137130000;
#10;x=137140000;
#10;x=137150000;
#10;x=137160000;
#10;x=137170000;
#10;x=137180000;
#10;x=137190000;
#10;x=137200000;
#10;x=137210000;
#10;x=137220000;
#10;x=137230000;
#10;x=137240000;
#10;x=137250000;
#10;x=137260000;
#10;x=137270000;
#10;x=137280000;
#10;x=137290000;
#10;x=137300000;
#10;x=137310000;
#10;x=137320000;
#10;x=137330000;
#10;x=137340000;
#10;x=137350000;
#10;x=137360000;
#10;x=137370000;
#10;x=137380000;
#10;x=137390000;
#10;x=137400000;
#10;x=137410000;
#10;x=137420000;
#10;x=137430000;
#10;x=137440000;
#10;x=137450000;
#10;x=137460000;
#10;x=137470000;
#10;x=137480000;
#10;x=137490000;
#10;x=137500000;
#10;x=137510000;
#10;x=137520000;
#10;x=137530000;
#10;x=137540000;
#10;x=137550000;
#10;x=137560000;
#10;x=137570000;
#10;x=137580000;
#10;x=137590000;
#10;x=137600000;
#10;x=137610000;
#10;x=137620000;
#10;x=137630000;
#10;x=137640000;
#10;x=137650000;
#10;x=137660000;
#10;x=137670000;
#10;x=137680000;
#10;x=137690000;
#10;x=137700000;
#10;x=137710000;
#10;x=137720000;
#10;x=137730000;
#10;x=137740000;
#10;x=137750000;
#10;x=137760000;
#10;x=137770000;
#10;x=137780000;
#10;x=137790000;
#10;x=137800000;
#10;x=137810000;
#10;x=137820000;
#10;x=137830000;
#10;x=137840000;
#10;x=137850000;
#10;x=137860000;
#10;x=137870000;
#10;x=137880000;
#10;x=137890000;
#10;x=137900000;
#10;x=137910000;
#10;x=137920000;
#10;x=137930000;
#10;x=137940000;
#10;x=137950000;
#10;x=137960000;
#10;x=137970000;
#10;x=137980000;
#10;x=137990000;
#10;x=138000000;
#10;x=138010000;
#10;x=138020000;
#10;x=138030000;
#10;x=138040000;
#10;x=138050000;
#10;x=138060000;
#10;x=138070000;
#10;x=138080000;
#10;x=138090000;
#10;x=138100000;
#10;x=138110000;
#10;x=138120000;
#10;x=138130000;
#10;x=138140000;
#10;x=138150000;
#10;x=138160000;
#10;x=138170000;
#10;x=138180000;
#10;x=138190000;
#10;x=138200000;
#10;x=138210000;
#10;x=138220000;
#10;x=138230000;
#10;x=138240000;
#10;x=138250000;
#10;x=138260000;
#10;x=138270000;
#10;x=138280000;
#10;x=138290000;
#10;x=138300000;
#10;x=138310000;
#10;x=138320000;
#10;x=138330000;
#10;x=138340000;
#10;x=138350000;
#10;x=138360000;
#10;x=138370000;
#10;x=138380000;
#10;x=138390000;
#10;x=138400000;
#10;x=138410000;
#10;x=138420000;
#10;x=138430000;
#10;x=138440000;
#10;x=138450000;
#10;x=138460000;
#10;x=138470000;
#10;x=138480000;
#10;x=138490000;
#10;x=138500000;
#10;x=138510000;
#10;x=138520000;
#10;x=138530000;
#10;x=138540000;
#10;x=138550000;
#10;x=138560000;
#10;x=138570000;
#10;x=138580000;
#10;x=138590000;
#10;x=138600000;
#10;x=138610000;
#10;x=138620000;
#10;x=138630000;
#10;x=138640000;
#10;x=138650000;
#10;x=138660000;
#10;x=138670000;
#10;x=138680000;
#10;x=138690000;
#10;x=138700000;
#10;x=138710000;
#10;x=138720000;
#10;x=138730000;
#10;x=138740000;
#10;x=138750000;
#10;x=138760000;
#10;x=138770000;
#10;x=138780000;
#10;x=138790000;
#10;x=138800000;
#10;x=138810000;
#10;x=138820000;
#10;x=138830000;
#10;x=138840000;
#10;x=138850000;
#10;x=138860000;
#10;x=138870000;
#10;x=138880000;
#10;x=138890000;
#10;x=138900000;
#10;x=138910000;
#10;x=138920000;
#10;x=138930000;
#10;x=138940000;
#10;x=138950000;
#10;x=138960000;
#10;x=138970000;
#10;x=138980000;
#10;x=138990000;
#10;x=139000000;
#10;x=139010000;
#10;x=139020000;
#10;x=139030000;
#10;x=139040000;
#10;x=139050000;
#10;x=139060000;
#10;x=139070000;
#10;x=139080000;
#10;x=139090000;
#10;x=139100000;
#10;x=139110000;
#10;x=139120000;
#10;x=139130000;
#10;x=139140000;
#10;x=139150000;
#10;x=139160000;
#10;x=139170000;
#10;x=139180000;
#10;x=139190000;
#10;x=139200000;
#10;x=139210000;
#10;x=139220000;
#10;x=139230000;
#10;x=139240000;
#10;x=139250000;
#10;x=139260000;
#10;x=139270000;
#10;x=139280000;
#10;x=139290000;
#10;x=139300000;
#10;x=139310000;
#10;x=139320000;
#10;x=139330000;
#10;x=139340000;
#10;x=139350000;
#10;x=139360000;
#10;x=139370000;
#10;x=139380000;
#10;x=139390000;
#10;x=139400000;
#10;x=139410000;
#10;x=139420000;
#10;x=139430000;
#10;x=139440000;
#10;x=139450000;
#10;x=139460000;
#10;x=139470000;
#10;x=139480000;
#10;x=139490000;
#10;x=139500000;
#10;x=139510000;
#10;x=139520000;
#10;x=139530000;
#10;x=139540000;
#10;x=139550000;
#10;x=139560000;
#10;x=139570000;
#10;x=139580000;
#10;x=139590000;
#10;x=139600000;
#10;x=139610000;
#10;x=139620000;
#10;x=139630000;
#10;x=139640000;
#10;x=139650000;
#10;x=139660000;
#10;x=139670000;
#10;x=139680000;
#10;x=139690000;
#10;x=139700000;
#10;x=139710000;
#10;x=139720000;
#10;x=139730000;
#10;x=139740000;
#10;x=139750000;
#10;x=139760000;
#10;x=139770000;
#10;x=139780000;
#10;x=139790000;
#10;x=139800000;
#10;x=139810000;
#10;x=139820000;
#10;x=139830000;
#10;x=139840000;
#10;x=139850000;
#10;x=139860000;
#10;x=139870000;
#10;x=139880000;
#10;x=139890000;
#10;x=139900000;
#10;x=139910000;
#10;x=139920000;
#10;x=139930000;
#10;x=139940000;
#10;x=139950000;
#10;x=139960000;
#10;x=139970000;
#10;x=139980000;
#10;x=139990000;
#10;x=140000000;
#10;x=140010000;
#10;x=140020000;
#10;x=140030000;
#10;x=140040000;
#10;x=140050000;
#10;x=140060000;
#10;x=140070000;
#10;x=140080000;
#10;x=140090000;
#10;x=140100000;
#10;x=140110000;
#10;x=140120000;
#10;x=140130000;
#10;x=140140000;
#10;x=140150000;
#10;x=140160000;
#10;x=140170000;
#10;x=140180000;
#10;x=140190000;
#10;x=140200000;
#10;x=140210000;
#10;x=140220000;
#10;x=140230000;
#10;x=140240000;
#10;x=140250000;
#10;x=140260000;
#10;x=140270000;
#10;x=140280000;
#10;x=140290000;
#10;x=140300000;
#10;x=140310000;
#10;x=140320000;
#10;x=140330000;
#10;x=140340000;
#10;x=140350000;
#10;x=140360000;
#10;x=140370000;
#10;x=140380000;
#10;x=140390000;
#10;x=140400000;
#10;x=140410000;
#10;x=140420000;
#10;x=140430000;
#10;x=140440000;
#10;x=140450000;
#10;x=140460000;
#10;x=140470000;
#10;x=140480000;
#10;x=140490000;
#10;x=140500000;
#10;x=140510000;
#10;x=140520000;
#10;x=140530000;
#10;x=140540000;
#10;x=140550000;
#10;x=140560000;
#10;x=140570000;
#10;x=140580000;
#10;x=140590000;
#10;x=140600000;
#10;x=140610000;
#10;x=140620000;
#10;x=140630000;
#10;x=140640000;
#10;x=140650000;
#10;x=140660000;
#10;x=140670000;
#10;x=140680000;
#10;x=140690000;
#10;x=140700000;
#10;x=140710000;
#10;x=140720000;
#10;x=140730000;
#10;x=140740000;
#10;x=140750000;
#10;x=140760000;
#10;x=140770000;
#10;x=140780000;
#10;x=140790000;
#10;x=140800000;
#10;x=140810000;
#10;x=140820000;
#10;x=140830000;
#10;x=140840000;
#10;x=140850000;
#10;x=140860000;
#10;x=140870000;
#10;x=140880000;
#10;x=140890000;
#10;x=140900000;
#10;x=140910000;
#10;x=140920000;
#10;x=140930000;
#10;x=140940000;
#10;x=140950000;
#10;x=140960000;
#10;x=140970000;
#10;x=140980000;
#10;x=140990000;
#10;x=141000000;
#10;x=141010000;
#10;x=141020000;
#10;x=141030000;
#10;x=141040000;
#10;x=141050000;
#10;x=141060000;
#10;x=141070000;
#10;x=141080000;
#10;x=141090000;
#10;x=141100000;
#10;x=141110000;
#10;x=141120000;
#10;x=141130000;
#10;x=141140000;
#10;x=141150000;
#10;x=141160000;
#10;x=141170000;
#10;x=141180000;
#10;x=141190000;
#10;x=141200000;
#10;x=141210000;
#10;x=141220000;
#10;x=141230000;
#10;x=141240000;
#10;x=141250000;
#10;x=141260000;
#10;x=141270000;
#10;x=141280000;
#10;x=141290000;
#10;x=141300000;
#10;x=141310000;
#10;x=141320000;
#10;x=141330000;
#10;x=141340000;
#10;x=141350000;
#10;x=141360000;
#10;x=141370000;
#10;x=141380000;
#10;x=141390000;
#10;x=141400000;
#10;x=141410000;
#10;x=141420000;
#10;x=141430000;
#10;x=141440000;
#10;x=141450000;
#10;x=141460000;
#10;x=141470000;
#10;x=141480000;
#10;x=141490000;
#10;x=141500000;
#10;x=141510000;
#10;x=141520000;
#10;x=141530000;
#10;x=141540000;
#10;x=141550000;
#10;x=141560000;
#10;x=141570000;
#10;x=141580000;
#10;x=141590000;
#10;x=141600000;
#10;x=141610000;
#10;x=141620000;
#10;x=141630000;
#10;x=141640000;
#10;x=141650000;
#10;x=141660000;
#10;x=141670000;
#10;x=141680000;
#10;x=141690000;
#10;x=141700000;
#10;x=141710000;
#10;x=141720000;
#10;x=141730000;
#10;x=141740000;
#10;x=141750000;
#10;x=141760000;
#10;x=141770000;
#10;x=141780000;
#10;x=141790000;
#10;x=141800000;
#10;x=141810000;
#10;x=141820000;
#10;x=141830000;
#10;x=141840000;
#10;x=141850000;
#10;x=141860000;
#10;x=141870000;
#10;x=141880000;
#10;x=141890000;
#10;x=141900000;
#10;x=141910000;
#10;x=141920000;
#10;x=141930000;
#10;x=141940000;
#10;x=141950000;
#10;x=141960000;
#10;x=141970000;
#10;x=141980000;
#10;x=141990000;
#10;x=142000000;
#10;x=142010000;
#10;x=142020000;
#10;x=142030000;
#10;x=142040000;
#10;x=142050000;
#10;x=142060000;
#10;x=142070000;
#10;x=142080000;
#10;x=142090000;
#10;x=142100000;
#10;x=142110000;
#10;x=142120000;
#10;x=142130000;
#10;x=142140000;
#10;x=142150000;
#10;x=142160000;
#10;x=142170000;
#10;x=142180000;
#10;x=142190000;
#10;x=142200000;
#10;x=142210000;
#10;x=142220000;
#10;x=142230000;
#10;x=142240000;
#10;x=142250000;
#10;x=142260000;
#10;x=142270000;
#10;x=142280000;
#10;x=142290000;
#10;x=142300000;
#10;x=142310000;
#10;x=142320000;
#10;x=142330000;
#10;x=142340000;
#10;x=142350000;
#10;x=142360000;
#10;x=142370000;
#10;x=142380000;
#10;x=142390000;
#10;x=142400000;
#10;x=142410000;
#10;x=142420000;
#10;x=142430000;
#10;x=142440000;
#10;x=142450000;
#10;x=142460000;
#10;x=142470000;
#10;x=142480000;
#10;x=142490000;
#10;x=142500000;
#10;x=142510000;
#10;x=142520000;
#10;x=142530000;
#10;x=142540000;
#10;x=142550000;
#10;x=142560000;
#10;x=142570000;
#10;x=142580000;
#10;x=142590000;
#10;x=142600000;
#10;x=142610000;
#10;x=142620000;
#10;x=142630000;
#10;x=142640000;
#10;x=142650000;
#10;x=142660000;
#10;x=142670000;
#10;x=142680000;
#10;x=142690000;
#10;x=142700000;
#10;x=142710000;
#10;x=142720000;
#10;x=142730000;
#10;x=142740000;
#10;x=142750000;
#10;x=142760000;
#10;x=142770000;
#10;x=142780000;
#10;x=142790000;
#10;x=142800000;
#10;x=142810000;
#10;x=142820000;
#10;x=142830000;
#10;x=142840000;
#10;x=142850000;
#10;x=142860000;
#10;x=142870000;
#10;x=142880000;
#10;x=142890000;
#10;x=142900000;
#10;x=142910000;
#10;x=142920000;
#10;x=142930000;
#10;x=142940000;
#10;x=142950000;
#10;x=142960000;
#10;x=142970000;
#10;x=142980000;
#10;x=142990000;
#10;x=143000000;
#10;x=143010000;
#10;x=143020000;
#10;x=143030000;
#10;x=143040000;
#10;x=143050000;
#10;x=143060000;
#10;x=143070000;
#10;x=143080000;
#10;x=143090000;
#10;x=143100000;
#10;x=143110000;
#10;x=143120000;
#10;x=143130000;
#10;x=143140000;
#10;x=143150000;
#10;x=143160000;
#10;x=143170000;
#10;x=143180000;
#10;x=143190000;
#10;x=143200000;
#10;x=143210000;
#10;x=143220000;
#10;x=143230000;
#10;x=143240000;
#10;x=143250000;
#10;x=143260000;
#10;x=143270000;
#10;x=143280000;
#10;x=143290000;
#10;x=143300000;
#10;x=143310000;
#10;x=143320000;
#10;x=143330000;
#10;x=143340000;
#10;x=143350000;
#10;x=143360000;
#10;x=143370000;
#10;x=143380000;
#10;x=143390000;
#10;x=143400000;
#10;x=143410000;
#10;x=143420000;
#10;x=143430000;
#10;x=143440000;
#10;x=143450000;
#10;x=143460000;
#10;x=143470000;
#10;x=143480000;
#10;x=143490000;
#10;x=143500000;
#10;x=143510000;
#10;x=143520000;
#10;x=143530000;
#10;x=143540000;
#10;x=143550000;
#10;x=143560000;
#10;x=143570000;
#10;x=143580000;
#10;x=143590000;
#10;x=143600000;
#10;x=143610000;
#10;x=143620000;
#10;x=143630000;
#10;x=143640000;
#10;x=143650000;
#10;x=143660000;
#10;x=143670000;
#10;x=143680000;
#10;x=143690000;
#10;x=143700000;
#10;x=143710000;
#10;x=143720000;
#10;x=143730000;
#10;x=143740000;
#10;x=143750000;
#10;x=143760000;
#10;x=143770000;
#10;x=143780000;
#10;x=143790000;
#10;x=143800000;
#10;x=143810000;
#10;x=143820000;
#10;x=143830000;
#10;x=143840000;
#10;x=143850000;
#10;x=143860000;
#10;x=143870000;
#10;x=143880000;
#10;x=143890000;
#10;x=143900000;
#10;x=143910000;
#10;x=143920000;
#10;x=143930000;
#10;x=143940000;
#10;x=143950000;
#10;x=143960000;
#10;x=143970000;
#10;x=143980000;
#10;x=143990000;
#10;x=144000000;
#10;x=144010000;
#10;x=144020000;
#10;x=144030000;
#10;x=144040000;
#10;x=144050000;
#10;x=144060000;
#10;x=144070000;
#10;x=144080000;
#10;x=144090000;
#10;x=144100000;
#10;x=144110000;
#10;x=144120000;
#10;x=144130000;
#10;x=144140000;
#10;x=144150000;
#10;x=144160000;
#10;x=144170000;
#10;x=144180000;
#10;x=144190000;
#10;x=144200000;
#10;x=144210000;
#10;x=144220000;
#10;x=144230000;
#10;x=144240000;
#10;x=144250000;
#10;x=144260000;
#10;x=144270000;
#10;x=144280000;
#10;x=144290000;
#10;x=144300000;
#10;x=144310000;
#10;x=144320000;
#10;x=144330000;
#10;x=144340000;
#10;x=144350000;
#10;x=144360000;
#10;x=144370000;
#10;x=144380000;
#10;x=144390000;
#10;x=144400000;
#10;x=144410000;
#10;x=144420000;
#10;x=144430000;
#10;x=144440000;
#10;x=144450000;
#10;x=144460000;
#10;x=144470000;
#10;x=144480000;
#10;x=144490000;
#10;x=144500000;
#10;x=144510000;
#10;x=144520000;
#10;x=144530000;
#10;x=144540000;
#10;x=144550000;
#10;x=144560000;
#10;x=144570000;
#10;x=144580000;
#10;x=144590000;
#10;x=144600000;
#10;x=144610000;
#10;x=144620000;
#10;x=144630000;
#10;x=144640000;
#10;x=144650000;
#10;x=144660000;
#10;x=144670000;
#10;x=144680000;
#10;x=144690000;
#10;x=144700000;
#10;x=144710000;
#10;x=144720000;
#10;x=144730000;
#10;x=144740000;
#10;x=144750000;
#10;x=144760000;
#10;x=144770000;
#10;x=144780000;
#10;x=144790000;
#10;x=144800000;
#10;x=144810000;
#10;x=144820000;
#10;x=144830000;
#10;x=144840000;
#10;x=144850000;
#10;x=144860000;
#10;x=144870000;
#10;x=144880000;
#10;x=144890000;
#10;x=144900000;
#10;x=144910000;
#10;x=144920000;
#10;x=144930000;
#10;x=144940000;
#10;x=144950000;
#10;x=144960000;
#10;x=144970000;
#10;x=144980000;
#10;x=144990000;
#10;x=145000000;
#10;x=145010000;
#10;x=145020000;
#10;x=145030000;
#10;x=145040000;
#10;x=145050000;
#10;x=145060000;
#10;x=145070000;
#10;x=145080000;
#10;x=145090000;
#10;x=145100000;
#10;x=145110000;
#10;x=145120000;
#10;x=145130000;
#10;x=145140000;
#10;x=145150000;
#10;x=145160000;
#10;x=145170000;
#10;x=145180000;
#10;x=145190000;
#10;x=145200000;
#10;x=145210000;
#10;x=145220000;
#10;x=145230000;
#10;x=145240000;
#10;x=145250000;
#10;x=145260000;
#10;x=145270000;
#10;x=145280000;
#10;x=145290000;
#10;x=145300000;
#10;x=145310000;
#10;x=145320000;
#10;x=145330000;
#10;x=145340000;
#10;x=145350000;
#10;x=145360000;
#10;x=145370000;
#10;x=145380000;
#10;x=145390000;
#10;x=145400000;
#10;x=145410000;
#10;x=145420000;
#10;x=145430000;
#10;x=145440000;
#10;x=145450000;
#10;x=145460000;
#10;x=145470000;
#10;x=145480000;
#10;x=145490000;
#10;x=145500000;
#10;x=145510000;
#10;x=145520000;
#10;x=145530000;
#10;x=145540000;
#10;x=145550000;
#10;x=145560000;
#10;x=145570000;
#10;x=145580000;
#10;x=145590000;
#10;x=145600000;
#10;x=145610000;
#10;x=145620000;
#10;x=145630000;
#10;x=145640000;
#10;x=145650000;
#10;x=145660000;
#10;x=145670000;
#10;x=145680000;
#10;x=145690000;
#10;x=145700000;
#10;x=145710000;
#10;x=145720000;
#10;x=145730000;
#10;x=145740000;
#10;x=145750000;
#10;x=145760000;
#10;x=145770000;
#10;x=145780000;
#10;x=145790000;
#10;x=145800000;
#10;x=145810000;
#10;x=145820000;
#10;x=145830000;
#10;x=145840000;
#10;x=145850000;
#10;x=145860000;
#10;x=145870000;
#10;x=145880000;
#10;x=145890000;
#10;x=145900000;
#10;x=145910000;
#10;x=145920000;
#10;x=145930000;
#10;x=145940000;
#10;x=145950000;
#10;x=145960000;
#10;x=145970000;
#10;x=145980000;
#10;x=145990000;
#10;x=146000000;
#10;x=146010000;
#10;x=146020000;
#10;x=146030000;
#10;x=146040000;
#10;x=146050000;
#10;x=146060000;
#10;x=146070000;
#10;x=146080000;
#10;x=146090000;
#10;x=146100000;
#10;x=146110000;
#10;x=146120000;
#10;x=146130000;
#10;x=146140000;
#10;x=146150000;
#10;x=146160000;
#10;x=146170000;
#10;x=146180000;
#10;x=146190000;
#10;x=146200000;
#10;x=146210000;
#10;x=146220000;
#10;x=146230000;
#10;x=146240000;
#10;x=146250000;
#10;x=146260000;
#10;x=146270000;
#10;x=146280000;
#10;x=146290000;
#10;x=146300000;
#10;x=146310000;
#10;x=146320000;
#10;x=146330000;
#10;x=146340000;
#10;x=146350000;
#10;x=146360000;
#10;x=146370000;
#10;x=146380000;
#10;x=146390000;
#10;x=146400000;
#10;x=146410000;
#10;x=146420000;
#10;x=146430000;
#10;x=146440000;
#10;x=146450000;
#10;x=146460000;
#10;x=146470000;
#10;x=146480000;
#10;x=146490000;
#10;x=146500000;
#10;x=146510000;
#10;x=146520000;
#10;x=146530000;
#10;x=146540000;
#10;x=146550000;
#10;x=146560000;
#10;x=146570000;
#10;x=146580000;
#10;x=146590000;
#10;x=146600000;
#10;x=146610000;
#10;x=146620000;
#10;x=146630000;
#10;x=146640000;
#10;x=146650000;
#10;x=146660000;
#10;x=146670000;
#10;x=146680000;
#10;x=146690000;
#10;x=146700000;
#10;x=146710000;
#10;x=146720000;
#10;x=146730000;
#10;x=146740000;
#10;x=146750000;
#10;x=146760000;
#10;x=146770000;
#10;x=146780000;
#10;x=146790000;
#10;x=146800000;
#10;x=146810000;
#10;x=146820000;
#10;x=146830000;
#10;x=146840000;
#10;x=146850000;
#10;x=146860000;
#10;x=146870000;
#10;x=146880000;
#10;x=146890000;
#10;x=146900000;
#10;x=146910000;
#10;x=146920000;
#10;x=146930000;
#10;x=146940000;
#10;x=146950000;
#10;x=146960000;
#10;x=146970000;
#10;x=146980000;
#10;x=146990000;
#10;x=147000000;
#10;x=147010000;
#10;x=147020000;
#10;x=147030000;
#10;x=147040000;
#10;x=147050000;
#10;x=147060000;
#10;x=147070000;
#10;x=147080000;
#10;x=147090000;
#10;x=147100000;
#10;x=147110000;
#10;x=147120000;
#10;x=147130000;
#10;x=147140000;
#10;x=147150000;
#10;x=147160000;
#10;x=147170000;
#10;x=147180000;
#10;x=147190000;
#10;x=147200000;
#10;x=147210000;
#10;x=147220000;
#10;x=147230000;
#10;x=147240000;
#10;x=147250000;
#10;x=147260000;
#10;x=147270000;
#10;x=147280000;
#10;x=147290000;
#10;x=147300000;
#10;x=147310000;
#10;x=147320000;
#10;x=147330000;
#10;x=147340000;
#10;x=147350000;
#10;x=147360000;
#10;x=147370000;
#10;x=147380000;
#10;x=147390000;
#10;x=147400000;
#10;x=147410000;
#10;x=147420000;
#10;x=147430000;
#10;x=147440000;
#10;x=147450000;
#10;x=147460000;
#10;x=147470000;
#10;x=147480000;
#10;x=147490000;
#10;x=147500000;
#10;x=147510000;
#10;x=147520000;
#10;x=147530000;
#10;x=147540000;
#10;x=147550000;
#10;x=147560000;
#10;x=147570000;
#10;x=147580000;
#10;x=147590000;
#10;x=147600000;
#10;x=147610000;
#10;x=147620000;
#10;x=147630000;
#10;x=147640000;
#10;x=147650000;
#10;x=147660000;
#10;x=147670000;
#10;x=147680000;
#10;x=147690000;
#10;x=147700000;
#10;x=147710000;
#10;x=147720000;
#10;x=147730000;
#10;x=147740000;
#10;x=147750000;
#10;x=147760000;
#10;x=147770000;
#10;x=147780000;
#10;x=147790000;
#10;x=147800000;
#10;x=147810000;
#10;x=147820000;
#10;x=147830000;
#10;x=147840000;
#10;x=147850000;
#10;x=147860000;
#10;x=147870000;
#10;x=147880000;
#10;x=147890000;
#10;x=147900000;
#10;x=147910000;
#10;x=147920000;
#10;x=147930000;
#10;x=147940000;
#10;x=147950000;
#10;x=147960000;
#10;x=147970000;
#10;x=147980000;
#10;x=147990000;
#10;x=148000000;
#10;x=148010000;
#10;x=148020000;
#10;x=148030000;
#10;x=148040000;
#10;x=148050000;
#10;x=148060000;
#10;x=148070000;
#10;x=148080000;
#10;x=148090000;
#10;x=148100000;
#10;x=148110000;
#10;x=148120000;
#10;x=148130000;
#10;x=148140000;
#10;x=148150000;
#10;x=148160000;
#10;x=148170000;
#10;x=148180000;
#10;x=148190000;
#10;x=148200000;
#10;x=148210000;
#10;x=148220000;
#10;x=148230000;
#10;x=148240000;
#10;x=148250000;
#10;x=148260000;
#10;x=148270000;
#10;x=148280000;
#10;x=148290000;
#10;x=148300000;
#10;x=148310000;
#10;x=148320000;
#10;x=148330000;
#10;x=148340000;
#10;x=148350000;
#10;x=148360000;
#10;x=148370000;
#10;x=148380000;
#10;x=148390000;
#10;x=148400000;
#10;x=148410000;
#10;x=148420000;
#10;x=148430000;
#10;x=148440000;
#10;x=148450000;
#10;x=148460000;
#10;x=148470000;
#10;x=148480000;
#10;x=148490000;
#10;x=148500000;
#10;x=148510000;
#10;x=148520000;
#10;x=148530000;
#10;x=148540000;
#10;x=148550000;
#10;x=148560000;
#10;x=148570000;
#10;x=148580000;
#10;x=148590000;
#10;x=148600000;
#10;x=148610000;
#10;x=148620000;
#10;x=148630000;
#10;x=148640000;
#10;x=148650000;
#10;x=148660000;
#10;x=148670000;
#10;x=148680000;
#10;x=148690000;
#10;x=148700000;
#10;x=148710000;
#10;x=148720000;
#10;x=148730000;
#10;x=148740000;
#10;x=148750000;
#10;x=148760000;
#10;x=148770000;
#10;x=148780000;
#10;x=148790000;
#10;x=148800000;
#10;x=148810000;
#10;x=148820000;
#10;x=148830000;
#10;x=148840000;
#10;x=148850000;
#10;x=148860000;
#10;x=148870000;
#10;x=148880000;
#10;x=148890000;
#10;x=148900000;
#10;x=148910000;
#10;x=148920000;
#10;x=148930000;
#10;x=148940000;
#10;x=148950000;
#10;x=148960000;
#10;x=148970000;
#10;x=148980000;
#10;x=148990000;
#10;x=149000000;
#10;x=149010000;
#10;x=149020000;
#10;x=149030000;
#10;x=149040000;
#10;x=149050000;
#10;x=149060000;
#10;x=149070000;
#10;x=149080000;
#10;x=149090000;
#10;x=149100000;
#10;x=149110000;
#10;x=149120000;
#10;x=149130000;
#10;x=149140000;
#10;x=149150000;
#10;x=149160000;
#10;x=149170000;
#10;x=149180000;
#10;x=149190000;
#10;x=149200000;
#10;x=149210000;
#10;x=149220000;
#10;x=149230000;
#10;x=149240000;
#10;x=149250000;
#10;x=149260000;
#10;x=149270000;
#10;x=149280000;
#10;x=149290000;
#10;x=149300000;
#10;x=149310000;
#10;x=149320000;
#10;x=149330000;
#10;x=149340000;
#10;x=149350000;
#10;x=149360000;
#10;x=149370000;
#10;x=149380000;
#10;x=149390000;
#10;x=149400000;
#10;x=149410000;
#10;x=149420000;
#10;x=149430000;
#10;x=149440000;
#10;x=149450000;
#10;x=149460000;
#10;x=149470000;
#10;x=149480000;
#10;x=149490000;
#10;x=149500000;
#10;x=149510000;
#10;x=149520000;
#10;x=149530000;
#10;x=149540000;
#10;x=149550000;
#10;x=149560000;
#10;x=149570000;
#10;x=149580000;
#10;x=149590000;
#10;x=149600000;
#10;x=149610000;
#10;x=149620000;
#10;x=149630000;
#10;x=149640000;
#10;x=149650000;
#10;x=149660000;
#10;x=149670000;
#10;x=149680000;
#10;x=149690000;
#10;x=149700000;
#10;x=149710000;
#10;x=149720000;
#10;x=149730000;
#10;x=149740000;
#10;x=149750000;
#10;x=149760000;
#10;x=149770000;
#10;x=149780000;
#10;x=149790000;
#10;x=149800000;
#10;x=149810000;
#10;x=149820000;
#10;x=149830000;
#10;x=149840000;
#10;x=149850000;
#10;x=149860000;
#10;x=149870000;
#10;x=149880000;
#10;x=149890000;
#10;x=149900000;
#10;x=149910000;
#10;x=149920000;
#10;x=149930000;
#10;x=149940000;
#10;x=149950000;
#10;x=149960000;
#10;x=149970000;
#10;x=149980000;
#10;x=149990000;
#10;x=150000000;
#10;x=150010000;
#10;x=150020000;
#10;x=150030000;
#10;x=150040000;
#10;x=150050000;
#10;x=150060000;
#10;x=150070000;
#10;x=150080000;
#10;x=150090000;
#10;x=150100000;
#10;x=150110000;
#10;x=150120000;
#10;x=150130000;
#10;x=150140000;
#10;x=150150000;
#10;x=150160000;
#10;x=150170000;
#10;x=150180000;
#10;x=150190000;
#10;x=150200000;
#10;x=150210000;
#10;x=150220000;
#10;x=150230000;
#10;x=150240000;
#10;x=150250000;
#10;x=150260000;
#10;x=150270000;
#10;x=150280000;
#10;x=150290000;
#10;x=150300000;
#10;x=150310000;
#10;x=150320000;
#10;x=150330000;
#10;x=150340000;
#10;x=150350000;
#10;x=150360000;
#10;x=150370000;
#10;x=150380000;
#10;x=150390000;
#10;x=150400000;
#10;x=150410000;
#10;x=150420000;
#10;x=150430000;
#10;x=150440000;
#10;x=150450000;
#10;x=150460000;
#10;x=150470000;
#10;x=150480000;
#10;x=150490000;
#10;x=150500000;
#10;x=150510000;
#10;x=150520000;
#10;x=150530000;
#10;x=150540000;
#10;x=150550000;
#10;x=150560000;
#10;x=150570000;
#10;x=150580000;
#10;x=150590000;
#10;x=150600000;
#10;x=150610000;
#10;x=150620000;
#10;x=150630000;
#10;x=150640000;
#10;x=150650000;
#10;x=150660000;
#10;x=150670000;
#10;x=150680000;
#10;x=150690000;
#10;x=150700000;
#10;x=150710000;
#10;x=150720000;
#10;x=150730000;
#10;x=150740000;
#10;x=150750000;
#10;x=150760000;
#10;x=150770000;
#10;x=150780000;
#10;x=150790000;
#10;x=150800000;
#10;x=150810000;
#10;x=150820000;
#10;x=150830000;
#10;x=150840000;
#10;x=150850000;
#10;x=150860000;
#10;x=150870000;
#10;x=150880000;
#10;x=150890000;
#10;x=150900000;
#10;x=150910000;
#10;x=150920000;
#10;x=150930000;
#10;x=150940000;
#10;x=150950000;
#10;x=150960000;
#10;x=150970000;
#10;x=150980000;
#10;x=150990000;
#10;x=151000000;
#10;x=151010000;
#10;x=151020000;
#10;x=151030000;
#10;x=151040000;
#10;x=151050000;
#10;x=151060000;
#10;x=151070000;
#10;x=151080000;
#10;x=151090000;
#10;x=151100000;
#10;x=151110000;
#10;x=151120000;
#10;x=151130000;
#10;x=151140000;
#10;x=151150000;
#10;x=151160000;
#10;x=151170000;
#10;x=151180000;
#10;x=151190000;
#10;x=151200000;
#10;x=151210000;
#10;x=151220000;
#10;x=151230000;
#10;x=151240000;
#10;x=151250000;
#10;x=151260000;
#10;x=151270000;
#10;x=151280000;
#10;x=151290000;
#10;x=151300000;
#10;x=151310000;
#10;x=151320000;
#10;x=151330000;
#10;x=151340000;
#10;x=151350000;
#10;x=151360000;
#10;x=151370000;
#10;x=151380000;
#10;x=151390000;
#10;x=151400000;
#10;x=151410000;
#10;x=151420000;
#10;x=151430000;
#10;x=151440000;
#10;x=151450000;
#10;x=151460000;
#10;x=151470000;
#10;x=151480000;
#10;x=151490000;
#10;x=151500000;
#10;x=151510000;
#10;x=151520000;
#10;x=151530000;
#10;x=151540000;
#10;x=151550000;
#10;x=151560000;
#10;x=151570000;
#10;x=151580000;
#10;x=151590000;
#10;x=151600000;
#10;x=151610000;
#10;x=151620000;
#10;x=151630000;
#10;x=151640000;
#10;x=151650000;
#10;x=151660000;
#10;x=151670000;
#10;x=151680000;
#10;x=151690000;
#10;x=151700000;
#10;x=151710000;
#10;x=151720000;
#10;x=151730000;
#10;x=151740000;
#10;x=151750000;
#10;x=151760000;
#10;x=151770000;
#10;x=151780000;
#10;x=151790000;
#10;x=151800000;
#10;x=151810000;
#10;x=151820000;
#10;x=151830000;
#10;x=151840000;
#10;x=151850000;
#10;x=151860000;
#10;x=151870000;
#10;x=151880000;
#10;x=151890000;
#10;x=151900000;
#10;x=151910000;
#10;x=151920000;
#10;x=151930000;
#10;x=151940000;
#10;x=151950000;
#10;x=151960000;
#10;x=151970000;
#10;x=151980000;
#10;x=151990000;
#10;x=152000000;
#10;x=152010000;
#10;x=152020000;
#10;x=152030000;
#10;x=152040000;
#10;x=152050000;
#10;x=152060000;
#10;x=152070000;
#10;x=152080000;
#10;x=152090000;
#10;x=152100000;
#10;x=152110000;
#10;x=152120000;
#10;x=152130000;
#10;x=152140000;
#10;x=152150000;
#10;x=152160000;
#10;x=152170000;
#10;x=152180000;
#10;x=152190000;
#10;x=152200000;
#10;x=152210000;
#10;x=152220000;
#10;x=152230000;
#10;x=152240000;
#10;x=152250000;
#10;x=152260000;
#10;x=152270000;
#10;x=152280000;
#10;x=152290000;
#10;x=152300000;
#10;x=152310000;
#10;x=152320000;
#10;x=152330000;
#10;x=152340000;
#10;x=152350000;
#10;x=152360000;
#10;x=152370000;
#10;x=152380000;
#10;x=152390000;
#10;x=152400000;
#10;x=152410000;
#10;x=152420000;
#10;x=152430000;
#10;x=152440000;
#10;x=152450000;
#10;x=152460000;
#10;x=152470000;
#10;x=152480000;
#10;x=152490000;
#10;x=152500000;
#10;x=152510000;
#10;x=152520000;
#10;x=152530000;
#10;x=152540000;
#10;x=152550000;
#10;x=152560000;
#10;x=152570000;
#10;x=152580000;
#10;x=152590000;
#10;x=152600000;
#10;x=152610000;
#10;x=152620000;
#10;x=152630000;
#10;x=152640000;
#10;x=152650000;
#10;x=152660000;
#10;x=152670000;
#10;x=152680000;
#10;x=152690000;
#10;x=152700000;
#10;x=152710000;
#10;x=152720000;
#10;x=152730000;
#10;x=152740000;
#10;x=152750000;
#10;x=152760000;
#10;x=152770000;
#10;x=152780000;
#10;x=152790000;
#10;x=152800000;
#10;x=152810000;
#10;x=152820000;
#10;x=152830000;
#10;x=152840000;
#10;x=152850000;
#10;x=152860000;
#10;x=152870000;
#10;x=152880000;
#10;x=152890000;
#10;x=152900000;
#10;x=152910000;
#10;x=152920000;
#10;x=152930000;
#10;x=152940000;
#10;x=152950000;
#10;x=152960000;
#10;x=152970000;
#10;x=152980000;
#10;x=152990000;
#10;x=153000000;
#10;x=153010000;
#10;x=153020000;
#10;x=153030000;
#10;x=153040000;
#10;x=153050000;
#10;x=153060000;
#10;x=153070000;
#10;x=153080000;
#10;x=153090000;
#10;x=153100000;
#10;x=153110000;
#10;x=153120000;
#10;x=153130000;
#10;x=153140000;
#10;x=153150000;
#10;x=153160000;
#10;x=153170000;
#10;x=153180000;
#10;x=153190000;
#10;x=153200000;
#10;x=153210000;
#10;x=153220000;
#10;x=153230000;
#10;x=153240000;
#10;x=153250000;
#10;x=153260000;
#10;x=153270000;
#10;x=153280000;
#10;x=153290000;
#10;x=153300000;
#10;x=153310000;
#10;x=153320000;
#10;x=153330000;
#10;x=153340000;
#10;x=153350000;
#10;x=153360000;
#10;x=153370000;
#10;x=153380000;
#10;x=153390000;
#10;x=153400000;
#10;x=153410000;
#10;x=153420000;
#10;x=153430000;
#10;x=153440000;
#10;x=153450000;
#10;x=153460000;
#10;x=153470000;
#10;x=153480000;
#10;x=153490000;
#10;x=153500000;
#10;x=153510000;
#10;x=153520000;
#10;x=153530000;
#10;x=153540000;
#10;x=153550000;
#10;x=153560000;
#10;x=153570000;
#10;x=153580000;
#10;x=153590000;
#10;x=153600000;
#10;x=153610000;
#10;x=153620000;
#10;x=153630000;
#10;x=153640000;
#10;x=153650000;
#10;x=153660000;
#10;x=153670000;
#10;x=153680000;
#10;x=153690000;
#10;x=153700000;
#10;x=153710000;
#10;x=153720000;
#10;x=153730000;
#10;x=153740000;
#10;x=153750000;
#10;x=153760000;
#10;x=153770000;
#10;x=153780000;
#10;x=153790000;
#10;x=153800000;
#10;x=153810000;
#10;x=153820000;
#10;x=153830000;
#10;x=153840000;
#10;x=153850000;
#10;x=153860000;
#10;x=153870000;
#10;x=153880000;
#10;x=153890000;
#10;x=153900000;
#10;x=153910000;
#10;x=153920000;
#10;x=153930000;
#10;x=153940000;
#10;x=153950000;
#10;x=153960000;
#10;x=153970000;
#10;x=153980000;
#10;x=153990000;
#10;x=154000000;
#10;x=154010000;
#10;x=154020000;
#10;x=154030000;
#10;x=154040000;
#10;x=154050000;
#10;x=154060000;
#10;x=154070000;
#10;x=154080000;
#10;x=154090000;
#10;x=154100000;
#10;x=154110000;
#10;x=154120000;
#10;x=154130000;
#10;x=154140000;
#10;x=154150000;
#10;x=154160000;
#10;x=154170000;
#10;x=154180000;
#10;x=154190000;
#10;x=154200000;
#10;x=154210000;
#10;x=154220000;
#10;x=154230000;
#10;x=154240000;
#10;x=154250000;
#10;x=154260000;
#10;x=154270000;
#10;x=154280000;
#10;x=154290000;
#10;x=154300000;
#10;x=154310000;
#10;x=154320000;
#10;x=154330000;
#10;x=154340000;
#10;x=154350000;
#10;x=154360000;
#10;x=154370000;
#10;x=154380000;
#10;x=154390000;
#10;x=154400000;
#10;x=154410000;
#10;x=154420000;
#10;x=154430000;
#10;x=154440000;
#10;x=154450000;
#10;x=154460000;
#10;x=154470000;
#10;x=154480000;
#10;x=154490000;
#10;x=154500000;
#10;x=154510000;
#10;x=154520000;
#10;x=154530000;
#10;x=154540000;
#10;x=154550000;
#10;x=154560000;
#10;x=154570000;
#10;x=154580000;
#10;x=154590000;
#10;x=154600000;
#10;x=154610000;
#10;x=154620000;
#10;x=154630000;
#10;x=154640000;
#10;x=154650000;
#10;x=154660000;
#10;x=154670000;
#10;x=154680000;
#10;x=154690000;
#10;x=154700000;
#10;x=154710000;
#10;x=154720000;
#10;x=154730000;
#10;x=154740000;
#10;x=154750000;
#10;x=154760000;
#10;x=154770000;
#10;x=154780000;
#10;x=154790000;
#10;x=154800000;
#10;x=154810000;
#10;x=154820000;
#10;x=154830000;
#10;x=154840000;
#10;x=154850000;
#10;x=154860000;
#10;x=154870000;
#10;x=154880000;
#10;x=154890000;
#10;x=154900000;
#10;x=154910000;
#10;x=154920000;
#10;x=154930000;
#10;x=154940000;
#10;x=154950000;
#10;x=154960000;
#10;x=154970000;
#10;x=154980000;
#10;x=154990000;
#10;x=155000000;
#10;x=155010000;
#10;x=155020000;
#10;x=155030000;
#10;x=155040000;
#10;x=155050000;
#10;x=155060000;
#10;x=155070000;
#10;x=155080000;
#10;x=155090000;
#10;x=155100000;
#10;x=155110000;
#10;x=155120000;
#10;x=155130000;
#10;x=155140000;
#10;x=155150000;
#10;x=155160000;
#10;x=155170000;
#10;x=155180000;
#10;x=155190000;
#10;x=155200000;
#10;x=155210000;
#10;x=155220000;
#10;x=155230000;
#10;x=155240000;
#10;x=155250000;
#10;x=155260000;
#10;x=155270000;
#10;x=155280000;
#10;x=155290000;
#10;x=155300000;
#10;x=155310000;
#10;x=155320000;
#10;x=155330000;
#10;x=155340000;
#10;x=155350000;
#10;x=155360000;
#10;x=155370000;
#10;x=155380000;
#10;x=155390000;
#10;x=155400000;
#10;x=155410000;
#10;x=155420000;
#10;x=155430000;
#10;x=155440000;
#10;x=155450000;
#10;x=155460000;
#10;x=155470000;
#10;x=155480000;
#10;x=155490000;
#10;x=155500000;
#10;x=155510000;
#10;x=155520000;
#10;x=155530000;
#10;x=155540000;
#10;x=155550000;
#10;x=155560000;
#10;x=155570000;
#10;x=155580000;
#10;x=155590000;
#10;x=155600000;
#10;x=155610000;
#10;x=155620000;
#10;x=155630000;
#10;x=155640000;
#10;x=155650000;
#10;x=155660000;
#10;x=155670000;
#10;x=155680000;
#10;x=155690000;
#10;x=155700000;
#10;x=155710000;
#10;x=155720000;
#10;x=155730000;
#10;x=155740000;
#10;x=155750000;
#10;x=155760000;
#10;x=155770000;
#10;x=155780000;
#10;x=155790000;
#10;x=155800000;
#10;x=155810000;
#10;x=155820000;
#10;x=155830000;
#10;x=155840000;
#10;x=155850000;
#10;x=155860000;
#10;x=155870000;
#10;x=155880000;
#10;x=155890000;
#10;x=155900000;
#10;x=155910000;
#10;x=155920000;
#10;x=155930000;
#10;x=155940000;
#10;x=155950000;
#10;x=155960000;
#10;x=155970000;
#10;x=155980000;
#10;x=155990000;
#10;x=156000000;
#10;x=156010000;
#10;x=156020000;
#10;x=156030000;
#10;x=156040000;
#10;x=156050000;
#10;x=156060000;
#10;x=156070000;
#10;x=156080000;
#10;x=156090000;
#10;x=156100000;
#10;x=156110000;
#10;x=156120000;
#10;x=156130000;
#10;x=156140000;
#10;x=156150000;
#10;x=156160000;
#10;x=156170000;
#10;x=156180000;
#10;x=156190000;
#10;x=156200000;
#10;x=156210000;
#10;x=156220000;
#10;x=156230000;
#10;x=156240000;
#10;x=156250000;
#10;x=156260000;
#10;x=156270000;
#10;x=156280000;
#10;x=156290000;
#10;x=156300000;
#10;x=156310000;
#10;x=156320000;
#10;x=156330000;
#10;x=156340000;
#10;x=156350000;
#10;x=156360000;
#10;x=156370000;
#10;x=156380000;
#10;x=156390000;
#10;x=156400000;
#10;x=156410000;
#10;x=156420000;
#10;x=156430000;
#10;x=156440000;
#10;x=156450000;
#10;x=156460000;
#10;x=156470000;
#10;x=156480000;
#10;x=156490000;
#10;x=156500000;
#10;x=156510000;
#10;x=156520000;
#10;x=156530000;
#10;x=156540000;
#10;x=156550000;
#10;x=156560000;
#10;x=156570000;
#10;x=156580000;
#10;x=156590000;
#10;x=156600000;
#10;x=156610000;
#10;x=156620000;
#10;x=156630000;
#10;x=156640000;
#10;x=156650000;
#10;x=156660000;
#10;x=156670000;
#10;x=156680000;
#10;x=156690000;
#10;x=156700000;
#10;x=156710000;
#10;x=156720000;
#10;x=156730000;
#10;x=156740000;
#10;x=156750000;
#10;x=156760000;
#10;x=156770000;
#10;x=156780000;
#10;x=156790000;
#10;x=156800000;
#10;x=156810000;
#10;x=156820000;
#10;x=156830000;
#10;x=156840000;
#10;x=156850000;
#10;x=156860000;
#10;x=156870000;
#10;x=156880000;
#10;x=156890000;
#10;x=156900000;
#10;x=156910000;
#10;x=156920000;
#10;x=156930000;
#10;x=156940000;
#10;x=156950000;
#10;x=156960000;
#10;x=156970000;
#10;x=156980000;
#10;x=156990000;
#10;x=157000000;
#10;x=157010000;
#10;x=157020000;
#10;x=157030000;
#10;x=157040000;
#10;x=157050000;
#10;x=157060000;
#10;x=157070000;
#10;x=157080000;
#10;x=157090000;
#10;x=157100000;
#10;x=157110000;
#10;x=157120000;
#10;x=157130000;
#10;x=157140000;
#10;x=157150000;
#10;x=157160000;
#10;x=157170000;
#10;x=157180000;
#10;x=157190000;
#10;x=157200000;
#10;x=157210000;
#10;x=157220000;
#10;x=157230000;
#10;x=157240000;
#10;x=157250000;
#10;x=157260000;
#10;x=157270000;
#10;x=157280000;
#10;x=157290000;
#10;x=157300000;
#10;x=157310000;
#10;x=157320000;
#10;x=157330000;
#10;x=157340000;
#10;x=157350000;
#10;x=157360000;
#10;x=157370000;
#10;x=157380000;
#10;x=157390000;
#10;x=157400000;
#10;x=157410000;
#10;x=157420000;
#10;x=157430000;
#10;x=157440000;
#10;x=157450000;
#10;x=157460000;
#10;x=157470000;
#10;x=157480000;
#10;x=157490000;
#10;x=157500000;
#10;x=157510000;
#10;x=157520000;
#10;x=157530000;
#10;x=157540000;
#10;x=157550000;
#10;x=157560000;
#10;x=157570000;
#10;x=157580000;
#10;x=157590000;
#10;x=157600000;
#10;x=157610000;
#10;x=157620000;
#10;x=157630000;
#10;x=157640000;
#10;x=157650000;
#10;x=157660000;
#10;x=157670000;
#10;x=157680000;
#10;x=157690000;
#10;x=157700000;
#10;x=157710000;
#10;x=157720000;
#10;x=157730000;
#10;x=157740000;
#10;x=157750000;
#10;x=157760000;
#10;x=157770000;
#10;x=157780000;
#10;x=157790000;
#10;x=157800000;
#10;x=157810000;
#10;x=157820000;
#10;x=157830000;
#10;x=157840000;
#10;x=157850000;
#10;x=157860000;
#10;x=157870000;
#10;x=157880000;
#10;x=157890000;
#10;x=157900000;
#10;x=157910000;
#10;x=157920000;
#10;x=157930000;
#10;x=157940000;
#10;x=157950000;
#10;x=157960000;
#10;x=157970000;
#10;x=157980000;
#10;x=157990000;
#10;x=158000000;
#10;x=158010000;
#10;x=158020000;
#10;x=158030000;
#10;x=158040000;
#10;x=158050000;
#10;x=158060000;
#10;x=158070000;
#10;x=158080000;
#10;x=158090000;
#10;x=158100000;
#10;x=158110000;
#10;x=158120000;
#10;x=158130000;
#10;x=158140000;
#10;x=158150000;
#10;x=158160000;
#10;x=158170000;
#10;x=158180000;
#10;x=158190000;
#10;x=158200000;
#10;x=158210000;
#10;x=158220000;
#10;x=158230000;
#10;x=158240000;
#10;x=158250000;
#10;x=158260000;
#10;x=158270000;
#10;x=158280000;
#10;x=158290000;
#10;x=158300000;
#10;x=158310000;
#10;x=158320000;
#10;x=158330000;
#10;x=158340000;
#10;x=158350000;
#10;x=158360000;
#10;x=158370000;
#10;x=158380000;
#10;x=158390000;
#10;x=158400000;
#10;x=158410000;
#10;x=158420000;
#10;x=158430000;
#10;x=158440000;
#10;x=158450000;
#10;x=158460000;
#10;x=158470000;
#10;x=158480000;
#10;x=158490000;
#10;x=158500000;
#10;x=158510000;
#10;x=158520000;
#10;x=158530000;
#10;x=158540000;
#10;x=158550000;
#10;x=158560000;
#10;x=158570000;
#10;x=158580000;
#10;x=158590000;
#10;x=158600000;
#10;x=158610000;
#10;x=158620000;
#10;x=158630000;
#10;x=158640000;
#10;x=158650000;
#10;x=158660000;
#10;x=158670000;
#10;x=158680000;
#10;x=158690000;
#10;x=158700000;
#10;x=158710000;
#10;x=158720000;
#10;x=158730000;
#10;x=158740000;
#10;x=158750000;
#10;x=158760000;
#10;x=158770000;
#10;x=158780000;
#10;x=158790000;
#10;x=158800000;
#10;x=158810000;
#10;x=158820000;
#10;x=158830000;
#10;x=158840000;
#10;x=158850000;
#10;x=158860000;
#10;x=158870000;
#10;x=158880000;
#10;x=158890000;
#10;x=158900000;
#10;x=158910000;
#10;x=158920000;
#10;x=158930000;
#10;x=158940000;
#10;x=158950000;
#10;x=158960000;
#10;x=158970000;
#10;x=158980000;
#10;x=158990000;
#10;x=159000000;
#10;x=159010000;
#10;x=159020000;
#10;x=159030000;
#10;x=159040000;
#10;x=159050000;
#10;x=159060000;
#10;x=159070000;
#10;x=159080000;
#10;x=159090000;
#10;x=159100000;
#10;x=159110000;
#10;x=159120000;
#10;x=159130000;
#10;x=159140000;
#10;x=159150000;
#10;x=159160000;
#10;x=159170000;
#10;x=159180000;
#10;x=159190000;
#10;x=159200000;
#10;x=159210000;
#10;x=159220000;
#10;x=159230000;
#10;x=159240000;
#10;x=159250000;
#10;x=159260000;
#10;x=159270000;
#10;x=159280000;
#10;x=159290000;
#10;x=159300000;
#10;x=159310000;
#10;x=159320000;
#10;x=159330000;
#10;x=159340000;
#10;x=159350000;
#10;x=159360000;
#10;x=159370000;
#10;x=159380000;
#10;x=159390000;
#10;x=159400000;
#10;x=159410000;
#10;x=159420000;
#10;x=159430000;
#10;x=159440000;
#10;x=159450000;
#10;x=159460000;
#10;x=159470000;
#10;x=159480000;
#10;x=159490000;
#10;x=159500000;
#10;x=159510000;
#10;x=159520000;
#10;x=159530000;
#10;x=159540000;
#10;x=159550000;
#10;x=159560000;
#10;x=159570000;
#10;x=159580000;
#10;x=159590000;
#10;x=159600000;
#10;x=159610000;
#10;x=159620000;
#10;x=159630000;
#10;x=159640000;
#10;x=159650000;
#10;x=159660000;
#10;x=159670000;
#10;x=159680000;
#10;x=159690000;
#10;x=159700000;
#10;x=159710000;
#10;x=159720000;
#10;x=159730000;
#10;x=159740000;
#10;x=159750000;
#10;x=159760000;
#10;x=159770000;
#10;x=159780000;
#10;x=159790000;
#10;x=159800000;
#10;x=159810000;
#10;x=159820000;
#10;x=159830000;
#10;x=159840000;
#10;x=159850000;
#10;x=159860000;
#10;x=159870000;
#10;x=159880000;
#10;x=159890000;
#10;x=159900000;
#10;x=159910000;
#10;x=159920000;
#10;x=159930000;
#10;x=159940000;
#10;x=159950000;
#10;x=159960000;
#10;x=159970000;
#10;x=159980000;
#10;x=159990000;
#10;x=160000000;
#10;x=160010000;
#10;x=160020000;
#10;x=160030000;
#10;x=160040000;
#10;x=160050000;
#10;x=160060000;
#10;x=160070000;
#10;x=160080000;
#10;x=160090000;
#10;x=160100000;
#10;x=160110000;
#10;x=160120000;
#10;x=160130000;
#10;x=160140000;
#10;x=160150000;
#10;x=160160000;
#10;x=160170000;
#10;x=160180000;
#10;x=160190000;
#10;x=160200000;
#10;x=160210000;
#10;x=160220000;
#10;x=160230000;
#10;x=160240000;
#10;x=160250000;
#10;x=160260000;
#10;x=160270000;
#10;x=160280000;
#10;x=160290000;
#10;x=160300000;
#10;x=160310000;
#10;x=160320000;
#10;x=160330000;
#10;x=160340000;
#10;x=160350000;
#10;x=160360000;
#10;x=160370000;
#10;x=160380000;
#10;x=160390000;
#10;x=160400000;
#10;x=160410000;
#10;x=160420000;
#10;x=160430000;
#10;x=160440000;
#10;x=160450000;
#10;x=160460000;
#10;x=160470000;
#10;x=160480000;
#10;x=160490000;
#10;x=160500000;
#10;x=160510000;
#10;x=160520000;
#10;x=160530000;
#10;x=160540000;
#10;x=160550000;
#10;x=160560000;
#10;x=160570000;
#10;x=160580000;
#10;x=160590000;
#10;x=160600000;
#10;x=160610000;
#10;x=160620000;
#10;x=160630000;
#10;x=160640000;
#10;x=160650000;
#10;x=160660000;
#10;x=160670000;
#10;x=160680000;
#10;x=160690000;
#10;x=160700000;
#10;x=160710000;
#10;x=160720000;
#10;x=160730000;
#10;x=160740000;
#10;x=160750000;
#10;x=160760000;
#10;x=160770000;
#10;x=160780000;
#10;x=160790000;
#10;x=160800000;
#10;x=160810000;
#10;x=160820000;
#10;x=160830000;
#10;x=160840000;
#10;x=160850000;
#10;x=160860000;
#10;x=160870000;
#10;x=160880000;
#10;x=160890000;
#10;x=160900000;
#10;x=160910000;
#10;x=160920000;
#10;x=160930000;
#10;x=160940000;
#10;x=160950000;
#10;x=160960000;
#10;x=160970000;
#10;x=160980000;
#10;x=160990000;
#10;x=161000000;
#10;x=161010000;
#10;x=161020000;
#10;x=161030000;
#10;x=161040000;
#10;x=161050000;
#10;x=161060000;
#10;x=161070000;
#10;x=161080000;
#10;x=161090000;
#10;x=161100000;
#10;x=161110000;
#10;x=161120000;
#10;x=161130000;
#10;x=161140000;
#10;x=161150000;
#10;x=161160000;
#10;x=161170000;
#10;x=161180000;
#10;x=161190000;
#10;x=161200000;
#10;x=161210000;
#10;x=161220000;
#10;x=161230000;
#10;x=161240000;
#10;x=161250000;
#10;x=161260000;
#10;x=161270000;
#10;x=161280000;
#10;x=161290000;
#10;x=161300000;
#10;x=161310000;
#10;x=161320000;
#10;x=161330000;
#10;x=161340000;
#10;x=161350000;
#10;x=161360000;
#10;x=161370000;
#10;x=161380000;
#10;x=161390000;
#10;x=161400000;
#10;x=161410000;
#10;x=161420000;
#10;x=161430000;
#10;x=161440000;
#10;x=161450000;
#10;x=161460000;
#10;x=161470000;
#10;x=161480000;
#10;x=161490000;
#10;x=161500000;
#10;x=161510000;
#10;x=161520000;
#10;x=161530000;
#10;x=161540000;
#10;x=161550000;
#10;x=161560000;
#10;x=161570000;
#10;x=161580000;
#10;x=161590000;
#10;x=161600000;
#10;x=161610000;
#10;x=161620000;
#10;x=161630000;
#10;x=161640000;
#10;x=161650000;
#10;x=161660000;
#10;x=161670000;
#10;x=161680000;
#10;x=161690000;
#10;x=161700000;
#10;x=161710000;
#10;x=161720000;
#10;x=161730000;
#10;x=161740000;
#10;x=161750000;
#10;x=161760000;
#10;x=161770000;
#10;x=161780000;
#10;x=161790000;
#10;x=161800000;
#10;x=161810000;
#10;x=161820000;
#10;x=161830000;
#10;x=161840000;
#10;x=161850000;
#10;x=161860000;
#10;x=161870000;
#10;x=161880000;
#10;x=161890000;
#10;x=161900000;
#10;x=161910000;
#10;x=161920000;
#10;x=161930000;
#10;x=161940000;
#10;x=161950000;
#10;x=161960000;
#10;x=161970000;
#10;x=161980000;
#10;x=161990000;
#10;x=162000000;
#10;x=162010000;
#10;x=162020000;
#10;x=162030000;
#10;x=162040000;
#10;x=162050000;
#10;x=162060000;
#10;x=162070000;
#10;x=162080000;
#10;x=162090000;
#10;x=162100000;
#10;x=162110000;
#10;x=162120000;
#10;x=162130000;
#10;x=162140000;
#10;x=162150000;
#10;x=162160000;
#10;x=162170000;
#10;x=162180000;
#10;x=162190000;
#10;x=162200000;
#10;x=162210000;
#10;x=162220000;
#10;x=162230000;
#10;x=162240000;
#10;x=162250000;
#10;x=162260000;
#10;x=162270000;
#10;x=162280000;
#10;x=162290000;
#10;x=162300000;
#10;x=162310000;
#10;x=162320000;
#10;x=162330000;
#10;x=162340000;
#10;x=162350000;
#10;x=162360000;
#10;x=162370000;
#10;x=162380000;
#10;x=162390000;
#10;x=162400000;
#10;x=162410000;
#10;x=162420000;
#10;x=162430000;
#10;x=162440000;
#10;x=162450000;
#10;x=162460000;
#10;x=162470000;
#10;x=162480000;
#10;x=162490000;
#10;x=162500000;
#10;x=162510000;
#10;x=162520000;
#10;x=162530000;
#10;x=162540000;
#10;x=162550000;
#10;x=162560000;
#10;x=162570000;
#10;x=162580000;
#10;x=162590000;
#10;x=162600000;
#10;x=162610000;
#10;x=162620000;
#10;x=162630000;
#10;x=162640000;
#10;x=162650000;
#10;x=162660000;
#10;x=162670000;
#10;x=162680000;
#10;x=162690000;
#10;x=162700000;
#10;x=162710000;
#10;x=162720000;
#10;x=162730000;
#10;x=162740000;
#10;x=162750000;
#10;x=162760000;
#10;x=162770000;
#10;x=162780000;
#10;x=162790000;
#10;x=162800000;
#10;x=162810000;
#10;x=162820000;
#10;x=162830000;
#10;x=162840000;
#10;x=162850000;
#10;x=162860000;
#10;x=162870000;
#10;x=162880000;
#10;x=162890000;
#10;x=162900000;
#10;x=162910000;
#10;x=162920000;
#10;x=162930000;
#10;x=162940000;
#10;x=162950000;
#10;x=162960000;
#10;x=162970000;
#10;x=162980000;
#10;x=162990000;
#10;x=163000000;
#10;x=163010000;
#10;x=163020000;
#10;x=163030000;
#10;x=163040000;
#10;x=163050000;
#10;x=163060000;
#10;x=163070000;
#10;x=163080000;
#10;x=163090000;
#10;x=163100000;
#10;x=163110000;
#10;x=163120000;
#10;x=163130000;
#10;x=163140000;
#10;x=163150000;
#10;x=163160000;
#10;x=163170000;
#10;x=163180000;
#10;x=163190000;
#10;x=163200000;
#10;x=163210000;
#10;x=163220000;
#10;x=163230000;
#10;x=163240000;
#10;x=163250000;
#10;x=163260000;
#10;x=163270000;
#10;x=163280000;
#10;x=163290000;
#10;x=163300000;
#10;x=163310000;
#10;x=163320000;
#10;x=163330000;
#10;x=163340000;
#10;x=163350000;
#10;x=163360000;
#10;x=163370000;
#10;x=163380000;
#10;x=163390000;
#10;x=163400000;
#10;x=163410000;
#10;x=163420000;
#10;x=163430000;
#10;x=163440000;
#10;x=163450000;
#10;x=163460000;
#10;x=163470000;
#10;x=163480000;
#10;x=163490000;
#10;x=163500000;
#10;x=163510000;
#10;x=163520000;
#10;x=163530000;
#10;x=163540000;
#10;x=163550000;
#10;x=163560000;
#10;x=163570000;
#10;x=163580000;
#10;x=163590000;
#10;x=163600000;
#10;x=163610000;
#10;x=163620000;
#10;x=163630000;
#10;x=163640000;
#10;x=163650000;
#10;x=163660000;
#10;x=163670000;
#10;x=163680000;
#10;x=163690000;
#10;x=163700000;
#10;x=163710000;
#10;x=163720000;
#10;x=163730000;
#10;x=163740000;
#10;x=163750000;
#10;x=163760000;
#10;x=163770000;
#10;x=163780000;
#10;x=163790000;
#10;x=163800000;
#10;x=163810000;
#10;x=163820000;
#10;x=163830000;
#10;x=163840000;
#10;x=163850000;
#10;x=163860000;
#10;x=163870000;
#10;x=163880000;
#10;x=163890000;
#10;x=163900000;
#10;x=163910000;
#10;x=163920000;
#10;x=163930000;
#10;x=163940000;
#10;x=163950000;
#10;x=163960000;
#10;x=163970000;
#10;x=163980000;
#10;x=163990000;
#10;x=164000000;
#10;x=164010000;
#10;x=164020000;
#10;x=164030000;
#10;x=164040000;
#10;x=164050000;
#10;x=164060000;
#10;x=164070000;
#10;x=164080000;
#10;x=164090000;
#10;x=164100000;
#10;x=164110000;
#10;x=164120000;
#10;x=164130000;
#10;x=164140000;
#10;x=164150000;
#10;x=164160000;
#10;x=164170000;
#10;x=164180000;
#10;x=164190000;
#10;x=164200000;
#10;x=164210000;
#10;x=164220000;
#10;x=164230000;
#10;x=164240000;
#10;x=164250000;
#10;x=164260000;
#10;x=164270000;
#10;x=164280000;
#10;x=164290000;
#10;x=164300000;
#10;x=164310000;
#10;x=164320000;
#10;x=164330000;
#10;x=164340000;
#10;x=164350000;
#10;x=164360000;
#10;x=164370000;
#10;x=164380000;
#10;x=164390000;
#10;x=164400000;
#10;x=164410000;
#10;x=164420000;
#10;x=164430000;
#10;x=164440000;
#10;x=164450000;
#10;x=164460000;
#10;x=164470000;
#10;x=164480000;
#10;x=164490000;
#10;x=164500000;
#10;x=164510000;
#10;x=164520000;
#10;x=164530000;
#10;x=164540000;
#10;x=164550000;
#10;x=164560000;
#10;x=164570000;
#10;x=164580000;
#10;x=164590000;
#10;x=164600000;
#10;x=164610000;
#10;x=164620000;
#10;x=164630000;
#10;x=164640000;
#10;x=164650000;
#10;x=164660000;
#10;x=164670000;
#10;x=164680000;
#10;x=164690000;
#10;x=164700000;
#10;x=164710000;
#10;x=164720000;
#10;x=164730000;
#10;x=164740000;
#10;x=164750000;
#10;x=164760000;
#10;x=164770000;
#10;x=164780000;
#10;x=164790000;
#10;x=164800000;
#10;x=164810000;
#10;x=164820000;
#10;x=164830000;
#10;x=164840000;
#10;x=164850000;
#10;x=164860000;
#10;x=164870000;
#10;x=164880000;
#10;x=164890000;
#10;x=164900000;
#10;x=164910000;
#10;x=164920000;
#10;x=164930000;
#10;x=164940000;
#10;x=164950000;
#10;x=164960000;
#10;x=164970000;
#10;x=164980000;
#10;x=164990000;
#10;x=165000000;
#10;x=165010000;
#10;x=165020000;
#10;x=165030000;
#10;x=165040000;
#10;x=165050000;
#10;x=165060000;
#10;x=165070000;
#10;x=165080000;
#10;x=165090000;
#10;x=165100000;
#10;x=165110000;
#10;x=165120000;
#10;x=165130000;
#10;x=165140000;
#10;x=165150000;
#10;x=165160000;
#10;x=165170000;
#10;x=165180000;
#10;x=165190000;
#10;x=165200000;
#10;x=165210000;
#10;x=165220000;
#10;x=165230000;
#10;x=165240000;
#10;x=165250000;
#10;x=165260000;
#10;x=165270000;
#10;x=165280000;
#10;x=165290000;
#10;x=165300000;
#10;x=165310000;
#10;x=165320000;
#10;x=165330000;
#10;x=165340000;
#10;x=165350000;
#10;x=165360000;
#10;x=165370000;
#10;x=165380000;
#10;x=165390000;
#10;x=165400000;
#10;x=165410000;
#10;x=165420000;
#10;x=165430000;
#10;x=165440000;
#10;x=165450000;
#10;x=165460000;
#10;x=165470000;
#10;x=165480000;
#10;x=165490000;
#10;x=165500000;
#10;x=165510000;
#10;x=165520000;
#10;x=165530000;
#10;x=165540000;
#10;x=165550000;
#10;x=165560000;
#10;x=165570000;
#10;x=165580000;
#10;x=165590000;
#10;x=165600000;
#10;x=165610000;
#10;x=165620000;
#10;x=165630000;
#10;x=165640000;
#10;x=165650000;
#10;x=165660000;
#10;x=165670000;
#10;x=165680000;
#10;x=165690000;
#10;x=165700000;
#10;x=165710000;
#10;x=165720000;
#10;x=165730000;
#10;x=165740000;
#10;x=165750000;
#10;x=165760000;
#10;x=165770000;
#10;x=165780000;
#10;x=165790000;
#10;x=165800000;
#10;x=165810000;
#10;x=165820000;
#10;x=165830000;
#10;x=165840000;
#10;x=165850000;
#10;x=165860000;
#10;x=165870000;
#10;x=165880000;
#10;x=165890000;
#10;x=165900000;
#10;x=165910000;
#10;x=165920000;
#10;x=165930000;
#10;x=165940000;
#10;x=165950000;
#10;x=165960000;
#10;x=165970000;
#10;x=165980000;
#10;x=165990000;
#10;x=166000000;
#10;x=166010000;
#10;x=166020000;
#10;x=166030000;
#10;x=166040000;
#10;x=166050000;
#10;x=166060000;
#10;x=166070000;
#10;x=166080000;
#10;x=166090000;
#10;x=166100000;
#10;x=166110000;
#10;x=166120000;
#10;x=166130000;
#10;x=166140000;
#10;x=166150000;
#10;x=166160000;
#10;x=166170000;
#10;x=166180000;
#10;x=166190000;
#10;x=166200000;
#10;x=166210000;
#10;x=166220000;
#10;x=166230000;
#10;x=166240000;
#10;x=166250000;
#10;x=166260000;
#10;x=166270000;
#10;x=166280000;
#10;x=166290000;
#10;x=166300000;
#10;x=166310000;
#10;x=166320000;
#10;x=166330000;
#10;x=166340000;
#10;x=166350000;
#10;x=166360000;
#10;x=166370000;
#10;x=166380000;
#10;x=166390000;
#10;x=166400000;
#10;x=166410000;
#10;x=166420000;
#10;x=166430000;
#10;x=166440000;
#10;x=166450000;
#10;x=166460000;
#10;x=166470000;
#10;x=166480000;
#10;x=166490000;
#10;x=166500000;
#10;x=166510000;
#10;x=166520000;
#10;x=166530000;
#10;x=166540000;
#10;x=166550000;
#10;x=166560000;
#10;x=166570000;
#10;x=166580000;
#10;x=166590000;
#10;x=166600000;
#10;x=166610000;
#10;x=166620000;
#10;x=166630000;
#10;x=166640000;
#10;x=166650000;
#10;x=166660000;
#10;x=166670000;
#10;x=166680000;
#10;x=166690000;
#10;x=166700000;
#10;x=166710000;
#10;x=166720000;
#10;x=166730000;
#10;x=166740000;
#10;x=166750000;
#10;x=166760000;
#10;x=166770000;
#10;x=166780000;
#10;x=166790000;
#10;x=166800000;
#10;x=166810000;
#10;x=166820000;
#10;x=166830000;
#10;x=166840000;
#10;x=166850000;
#10;x=166860000;
#10;x=166870000;
#10;x=166880000;
#10;x=166890000;
#10;x=166900000;
#10;x=166910000;
#10;x=166920000;
#10;x=166930000;
#10;x=166940000;
#10;x=166950000;
#10;x=166960000;
#10;x=166970000;
#10;x=166980000;
#10;x=166990000;
#10;x=167000000;
#10;x=167010000;
#10;x=167020000;
#10;x=167030000;
#10;x=167040000;
#10;x=167050000;
#10;x=167060000;
#10;x=167070000;
#10;x=167080000;
#10;x=167090000;
#10;x=167100000;
#10;x=167110000;
#10;x=167120000;
#10;x=167130000;
#10;x=167140000;
#10;x=167150000;
#10;x=167160000;
#10;x=167170000;
#10;x=167180000;
#10;x=167190000;
#10;x=167200000;
#10;x=167210000;
#10;x=167220000;
#10;x=167230000;
#10;x=167240000;
#10;x=167250000;
#10;x=167260000;
#10;x=167270000;
#10;x=167280000;
#10;x=167290000;
#10;x=167300000;
#10;x=167310000;
#10;x=167320000;
#10;x=167330000;
#10;x=167340000;
#10;x=167350000;
#10;x=167360000;
#10;x=167370000;
#10;x=167380000;
#10;x=167390000;
#10;x=167400000;
#10;x=167410000;
#10;x=167420000;
#10;x=167430000;
#10;x=167440000;
#10;x=167450000;
#10;x=167460000;
#10;x=167470000;
#10;x=167480000;
#10;x=167490000;
#10;x=167500000;
#10;x=167510000;
#10;x=167520000;
#10;x=167530000;
#10;x=167540000;
#10;x=167550000;
#10;x=167560000;
#10;x=167570000;
#10;x=167580000;
#10;x=167590000;
#10;x=167600000;
#10;x=167610000;
#10;x=167620000;
#10;x=167630000;
#10;x=167640000;
#10;x=167650000;
#10;x=167660000;
#10;x=167670000;
#10;x=167680000;
#10;x=167690000;
#10;x=167700000;
#10;x=167710000;
#10;x=167720000;
#10;x=167730000;
#10;x=167740000;
#10;x=167750000;
#10;x=167760000;
#10;x=167770000;
#10;x=167780000;
#10;x=167790000;
#10;x=167800000;
#10;x=167810000;
#10;x=167820000;
#10;x=167830000;
#10;x=167840000;
#10;x=167850000;
#10;x=167860000;
#10;x=167870000;
#10;x=167880000;
#10;x=167890000;
#10;x=167900000;
#10;x=167910000;
#10;x=167920000;
#10;x=167930000;
#10;x=167940000;
#10;x=167950000;
#10;x=167960000;
#10;x=167970000;
#10;x=167980000;
#10;x=167990000;
#10;x=168000000;
#10;x=168010000;
#10;x=168020000;
#10;x=168030000;
#10;x=168040000;
#10;x=168050000;
#10;x=168060000;
#10;x=168070000;
#10;x=168080000;
#10;x=168090000;
#10;x=168100000;
#10;x=168110000;
#10;x=168120000;
#10;x=168130000;
#10;x=168140000;
#10;x=168150000;
#10;x=168160000;
#10;x=168170000;
#10;x=168180000;
#10;x=168190000;
#10;x=168200000;
#10;x=168210000;
#10;x=168220000;
#10;x=168230000;
#10;x=168240000;
#10;x=168250000;
#10;x=168260000;
#10;x=168270000;
#10;x=168280000;
#10;x=168290000;
#10;x=168300000;
#10;x=168310000;
#10;x=168320000;
#10;x=168330000;
#10;x=168340000;
#10;x=168350000;
#10;x=168360000;
#10;x=168370000;
#10;x=168380000;
#10;x=168390000;
#10;x=168400000;
#10;x=168410000;
#10;x=168420000;
#10;x=168430000;
#10;x=168440000;
#10;x=168450000;
#10;x=168460000;
#10;x=168470000;
#10;x=168480000;
#10;x=168490000;
#10;x=168500000;
#10;x=168510000;
#10;x=168520000;
#10;x=168530000;
#10;x=168540000;
#10;x=168550000;
#10;x=168560000;
#10;x=168570000;
#10;x=168580000;
#10;x=168590000;
#10;x=168600000;
#10;x=168610000;
#10;x=168620000;
#10;x=168630000;
#10;x=168640000;
#10;x=168650000;
#10;x=168660000;
#10;x=168670000;
#10;x=168680000;
#10;x=168690000;
#10;x=168700000;
#10;x=168710000;
#10;x=168720000;
#10;x=168730000;
#10;x=168740000;
#10;x=168750000;
#10;x=168760000;
#10;x=168770000;
#10;x=168780000;
#10;x=168790000;
#10;x=168800000;
#10;x=168810000;
#10;x=168820000;
#10;x=168830000;
#10;x=168840000;
#10;x=168850000;
#10;x=168860000;
#10;x=168870000;
#10;x=168880000;
#10;x=168890000;
#10;x=168900000;
#10;x=168910000;
#10;x=168920000;
#10;x=168930000;
#10;x=168940000;
#10;x=168950000;
#10;x=168960000;
#10;x=168970000;
#10;x=168980000;
#10;x=168990000;
#10;x=169000000;
#10;x=169010000;
#10;x=169020000;
#10;x=169030000;
#10;x=169040000;
#10;x=169050000;
#10;x=169060000;
#10;x=169070000;
#10;x=169080000;
#10;x=169090000;
#10;x=169100000;
#10;x=169110000;
#10;x=169120000;
#10;x=169130000;
#10;x=169140000;
#10;x=169150000;
#10;x=169160000;
#10;x=169170000;
#10;x=169180000;
#10;x=169190000;
#10;x=169200000;
#10;x=169210000;
#10;x=169220000;
#10;x=169230000;
#10;x=169240000;
#10;x=169250000;
#10;x=169260000;
#10;x=169270000;
#10;x=169280000;
#10;x=169290000;
#10;x=169300000;
#10;x=169310000;
#10;x=169320000;
#10;x=169330000;
#10;x=169340000;
#10;x=169350000;
#10;x=169360000;
#10;x=169370000;
#10;x=169380000;
#10;x=169390000;
#10;x=169400000;
#10;x=169410000;
#10;x=169420000;
#10;x=169430000;
#10;x=169440000;
#10;x=169450000;
#10;x=169460000;
#10;x=169470000;
#10;x=169480000;
#10;x=169490000;
#10;x=169500000;
#10;x=169510000;
#10;x=169520000;
#10;x=169530000;
#10;x=169540000;
#10;x=169550000;
#10;x=169560000;
#10;x=169570000;
#10;x=169580000;
#10;x=169590000;
#10;x=169600000;
#10;x=169610000;
#10;x=169620000;
#10;x=169630000;
#10;x=169640000;
#10;x=169650000;
#10;x=169660000;
#10;x=169670000;
#10;x=169680000;
#10;x=169690000;
#10;x=169700000;
#10;x=169710000;
#10;x=169720000;
#10;x=169730000;
#10;x=169740000;
#10;x=169750000;
#10;x=169760000;
#10;x=169770000;
#10;x=169780000;
#10;x=169790000;
#10;x=169800000;
#10;x=169810000;
#10;x=169820000;
#10;x=169830000;
#10;x=169840000;
#10;x=169850000;
#10;x=169860000;
#10;x=169870000;
#10;x=169880000;
#10;x=169890000;
#10;x=169900000;
#10;x=169910000;
#10;x=169920000;
#10;x=169930000;
#10;x=169940000;
#10;x=169950000;
#10;x=169960000;
#10;x=169970000;
#10;x=169980000;
#10;x=169990000;
#10;x=170000000;
#10;x=170010000;
#10;x=170020000;
#10;x=170030000;
#10;x=170040000;
#10;x=170050000;
#10;x=170060000;
#10;x=170070000;
#10;x=170080000;
#10;x=170090000;
#10;x=170100000;
#10;x=170110000;
#10;x=170120000;
#10;x=170130000;
#10;x=170140000;
#10;x=170150000;
#10;x=170160000;
#10;x=170170000;
#10;x=170180000;
#10;x=170190000;
#10;x=170200000;
#10;x=170210000;
#10;x=170220000;
#10;x=170230000;
#10;x=170240000;
#10;x=170250000;
#10;x=170260000;
#10;x=170270000;
#10;x=170280000;
#10;x=170290000;
#10;x=170300000;
#10;x=170310000;
#10;x=170320000;
#10;x=170330000;
#10;x=170340000;
#10;x=170350000;
#10;x=170360000;
#10;x=170370000;
#10;x=170380000;
#10;x=170390000;
#10;x=170400000;
#10;x=170410000;
#10;x=170420000;
#10;x=170430000;
#10;x=170440000;
#10;x=170450000;
#10;x=170460000;
#10;x=170470000;
#10;x=170480000;
#10;x=170490000;
#10;x=170500000;
#10;x=170510000;
#10;x=170520000;
#10;x=170530000;
#10;x=170540000;
#10;x=170550000;
#10;x=170560000;
#10;x=170570000;
#10;x=170580000;
#10;x=170590000;
#10;x=170600000;
#10;x=170610000;
#10;x=170620000;
#10;x=170630000;
#10;x=170640000;
#10;x=170650000;
#10;x=170660000;
#10;x=170670000;
#10;x=170680000;
#10;x=170690000;
#10;x=170700000;
#10;x=170710000;
#10;x=170720000;
#10;x=170730000;
#10;x=170740000;
#10;x=170750000;
#10;x=170760000;
#10;x=170770000;
#10;x=170780000;
#10;x=170790000;
#10;x=170800000;
#10;x=170810000;
#10;x=170820000;
#10;x=170830000;
#10;x=170840000;
#10;x=170850000;
#10;x=170860000;
#10;x=170870000;
#10;x=170880000;
#10;x=170890000;
#10;x=170900000;
#10;x=170910000;
#10;x=170920000;
#10;x=170930000;
#10;x=170940000;
#10;x=170950000;
#10;x=170960000;
#10;x=170970000;
#10;x=170980000;
#10;x=170990000;
#10;x=171000000;
#10;x=171010000;
#10;x=171020000;
#10;x=171030000;
#10;x=171040000;
#10;x=171050000;
#10;x=171060000;
#10;x=171070000;
#10;x=171080000;
#10;x=171090000;
#10;x=171100000;
#10;x=171110000;
#10;x=171120000;
#10;x=171130000;
#10;x=171140000;
#10;x=171150000;
#10;x=171160000;
#10;x=171170000;
#10;x=171180000;
#10;x=171190000;
#10;x=171200000;
#10;x=171210000;
#10;x=171220000;
#10;x=171230000;
#10;x=171240000;
#10;x=171250000;
#10;x=171260000;
#10;x=171270000;
#10;x=171280000;
#10;x=171290000;
#10;x=171300000;
#10;x=171310000;
#10;x=171320000;
#10;x=171330000;
#10;x=171340000;
#10;x=171350000;
#10;x=171360000;
#10;x=171370000;
#10;x=171380000;
#10;x=171390000;
#10;x=171400000;
#10;x=171410000;
#10;x=171420000;
#10;x=171430000;
#10;x=171440000;
#10;x=171450000;
#10;x=171460000;
#10;x=171470000;
#10;x=171480000;
#10;x=171490000;
#10;x=171500000;
#10;x=171510000;
#10;x=171520000;
#10;x=171530000;
#10;x=171540000;
#10;x=171550000;
#10;x=171560000;
#10;x=171570000;
#10;x=171580000;
#10;x=171590000;
#10;x=171600000;
#10;x=171610000;
#10;x=171620000;
#10;x=171630000;
#10;x=171640000;
#10;x=171650000;
#10;x=171660000;
#10;x=171670000;
#10;x=171680000;
#10;x=171690000;
#10;x=171700000;
#10;x=171710000;
#10;x=171720000;
#10;x=171730000;
#10;x=171740000;
#10;x=171750000;
#10;x=171760000;
#10;x=171770000;
#10;x=171780000;
#10;x=171790000;
#10;x=171800000;
#10;x=171810000;
#10;x=171820000;
#10;x=171830000;
#10;x=171840000;
#10;x=171850000;
#10;x=171860000;
#10;x=171870000;
#10;x=171880000;
#10;x=171890000;
#10;x=171900000;
#10;x=171910000;
#10;x=171920000;
#10;x=171930000;
#10;x=171940000;
#10;x=171950000;
#10;x=171960000;
#10;x=171970000;
#10;x=171980000;
#10;x=171990000;
#10;x=172000000;
#10;x=172010000;
#10;x=172020000;
#10;x=172030000;
#10;x=172040000;
#10;x=172050000;
#10;x=172060000;
#10;x=172070000;
#10;x=172080000;
#10;x=172090000;
#10;x=172100000;
#10;x=172110000;
#10;x=172120000;
#10;x=172130000;
#10;x=172140000;
#10;x=172150000;
#10;x=172160000;
#10;x=172170000;
#10;x=172180000;
#10;x=172190000;
#10;x=172200000;
#10;x=172210000;
#10;x=172220000;
#10;x=172230000;
#10;x=172240000;
#10;x=172250000;
#10;x=172260000;
#10;x=172270000;
#10;x=172280000;
#10;x=172290000;
#10;x=172300000;
#10;x=172310000;
#10;x=172320000;
#10;x=172330000;
#10;x=172340000;
#10;x=172350000;
#10;x=172360000;
#10;x=172370000;
#10;x=172380000;
#10;x=172390000;
#10;x=172400000;
#10;x=172410000;
#10;x=172420000;
#10;x=172430000;
#10;x=172440000;
#10;x=172450000;
#10;x=172460000;
#10;x=172470000;
#10;x=172480000;
#10;x=172490000;
#10;x=172500000;
#10;x=172510000;
#10;x=172520000;
#10;x=172530000;
#10;x=172540000;
#10;x=172550000;
#10;x=172560000;
#10;x=172570000;
#10;x=172580000;
#10;x=172590000;
#10;x=172600000;
#10;x=172610000;
#10;x=172620000;
#10;x=172630000;
#10;x=172640000;
#10;x=172650000;
#10;x=172660000;
#10;x=172670000;
#10;x=172680000;
#10;x=172690000;
#10;x=172700000;
#10;x=172710000;
#10;x=172720000;
#10;x=172730000;
#10;x=172740000;
#10;x=172750000;
#10;x=172760000;
#10;x=172770000;
#10;x=172780000;
#10;x=172790000;
#10;x=172800000;
#10;x=172810000;
#10;x=172820000;
#10;x=172830000;
#10;x=172840000;
#10;x=172850000;
#10;x=172860000;
#10;x=172870000;
#10;x=172880000;
#10;x=172890000;
#10;x=172900000;
#10;x=172910000;
#10;x=172920000;
#10;x=172930000;
#10;x=172940000;
#10;x=172950000;
#10;x=172960000;
#10;x=172970000;
#10;x=172980000;
#10;x=172990000;
#10;x=173000000;
#10;x=173010000;
#10;x=173020000;
#10;x=173030000;
#10;x=173040000;
#10;x=173050000;
#10;x=173060000;
#10;x=173070000;
#10;x=173080000;
#10;x=173090000;
#10;x=173100000;
#10;x=173110000;
#10;x=173120000;
#10;x=173130000;
#10;x=173140000;
#10;x=173150000;
#10;x=173160000;
#10;x=173170000;
#10;x=173180000;
#10;x=173190000;
#10;x=173200000;
#10;x=173210000;
#10;x=173220000;
#10;x=173230000;
#10;x=173240000;
#10;x=173250000;
#10;x=173260000;
#10;x=173270000;
#10;x=173280000;
#10;x=173290000;
#10;x=173300000;
#10;x=173310000;
#10;x=173320000;
#10;x=173330000;
#10;x=173340000;
#10;x=173350000;
#10;x=173360000;
#10;x=173370000;
#10;x=173380000;
#10;x=173390000;
#10;x=173400000;
#10;x=173410000;
#10;x=173420000;
#10;x=173430000;
#10;x=173440000;
#10;x=173450000;
#10;x=173460000;
#10;x=173470000;
#10;x=173480000;
#10;x=173490000;
#10;x=173500000;
#10;x=173510000;
#10;x=173520000;
#10;x=173530000;
#10;x=173540000;
#10;x=173550000;
#10;x=173560000;
#10;x=173570000;
#10;x=173580000;
#10;x=173590000;
#10;x=173600000;
#10;x=173610000;
#10;x=173620000;
#10;x=173630000;
#10;x=173640000;
#10;x=173650000;
#10;x=173660000;
#10;x=173670000;
#10;x=173680000;
#10;x=173690000;
#10;x=173700000;
#10;x=173710000;
#10;x=173720000;
#10;x=173730000;
#10;x=173740000;
#10;x=173750000;
#10;x=173760000;
#10;x=173770000;
#10;x=173780000;
#10;x=173790000;
#10;x=173800000;
#10;x=173810000;
#10;x=173820000;
#10;x=173830000;
#10;x=173840000;
#10;x=173850000;
#10;x=173860000;
#10;x=173870000;
#10;x=173880000;
#10;x=173890000;
#10;x=173900000;
#10;x=173910000;
#10;x=173920000;
#10;x=173930000;
#10;x=173940000;
#10;x=173950000;
#10;x=173960000;
#10;x=173970000;
#10;x=173980000;
#10;x=173990000;
#10;x=174000000;
#10;x=174010000;
#10;x=174020000;
#10;x=174030000;
#10;x=174040000;
#10;x=174050000;
#10;x=174060000;
#10;x=174070000;
#10;x=174080000;
#10;x=174090000;
#10;x=174100000;
#10;x=174110000;
#10;x=174120000;
#10;x=174130000;
#10;x=174140000;
#10;x=174150000;
#10;x=174160000;
#10;x=174170000;
#10;x=174180000;
#10;x=174190000;
#10;x=174200000;
#10;x=174210000;
#10;x=174220000;
#10;x=174230000;
#10;x=174240000;
#10;x=174250000;
#10;x=174260000;
#10;x=174270000;
#10;x=174280000;
#10;x=174290000;
#10;x=174300000;
#10;x=174310000;
#10;x=174320000;
#10;x=174330000;
#10;x=174340000;
#10;x=174350000;
#10;x=174360000;
#10;x=174370000;
#10;x=174380000;
#10;x=174390000;
#10;x=174400000;
#10;x=174410000;
#10;x=174420000;
#10;x=174430000;
#10;x=174440000;
#10;x=174450000;
#10;x=174460000;
#10;x=174470000;
#10;x=174480000;
#10;x=174490000;
#10;x=174500000;
#10;x=174510000;
#10;x=174520000;
#10;x=174530000;
#10;x=174540000;
#10;x=174550000;
#10;x=174560000;
#10;x=174570000;
#10;x=174580000;
#10;x=174590000;
#10;x=174600000;
#10;x=174610000;
#10;x=174620000;
#10;x=174630000;
#10;x=174640000;
#10;x=174650000;
#10;x=174660000;
#10;x=174670000;
#10;x=174680000;
#10;x=174690000;
#10;x=174700000;
#10;x=174710000;
#10;x=174720000;
#10;x=174730000;
#10;x=174740000;
#10;x=174750000;
#10;x=174760000;
#10;x=174770000;
#10;x=174780000;
#10;x=174790000;
#10;x=174800000;
#10;x=174810000;
#10;x=174820000;
#10;x=174830000;
#10;x=174840000;
#10;x=174850000;
#10;x=174860000;
#10;x=174870000;
#10;x=174880000;
#10;x=174890000;
#10;x=174900000;
#10;x=174910000;
#10;x=174920000;
#10;x=174930000;
#10;x=174940000;
#10;x=174950000;
#10;x=174960000;
#10;x=174970000;
#10;x=174980000;
#10;x=174990000;
#10;x=175000000;
#10;x=175010000;
#10;x=175020000;
#10;x=175030000;
#10;x=175040000;
#10;x=175050000;
#10;x=175060000;
#10;x=175070000;
#10;x=175080000;
#10;x=175090000;
#10;x=175100000;
#10;x=175110000;
#10;x=175120000;
#10;x=175130000;
#10;x=175140000;
#10;x=175150000;
#10;x=175160000;
#10;x=175170000;
#10;x=175180000;
#10;x=175190000;
#10;x=175200000;
#10;x=175210000;
#10;x=175220000;
#10;x=175230000;
#10;x=175240000;
#10;x=175250000;
#10;x=175260000;
#10;x=175270000;
#10;x=175280000;
#10;x=175290000;
#10;x=175300000;
#10;x=175310000;
#10;x=175320000;
#10;x=175330000;
#10;x=175340000;
#10;x=175350000;
#10;x=175360000;
#10;x=175370000;
#10;x=175380000;
#10;x=175390000;
#10;x=175400000;
#10;x=175410000;
#10;x=175420000;
#10;x=175430000;
#10;x=175440000;
#10;x=175450000;
#10;x=175460000;
#10;x=175470000;
#10;x=175480000;
#10;x=175490000;
#10;x=175500000;
#10;x=175510000;
#10;x=175520000;
#10;x=175530000;
#10;x=175540000;
#10;x=175550000;
#10;x=175560000;
#10;x=175570000;
#10;x=175580000;
#10;x=175590000;
#10;x=175600000;
#10;x=175610000;
#10;x=175620000;
#10;x=175630000;
#10;x=175640000;
#10;x=175650000;
#10;x=175660000;
#10;x=175670000;
#10;x=175680000;
#10;x=175690000;
#10;x=175700000;
#10;x=175710000;
#10;x=175720000;
#10;x=175730000;
#10;x=175740000;
#10;x=175750000;
#10;x=175760000;
#10;x=175770000;
#10;x=175780000;
#10;x=175790000;
#10;x=175800000;
#10;x=175810000;
#10;x=175820000;
#10;x=175830000;
#10;x=175840000;
#10;x=175850000;
#10;x=175860000;
#10;x=175870000;
#10;x=175880000;
#10;x=175890000;
#10;x=175900000;
#10;x=175910000;
#10;x=175920000;
#10;x=175930000;
#10;x=175940000;
#10;x=175950000;
#10;x=175960000;
#10;x=175970000;
#10;x=175980000;
#10;x=175990000;
#10;x=176000000;
#10;x=176010000;
#10;x=176020000;
#10;x=176030000;
#10;x=176040000;
#10;x=176050000;
#10;x=176060000;
#10;x=176070000;
#10;x=176080000;
#10;x=176090000;
#10;x=176100000;
#10;x=176110000;
#10;x=176120000;
#10;x=176130000;
#10;x=176140000;
#10;x=176150000;
#10;x=176160000;
#10;x=176170000;
#10;x=176180000;
#10;x=176190000;
#10;x=176200000;
#10;x=176210000;
#10;x=176220000;
#10;x=176230000;
#10;x=176240000;
#10;x=176250000;
#10;x=176260000;
#10;x=176270000;
#10;x=176280000;
#10;x=176290000;
#10;x=176300000;
#10;x=176310000;
#10;x=176320000;
#10;x=176330000;
#10;x=176340000;
#10;x=176350000;
#10;x=176360000;
#10;x=176370000;
#10;x=176380000;
#10;x=176390000;
#10;x=176400000;
#10;x=176410000;
#10;x=176420000;
#10;x=176430000;
#10;x=176440000;
#10;x=176450000;
#10;x=176460000;
#10;x=176470000;
#10;x=176480000;
#10;x=176490000;
#10;x=176500000;
#10;x=176510000;
#10;x=176520000;
#10;x=176530000;
#10;x=176540000;
#10;x=176550000;
#10;x=176560000;
#10;x=176570000;
#10;x=176580000;
#10;x=176590000;
#10;x=176600000;
#10;x=176610000;
#10;x=176620000;
#10;x=176630000;
#10;x=176640000;
#10;x=176650000;
#10;x=176660000;
#10;x=176670000;
#10;x=176680000;
#10;x=176690000;
#10;x=176700000;
#10;x=176710000;
#10;x=176720000;
#10;x=176730000;
#10;x=176740000;
#10;x=176750000;
#10;x=176760000;
#10;x=176770000;
#10;x=176780000;
#10;x=176790000;
#10;x=176800000;
#10;x=176810000;
#10;x=176820000;
#10;x=176830000;
#10;x=176840000;
#10;x=176850000;
#10;x=176860000;
#10;x=176870000;
#10;x=176880000;
#10;x=176890000;
#10;x=176900000;
#10;x=176910000;
#10;x=176920000;
#10;x=176930000;
#10;x=176940000;
#10;x=176950000;
#10;x=176960000;
#10;x=176970000;
#10;x=176980000;
#10;x=176990000;
#10;x=177000000;
#10;x=177010000;
#10;x=177020000;
#10;x=177030000;
#10;x=177040000;
#10;x=177050000;
#10;x=177060000;
#10;x=177070000;
#10;x=177080000;
#10;x=177090000;
#10;x=177100000;
#10;x=177110000;
#10;x=177120000;
#10;x=177130000;
#10;x=177140000;
#10;x=177150000;
#10;x=177160000;
#10;x=177170000;
#10;x=177180000;
#10;x=177190000;
#10;x=177200000;
#10;x=177210000;
#10;x=177220000;
#10;x=177230000;
#10;x=177240000;
#10;x=177250000;
#10;x=177260000;
#10;x=177270000;
#10;x=177280000;
#10;x=177290000;
#10;x=177300000;
#10;x=177310000;
#10;x=177320000;
#10;x=177330000;
#10;x=177340000;
#10;x=177350000;
#10;x=177360000;
#10;x=177370000;
#10;x=177380000;
#10;x=177390000;
#10;x=177400000;
#10;x=177410000;
#10;x=177420000;
#10;x=177430000;
#10;x=177440000;
#10;x=177450000;
#10;x=177460000;
#10;x=177470000;
#10;x=177480000;
#10;x=177490000;
#10;x=177500000;
#10;x=177510000;
#10;x=177520000;
#10;x=177530000;
#10;x=177540000;
#10;x=177550000;
#10;x=177560000;
#10;x=177570000;
#10;x=177580000;
#10;x=177590000;
#10;x=177600000;
#10;x=177610000;
#10;x=177620000;
#10;x=177630000;
#10;x=177640000;
#10;x=177650000;
#10;x=177660000;
#10;x=177670000;
#10;x=177680000;
#10;x=177690000;
#10;x=177700000;
#10;x=177710000;
#10;x=177720000;
#10;x=177730000;
#10;x=177740000;
#10;x=177750000;
#10;x=177760000;
#10;x=177770000;
#10;x=177780000;
#10;x=177790000;
#10;x=177800000;
#10;x=177810000;
#10;x=177820000;
#10;x=177830000;
#10;x=177840000;
#10;x=177850000;
#10;x=177860000;
#10;x=177870000;
#10;x=177880000;
#10;x=177890000;
#10;x=177900000;
#10;x=177910000;
#10;x=177920000;
#10;x=177930000;
#10;x=177940000;
#10;x=177950000;
#10;x=177960000;
#10;x=177970000;
#10;x=177980000;
#10;x=177990000;
#10;x=178000000;
#10;x=178010000;
#10;x=178020000;
#10;x=178030000;
#10;x=178040000;
#10;x=178050000;
#10;x=178060000;
#10;x=178070000;
#10;x=178080000;
#10;x=178090000;
#10;x=178100000;
#10;x=178110000;
#10;x=178120000;
#10;x=178130000;
#10;x=178140000;
#10;x=178150000;
#10;x=178160000;
#10;x=178170000;
#10;x=178180000;
#10;x=178190000;
#10;x=178200000;
#10;x=178210000;
#10;x=178220000;
#10;x=178230000;
#10;x=178240000;
#10;x=178250000;
#10;x=178260000;
#10;x=178270000;
#10;x=178280000;
#10;x=178290000;
#10;x=178300000;
#10;x=178310000;
#10;x=178320000;
#10;x=178330000;
#10;x=178340000;
#10;x=178350000;
#10;x=178360000;
#10;x=178370000;
#10;x=178380000;
#10;x=178390000;
#10;x=178400000;
#10;x=178410000;
#10;x=178420000;
#10;x=178430000;
#10;x=178440000;
#10;x=178450000;
#10;x=178460000;
#10;x=178470000;
#10;x=178480000;
#10;x=178490000;
#10;x=178500000;
#10;x=178510000;
#10;x=178520000;
#10;x=178530000;
#10;x=178540000;
#10;x=178550000;
#10;x=178560000;
#10;x=178570000;
#10;x=178580000;
#10;x=178590000;
#10;x=178600000;
#10;x=178610000;
#10;x=178620000;
#10;x=178630000;
#10;x=178640000;
#10;x=178650000;
#10;x=178660000;
#10;x=178670000;
#10;x=178680000;
#10;x=178690000;
#10;x=178700000;
#10;x=178710000;
#10;x=178720000;
#10;x=178730000;
#10;x=178740000;
#10;x=178750000;
#10;x=178760000;
#10;x=178770000;
#10;x=178780000;
#10;x=178790000;
#10;x=178800000;
#10;x=178810000;
#10;x=178820000;
#10;x=178830000;
#10;x=178840000;
#10;x=178850000;
#10;x=178860000;
#10;x=178870000;
#10;x=178880000;
#10;x=178890000;
#10;x=178900000;
#10;x=178910000;
#10;x=178920000;
#10;x=178930000;
#10;x=178940000;
#10;x=178950000;
#10;x=178960000;
#10;x=178970000;
#10;x=178980000;
#10;x=178990000;
#10;x=179000000;
#10;x=179010000;
#10;x=179020000;
#10;x=179030000;
#10;x=179040000;
#10;x=179050000;
#10;x=179060000;
#10;x=179070000;
#10;x=179080000;
#10;x=179090000;
#10;x=179100000;
#10;x=179110000;
#10;x=179120000;
#10;x=179130000;
#10;x=179140000;
#10;x=179150000;
#10;x=179160000;
#10;x=179170000;
#10;x=179180000;
#10;x=179190000;
#10;x=179200000;
#10;x=179210000;
#10;x=179220000;
#10;x=179230000;
#10;x=179240000;
#10;x=179250000;
#10;x=179260000;
#10;x=179270000;
#10;x=179280000;
#10;x=179290000;
#10;x=179300000;
#10;x=179310000;
#10;x=179320000;
#10;x=179330000;
#10;x=179340000;
#10;x=179350000;
#10;x=179360000;
#10;x=179370000;
#10;x=179380000;
#10;x=179390000;
#10;x=179400000;
#10;x=179410000;
#10;x=179420000;
#10;x=179430000;
#10;x=179440000;
#10;x=179450000;
#10;x=179460000;
#10;x=179470000;
#10;x=179480000;
#10;x=179490000;
#10;x=179500000;
#10;x=179510000;
#10;x=179520000;
#10;x=179530000;
#10;x=179540000;
#10;x=179550000;
#10;x=179560000;
#10;x=179570000;
#10;x=179580000;
#10;x=179590000;
#10;x=179600000;
#10;x=179610000;
#10;x=179620000;
#10;x=179630000;
#10;x=179640000;
#10;x=179650000;
#10;x=179660000;
#10;x=179670000;
#10;x=179680000;
#10;x=179690000;
#10;x=179700000;
#10;x=179710000;
#10;x=179720000;
#10;x=179730000;
#10;x=179740000;
#10;x=179750000;
#10;x=179760000;
#10;x=179770000;
#10;x=179780000;
#10;x=179790000;
#10;x=179800000;
#10;x=179810000;
#10;x=179820000;
#10;x=179830000;
#10;x=179840000;
#10;x=179850000;
#10;x=179860000;
#10;x=179870000;
#10;x=179880000;
#10;x=179890000;
#10;x=179900000;
#10;x=179910000;
#10;x=179920000;
#10;x=179930000;
#10;x=179940000;
#10;x=179950000;
#10;x=179960000;
#10;x=179970000;
#10;x=179980000;
#10;x=179990000;
#10;x=180000000;
#10;x=180010000;
#10;x=180020000;
#10;x=180030000;
#10;x=180040000;
#10;x=180050000;
#10;x=180060000;
#10;x=180070000;
#10;x=180080000;
#10;x=180090000;
#10;x=180100000;
#10;x=180110000;
#10;x=180120000;
#10;x=180130000;
#10;x=180140000;
#10;x=180150000;
#10;x=180160000;
#10;x=180170000;
#10;x=180180000;
#10;x=180190000;
#10;x=180200000;
#10;x=180210000;
#10;x=180220000;
#10;x=180230000;
#10;x=180240000;
#10;x=180250000;
#10;x=180260000;
#10;x=180270000;
#10;x=180280000;
#10;x=180290000;
#10;x=180300000;
#10;x=180310000;
#10;x=180320000;
#10;x=180330000;
#10;x=180340000;
#10;x=180350000;
#10;x=180360000;
#10;x=180370000;
#10;x=180380000;
#10;x=180390000;
#10;x=180400000;
#10;x=180410000;
#10;x=180420000;
#10;x=180430000;
#10;x=180440000;
#10;x=180450000;
#10;x=180460000;
#10;x=180470000;
#10;x=180480000;
#10;x=180490000;
#10;x=180500000;
#10;x=180510000;
#10;x=180520000;
#10;x=180530000;
#10;x=180540000;
#10;x=180550000;
#10;x=180560000;
#10;x=180570000;
#10;x=180580000;
#10;x=180590000;
#10;x=180600000;
#10;x=180610000;
#10;x=180620000;
#10;x=180630000;
#10;x=180640000;
#10;x=180650000;
#10;x=180660000;
#10;x=180670000;
#10;x=180680000;
#10;x=180690000;
#10;x=180700000;
#10;x=180710000;
#10;x=180720000;
#10;x=180730000;
#10;x=180740000;
#10;x=180750000;
#10;x=180760000;
#10;x=180770000;
#10;x=180780000;
#10;x=180790000;
#10;x=180800000;
#10;x=180810000;
#10;x=180820000;
#10;x=180830000;
#10;x=180840000;
#10;x=180850000;
#10;x=180860000;
#10;x=180870000;
#10;x=180880000;
#10;x=180890000;
#10;x=180900000;
#10;x=180910000;
#10;x=180920000;
#10;x=180930000;
#10;x=180940000;
#10;x=180950000;
#10;x=180960000;
#10;x=180970000;
#10;x=180980000;
#10;x=180990000;
#10;x=181000000;
#10;x=181010000;
#10;x=181020000;
#10;x=181030000;
#10;x=181040000;
#10;x=181050000;
#10;x=181060000;
#10;x=181070000;
#10;x=181080000;
#10;x=181090000;
#10;x=181100000;
#10;x=181110000;
#10;x=181120000;
#10;x=181130000;
#10;x=181140000;
#10;x=181150000;
#10;x=181160000;
#10;x=181170000;
#10;x=181180000;
#10;x=181190000;
#10;x=181200000;
#10;x=181210000;
#10;x=181220000;
#10;x=181230000;
#10;x=181240000;
#10;x=181250000;
#10;x=181260000;
#10;x=181270000;
#10;x=181280000;
#10;x=181290000;
#10;x=181300000;
#10;x=181310000;
#10;x=181320000;
#10;x=181330000;
#10;x=181340000;
#10;x=181350000;
#10;x=181360000;
#10;x=181370000;
#10;x=181380000;
#10;x=181390000;
#10;x=181400000;
#10;x=181410000;
#10;x=181420000;
#10;x=181430000;
#10;x=181440000;
#10;x=181450000;
#10;x=181460000;
#10;x=181470000;
#10;x=181480000;
#10;x=181490000;
#10;x=181500000;
#10;x=181510000;
#10;x=181520000;
#10;x=181530000;
#10;x=181540000;
#10;x=181550000;
#10;x=181560000;
#10;x=181570000;
#10;x=181580000;
#10;x=181590000;
#10;x=181600000;
#10;x=181610000;
#10;x=181620000;
#10;x=181630000;
#10;x=181640000;
#10;x=181650000;
#10;x=181660000;
#10;x=181670000;
#10;x=181680000;
#10;x=181690000;
#10;x=181700000;
#10;x=181710000;
#10;x=181720000;
#10;x=181730000;
#10;x=181740000;
#10;x=181750000;
#10;x=181760000;
#10;x=181770000;
#10;x=181780000;
#10;x=181790000;
#10;x=181800000;
#10;x=181810000;
#10;x=181820000;
#10;x=181830000;
#10;x=181840000;
#10;x=181850000;
#10;x=181860000;
#10;x=181870000;
#10;x=181880000;
#10;x=181890000;
#10;x=181900000;
#10;x=181910000;
#10;x=181920000;
#10;x=181930000;
#10;x=181940000;
#10;x=181950000;
#10;x=181960000;
#10;x=181970000;
#10;x=181980000;
#10;x=181990000;
#10;x=182000000;
#10;x=182010000;
#10;x=182020000;
#10;x=182030000;
#10;x=182040000;
#10;x=182050000;
#10;x=182060000;
#10;x=182070000;
#10;x=182080000;
#10;x=182090000;
#10;x=182100000;
#10;x=182110000;
#10;x=182120000;
#10;x=182130000;
#10;x=182140000;
#10;x=182150000;
#10;x=182160000;
#10;x=182170000;
#10;x=182180000;
#10;x=182190000;
#10;x=182200000;
#10;x=182210000;
#10;x=182220000;
#10;x=182230000;
#10;x=182240000;
#10;x=182250000;
#10;x=182260000;
#10;x=182270000;
#10;x=182280000;
#10;x=182290000;
#10;x=182300000;
#10;x=182310000;
#10;x=182320000;
#10;x=182330000;
#10;x=182340000;
#10;x=182350000;
#10;x=182360000;
#10;x=182370000;
#10;x=182380000;
#10;x=182390000;
#10;x=182400000;
#10;x=182410000;
#10;x=182420000;
#10;x=182430000;
#10;x=182440000;
#10;x=182450000;
#10;x=182460000;
#10;x=182470000;
#10;x=182480000;
#10;x=182490000;
#10;x=182500000;
#10;x=182510000;
#10;x=182520000;
#10;x=182530000;
#10;x=182540000;
#10;x=182550000;
#10;x=182560000;
#10;x=182570000;
#10;x=182580000;
#10;x=182590000;
#10;x=182600000;
#10;x=182610000;
#10;x=182620000;
#10;x=182630000;
#10;x=182640000;
#10;x=182650000;
#10;x=182660000;
#10;x=182670000;
#10;x=182680000;
#10;x=182690000;
#10;x=182700000;
#10;x=182710000;
#10;x=182720000;
#10;x=182730000;
#10;x=182740000;
#10;x=182750000;
#10;x=182760000;
#10;x=182770000;
#10;x=182780000;
#10;x=182790000;
#10;x=182800000;
#10;x=182810000;
#10;x=182820000;
#10;x=182830000;
#10;x=182840000;
#10;x=182850000;
#10;x=182860000;
#10;x=182870000;
#10;x=182880000;
#10;x=182890000;
#10;x=182900000;
#10;x=182910000;
#10;x=182920000;
#10;x=182930000;
#10;x=182940000;
#10;x=182950000;
#10;x=182960000;
#10;x=182970000;
#10;x=182980000;
#10;x=182990000;
#10;x=183000000;
#10;x=183010000;
#10;x=183020000;
#10;x=183030000;
#10;x=183040000;
#10;x=183050000;
#10;x=183060000;
#10;x=183070000;
#10;x=183080000;
#10;x=183090000;
#10;x=183100000;
#10;x=183110000;
#10;x=183120000;
#10;x=183130000;
#10;x=183140000;
#10;x=183150000;
#10;x=183160000;
#10;x=183170000;
#10;x=183180000;
#10;x=183190000;
#10;x=183200000;
#10;x=183210000;
#10;x=183220000;
#10;x=183230000;
#10;x=183240000;
#10;x=183250000;
#10;x=183260000;
#10;x=183270000;
#10;x=183280000;
#10;x=183290000;
#10;x=183300000;
#10;x=183310000;
#10;x=183320000;
#10;x=183330000;
#10;x=183340000;
#10;x=183350000;
#10;x=183360000;
#10;x=183370000;
#10;x=183380000;
#10;x=183390000;
#10;x=183400000;
#10;x=183410000;
#10;x=183420000;
#10;x=183430000;
#10;x=183440000;
#10;x=183450000;
#10;x=183460000;
#10;x=183470000;
#10;x=183480000;
#10;x=183490000;
#10;x=183500000;
#10;x=183510000;
#10;x=183520000;
#10;x=183530000;
#10;x=183540000;
#10;x=183550000;
#10;x=183560000;
#10;x=183570000;
#10;x=183580000;
#10;x=183590000;
#10;x=183600000;
#10;x=183610000;
#10;x=183620000;
#10;x=183630000;
#10;x=183640000;
#10;x=183650000;
#10;x=183660000;
#10;x=183670000;
#10;x=183680000;
#10;x=183690000;
#10;x=183700000;
#10;x=183710000;
#10;x=183720000;
#10;x=183730000;
#10;x=183740000;
#10;x=183750000;
#10;x=183760000;
#10;x=183770000;
#10;x=183780000;
#10;x=183790000;
#10;x=183800000;
#10;x=183810000;
#10;x=183820000;
#10;x=183830000;
#10;x=183840000;
#10;x=183850000;
#10;x=183860000;
#10;x=183870000;
#10;x=183880000;
#10;x=183890000;
#10;x=183900000;
#10;x=183910000;
#10;x=183920000;
#10;x=183930000;
#10;x=183940000;
#10;x=183950000;
#10;x=183960000;
#10;x=183970000;
#10;x=183980000;
#10;x=183990000;
#10;x=184000000;
#10;x=184010000;
#10;x=184020000;
#10;x=184030000;
#10;x=184040000;
#10;x=184050000;
#10;x=184060000;
#10;x=184070000;
#10;x=184080000;
#10;x=184090000;
#10;x=184100000;
#10;x=184110000;
#10;x=184120000;
#10;x=184130000;
#10;x=184140000;
#10;x=184150000;
#10;x=184160000;
#10;x=184170000;
#10;x=184180000;
#10;x=184190000;
#10;x=184200000;
#10;x=184210000;
#10;x=184220000;
#10;x=184230000;
#10;x=184240000;
#10;x=184250000;
#10;x=184260000;
#10;x=184270000;
#10;x=184280000;
#10;x=184290000;
#10;x=184300000;
#10;x=184310000;
#10;x=184320000;
#10;x=184330000;
#10;x=184340000;
#10;x=184350000;
#10;x=184360000;
#10;x=184370000;
#10;x=184380000;
#10;x=184390000;
#10;x=184400000;
#10;x=184410000;
#10;x=184420000;
#10;x=184430000;
#10;x=184440000;
#10;x=184450000;
#10;x=184460000;
#10;x=184470000;
#10;x=184480000;
#10;x=184490000;
#10;x=184500000;
#10;x=184510000;
#10;x=184520000;
#10;x=184530000;
#10;x=184540000;
#10;x=184550000;
#10;x=184560000;
#10;x=184570000;
#10;x=184580000;
#10;x=184590000;
#10;x=184600000;
#10;x=184610000;
#10;x=184620000;
#10;x=184630000;
#10;x=184640000;
#10;x=184650000;
#10;x=184660000;
#10;x=184670000;
#10;x=184680000;
#10;x=184690000;
#10;x=184700000;
#10;x=184710000;
#10;x=184720000;
#10;x=184730000;
#10;x=184740000;
#10;x=184750000;
#10;x=184760000;
#10;x=184770000;
#10;x=184780000;
#10;x=184790000;
#10;x=184800000;
#10;x=184810000;
#10;x=184820000;
#10;x=184830000;
#10;x=184840000;
#10;x=184850000;
#10;x=184860000;
#10;x=184870000;
#10;x=184880000;
#10;x=184890000;
#10;x=184900000;
#10;x=184910000;
#10;x=184920000;
#10;x=184930000;
#10;x=184940000;
#10;x=184950000;
#10;x=184960000;
#10;x=184970000;
#10;x=184980000;
#10;x=184990000;
#10;x=185000000;
#10;x=185010000;
#10;x=185020000;
#10;x=185030000;
#10;x=185040000;
#10;x=185050000;
#10;x=185060000;
#10;x=185070000;
#10;x=185080000;
#10;x=185090000;
#10;x=185100000;
#10;x=185110000;
#10;x=185120000;
#10;x=185130000;
#10;x=185140000;
#10;x=185150000;
#10;x=185160000;
#10;x=185170000;
#10;x=185180000;
#10;x=185190000;
#10;x=185200000;
#10;x=185210000;
#10;x=185220000;
#10;x=185230000;
#10;x=185240000;
#10;x=185250000;
#10;x=185260000;
#10;x=185270000;
#10;x=185280000;
#10;x=185290000;
#10;x=185300000;
#10;x=185310000;
#10;x=185320000;
#10;x=185330000;
#10;x=185340000;
#10;x=185350000;
#10;x=185360000;
#10;x=185370000;
#10;x=185380000;
#10;x=185390000;
#10;x=185400000;
#10;x=185410000;
#10;x=185420000;
#10;x=185430000;
#10;x=185440000;
#10;x=185450000;
#10;x=185460000;
#10;x=185470000;
#10;x=185480000;
#10;x=185490000;
#10;x=185500000;
#10;x=185510000;
#10;x=185520000;
#10;x=185530000;
#10;x=185540000;
#10;x=185550000;
#10;x=185560000;
#10;x=185570000;
#10;x=185580000;
#10;x=185590000;
#10;x=185600000;
#10;x=185610000;
#10;x=185620000;
#10;x=185630000;
#10;x=185640000;
#10;x=185650000;
#10;x=185660000;
#10;x=185670000;
#10;x=185680000;
#10;x=185690000;
#10;x=185700000;
#10;x=185710000;
#10;x=185720000;
#10;x=185730000;
#10;x=185740000;
#10;x=185750000;
#10;x=185760000;
#10;x=185770000;
#10;x=185780000;
#10;x=185790000;
#10;x=185800000;
#10;x=185810000;
#10;x=185820000;
#10;x=185830000;
#10;x=185840000;
#10;x=185850000;
#10;x=185860000;
#10;x=185870000;
#10;x=185880000;
#10;x=185890000;
#10;x=185900000;
#10;x=185910000;
#10;x=185920000;
#10;x=185930000;
#10;x=185940000;
#10;x=185950000;
#10;x=185960000;
#10;x=185970000;
#10;x=185980000;
#10;x=185990000;
#10;x=186000000;
#10;x=186010000;
#10;x=186020000;
#10;x=186030000;
#10;x=186040000;
#10;x=186050000;
#10;x=186060000;
#10;x=186070000;
#10;x=186080000;
#10;x=186090000;
#10;x=186100000;
#10;x=186110000;
#10;x=186120000;
#10;x=186130000;
#10;x=186140000;
#10;x=186150000;
#10;x=186160000;
#10;x=186170000;
#10;x=186180000;
#10;x=186190000;
#10;x=186200000;
#10;x=186210000;
#10;x=186220000;
#10;x=186230000;
#10;x=186240000;
#10;x=186250000;
#10;x=186260000;
#10;x=186270000;
#10;x=186280000;
#10;x=186290000;
#10;x=186300000;
#10;x=186310000;
#10;x=186320000;
#10;x=186330000;
#10;x=186340000;
#10;x=186350000;
#10;x=186360000;
#10;x=186370000;
#10;x=186380000;
#10;x=186390000;
#10;x=186400000;
#10;x=186410000;
#10;x=186420000;
#10;x=186430000;
#10;x=186440000;
#10;x=186450000;
#10;x=186460000;
#10;x=186470000;
#10;x=186480000;
#10;x=186490000;
#10;x=186500000;
#10;x=186510000;
#10;x=186520000;
#10;x=186530000;
#10;x=186540000;
#10;x=186550000;
#10;x=186560000;
#10;x=186570000;
#10;x=186580000;
#10;x=186590000;
#10;x=186600000;
#10;x=186610000;
#10;x=186620000;
#10;x=186630000;
#10;x=186640000;
#10;x=186650000;
#10;x=186660000;
#10;x=186670000;
#10;x=186680000;
#10;x=186690000;
#10;x=186700000;
#10;x=186710000;
#10;x=186720000;
#10;x=186730000;
#10;x=186740000;
#10;x=186750000;
#10;x=186760000;
#10;x=186770000;
#10;x=186780000;
#10;x=186790000;
#10;x=186800000;
#10;x=186810000;
#10;x=186820000;
#10;x=186830000;
#10;x=186840000;
#10;x=186850000;
#10;x=186860000;
#10;x=186870000;
#10;x=186880000;
#10;x=186890000;
#10;x=186900000;
#10;x=186910000;
#10;x=186920000;
#10;x=186930000;
#10;x=186940000;
#10;x=186950000;
#10;x=186960000;
#10;x=186970000;
#10;x=186980000;
#10;x=186990000;
#10;x=187000000;
#10;x=187010000;
#10;x=187020000;
#10;x=187030000;
#10;x=187040000;
#10;x=187050000;
#10;x=187060000;
#10;x=187070000;
#10;x=187080000;
#10;x=187090000;
#10;x=187100000;
#10;x=187110000;
#10;x=187120000;
#10;x=187130000;
#10;x=187140000;
#10;x=187150000;
#10;x=187160000;
#10;x=187170000;
#10;x=187180000;
#10;x=187190000;
#10;x=187200000;
#10;x=187210000;
#10;x=187220000;
#10;x=187230000;
#10;x=187240000;
#10;x=187250000;
#10;x=187260000;
#10;x=187270000;
#10;x=187280000;
#10;x=187290000;
#10;x=187300000;
#10;x=187310000;
#10;x=187320000;
#10;x=187330000;
#10;x=187340000;
#10;x=187350000;
#10;x=187360000;
#10;x=187370000;
#10;x=187380000;
#10;x=187390000;
#10;x=187400000;
#10;x=187410000;
#10;x=187420000;
#10;x=187430000;
#10;x=187440000;
#10;x=187450000;
#10;x=187460000;
#10;x=187470000;
#10;x=187480000;
#10;x=187490000;
#10;x=187500000;
#10;x=187510000;
#10;x=187520000;
#10;x=187530000;
#10;x=187540000;
#10;x=187550000;
#10;x=187560000;
#10;x=187570000;
#10;x=187580000;
#10;x=187590000;
#10;x=187600000;
#10;x=187610000;
#10;x=187620000;
#10;x=187630000;
#10;x=187640000;
#10;x=187650000;
#10;x=187660000;
#10;x=187670000;
#10;x=187680000;
#10;x=187690000;
#10;x=187700000;
#10;x=187710000;
#10;x=187720000;
#10;x=187730000;
#10;x=187740000;
#10;x=187750000;
#10;x=187760000;
#10;x=187770000;
#10;x=187780000;
#10;x=187790000;
#10;x=187800000;
#10;x=187810000;
#10;x=187820000;
#10;x=187830000;
#10;x=187840000;
#10;x=187850000;
#10;x=187860000;
#10;x=187870000;
#10;x=187880000;
#10;x=187890000;
#10;x=187900000;
#10;x=187910000;
#10;x=187920000;
#10;x=187930000;
#10;x=187940000;
#10;x=187950000;
#10;x=187960000;
#10;x=187970000;
#10;x=187980000;
#10;x=187990000;
#10;x=188000000;
#10;x=188010000;
#10;x=188020000;
#10;x=188030000;
#10;x=188040000;
#10;x=188050000;
#10;x=188060000;
#10;x=188070000;
#10;x=188080000;
#10;x=188090000;
#10;x=188100000;
#10;x=188110000;
#10;x=188120000;
#10;x=188130000;
#10;x=188140000;
#10;x=188150000;
#10;x=188160000;
#10;x=188170000;
#10;x=188180000;
#10;x=188190000;
#10;x=188200000;
#10;x=188210000;
#10;x=188220000;
#10;x=188230000;
#10;x=188240000;
#10;x=188250000;
#10;x=188260000;
#10;x=188270000;
#10;x=188280000;
#10;x=188290000;
#10;x=188300000;
#10;x=188310000;
#10;x=188320000;
#10;x=188330000;
#10;x=188340000;
#10;x=188350000;
#10;x=188360000;
#10;x=188370000;
#10;x=188380000;
#10;x=188390000;
#10;x=188400000;
#10;x=188410000;
#10;x=188420000;
#10;x=188430000;
#10;x=188440000;
#10;x=188450000;
#10;x=188460000;
#10;x=188470000;
#10;x=188480000;
#10;x=188490000;
#10;x=188500000;
#10;x=188510000;
#10;x=188520000;
#10;x=188530000;
#10;x=188540000;
#10;x=188550000;
#10;x=188560000;
#10;x=188570000;
#10;x=188580000;
#10;x=188590000;
#10;x=188600000;
#10;x=188610000;
#10;x=188620000;
#10;x=188630000;
#10;x=188640000;
#10;x=188650000;
#10;x=188660000;
#10;x=188670000;
#10;x=188680000;
#10;x=188690000;
#10;x=188700000;
#10;x=188710000;
#10;x=188720000;
#10;x=188730000;
#10;x=188740000;
#10;x=188750000;
#10;x=188760000;
#10;x=188770000;
#10;x=188780000;
#10;x=188790000;
#10;x=188800000;
#10;x=188810000;
#10;x=188820000;
#10;x=188830000;
#10;x=188840000;
#10;x=188850000;
#10;x=188860000;
#10;x=188870000;
#10;x=188880000;
#10;x=188890000;
#10;x=188900000;
#10;x=188910000;
#10;x=188920000;
#10;x=188930000;
#10;x=188940000;
#10;x=188950000;
#10;x=188960000;
#10;x=188970000;
#10;x=188980000;
#10;x=188990000;
#10;x=189000000;
#10;x=189010000;
#10;x=189020000;
#10;x=189030000;
#10;x=189040000;
#10;x=189050000;
#10;x=189060000;
#10;x=189070000;
#10;x=189080000;
#10;x=189090000;
#10;x=189100000;
#10;x=189110000;
#10;x=189120000;
#10;x=189130000;
#10;x=189140000;
#10;x=189150000;
#10;x=189160000;
#10;x=189170000;
#10;x=189180000;
#10;x=189190000;
#10;x=189200000;
#10;x=189210000;
#10;x=189220000;
#10;x=189230000;
#10;x=189240000;
#10;x=189250000;
#10;x=189260000;
#10;x=189270000;
#10;x=189280000;
#10;x=189290000;
#10;x=189300000;
#10;x=189310000;
#10;x=189320000;
#10;x=189330000;
#10;x=189340000;
#10;x=189350000;
#10;x=189360000;
#10;x=189370000;
#10;x=189380000;
#10;x=189390000;
#10;x=189400000;
#10;x=189410000;
#10;x=189420000;
#10;x=189430000;
#10;x=189440000;
#10;x=189450000;
#10;x=189460000;
#10;x=189470000;
#10;x=189480000;
#10;x=189490000;
#10;x=189500000;
#10;x=189510000;
#10;x=189520000;
#10;x=189530000;
#10;x=189540000;
#10;x=189550000;
#10;x=189560000;
#10;x=189570000;
#10;x=189580000;
#10;x=189590000;
#10;x=189600000;
#10;x=189610000;
#10;x=189620000;
#10;x=189630000;
#10;x=189640000;
#10;x=189650000;
#10;x=189660000;
#10;x=189670000;
#10;x=189680000;
#10;x=189690000;
#10;x=189700000;
#10;x=189710000;
#10;x=189720000;
#10;x=189730000;
#10;x=189740000;
#10;x=189750000;
#10;x=189760000;
#10;x=189770000;
#10;x=189780000;
#10;x=189790000;
#10;x=189800000;
#10;x=189810000;
#10;x=189820000;
#10;x=189830000;
#10;x=189840000;
#10;x=189850000;
#10;x=189860000;
#10;x=189870000;
#10;x=189880000;
#10;x=189890000;
#10;x=189900000;
#10;x=189910000;
#10;x=189920000;
#10;x=189930000;
#10;x=189940000;
#10;x=189950000;
#10;x=189960000;
#10;x=189970000;
#10;x=189980000;
#10;x=189990000;
#10;x=190000000;
#10;x=190010000;
#10;x=190020000;
#10;x=190030000;
#10;x=190040000;
#10;x=190050000;
#10;x=190060000;
#10;x=190070000;
#10;x=190080000;
#10;x=190090000;
#10;x=190100000;
#10;x=190110000;
#10;x=190120000;
#10;x=190130000;
#10;x=190140000;
#10;x=190150000;
#10;x=190160000;
#10;x=190170000;
#10;x=190180000;
#10;x=190190000;
#10;x=190200000;
#10;x=190210000;
#10;x=190220000;
#10;x=190230000;
#10;x=190240000;
#10;x=190250000;
#10;x=190260000;
#10;x=190270000;
#10;x=190280000;
#10;x=190290000;
#10;x=190300000;
#10;x=190310000;
#10;x=190320000;
#10;x=190330000;
#10;x=190340000;
#10;x=190350000;
#10;x=190360000;
#10;x=190370000;
#10;x=190380000;
#10;x=190390000;
#10;x=190400000;
#10;x=190410000;
#10;x=190420000;
#10;x=190430000;
#10;x=190440000;
#10;x=190450000;
#10;x=190460000;
#10;x=190470000;
#10;x=190480000;
#10;x=190490000;
#10;x=190500000;
#10;x=190510000;
#10;x=190520000;
#10;x=190530000;
#10;x=190540000;
#10;x=190550000;
#10;x=190560000;
#10;x=190570000;
#10;x=190580000;
#10;x=190590000;
#10;x=190600000;
#10;x=190610000;
#10;x=190620000;
#10;x=190630000;
#10;x=190640000;
#10;x=190650000;
#10;x=190660000;
#10;x=190670000;
#10;x=190680000;
#10;x=190690000;
#10;x=190700000;
#10;x=190710000;
#10;x=190720000;
#10;x=190730000;
#10;x=190740000;
#10;x=190750000;
#10;x=190760000;
#10;x=190770000;
#10;x=190780000;
#10;x=190790000;
#10;x=190800000;
#10;x=190810000;
#10;x=190820000;
#10;x=190830000;
#10;x=190840000;
#10;x=190850000;
#10;x=190860000;
#10;x=190870000;
#10;x=190880000;
#10;x=190890000;
#10;x=190900000;
#10;x=190910000;
#10;x=190920000;
#10;x=190930000;
#10;x=190940000;
#10;x=190950000;
#10;x=190960000;
#10;x=190970000;
#10;x=190980000;
#10;x=190990000;
#10;x=191000000;
#10;x=191010000;
#10;x=191020000;
#10;x=191030000;
#10;x=191040000;
#10;x=191050000;
#10;x=191060000;
#10;x=191070000;
#10;x=191080000;
#10;x=191090000;
#10;x=191100000;
#10;x=191110000;
#10;x=191120000;
#10;x=191130000;
#10;x=191140000;
#10;x=191150000;
#10;x=191160000;
#10;x=191170000;
#10;x=191180000;
#10;x=191190000;
#10;x=191200000;
#10;x=191210000;
#10;x=191220000;
#10;x=191230000;
#10;x=191240000;
#10;x=191250000;
#10;x=191260000;
#10;x=191270000;
#10;x=191280000;
#10;x=191290000;
#10;x=191300000;
#10;x=191310000;
#10;x=191320000;
#10;x=191330000;
#10;x=191340000;
#10;x=191350000;
#10;x=191360000;
#10;x=191370000;
#10;x=191380000;
#10;x=191390000;
#10;x=191400000;
#10;x=191410000;
#10;x=191420000;
#10;x=191430000;
#10;x=191440000;
#10;x=191450000;
#10;x=191460000;
#10;x=191470000;
#10;x=191480000;
#10;x=191490000;
#10;x=191500000;
#10;x=191510000;
#10;x=191520000;
#10;x=191530000;
#10;x=191540000;
#10;x=191550000;
#10;x=191560000;
#10;x=191570000;
#10;x=191580000;
#10;x=191590000;
#10;x=191600000;
#10;x=191610000;
#10;x=191620000;
#10;x=191630000;
#10;x=191640000;
#10;x=191650000;
#10;x=191660000;
#10;x=191670000;
#10;x=191680000;
#10;x=191690000;
#10;x=191700000;
#10;x=191710000;
#10;x=191720000;
#10;x=191730000;
#10;x=191740000;
#10;x=191750000;
#10;x=191760000;
#10;x=191770000;
#10;x=191780000;
#10;x=191790000;
#10;x=191800000;
#10;x=191810000;
#10;x=191820000;
#10;x=191830000;
#10;x=191840000;
#10;x=191850000;
#10;x=191860000;
#10;x=191870000;
#10;x=191880000;
#10;x=191890000;
#10;x=191900000;
#10;x=191910000;
#10;x=191920000;
#10;x=191930000;
#10;x=191940000;
#10;x=191950000;
#10;x=191960000;
#10;x=191970000;
#10;x=191980000;
#10;x=191990000;
#10;x=192000000;
#10;x=192010000;
#10;x=192020000;
#10;x=192030000;
#10;x=192040000;
#10;x=192050000;
#10;x=192060000;
#10;x=192070000;
#10;x=192080000;
#10;x=192090000;
#10;x=192100000;
#10;x=192110000;
#10;x=192120000;
#10;x=192130000;
#10;x=192140000;
#10;x=192150000;
#10;x=192160000;
#10;x=192170000;
#10;x=192180000;
#10;x=192190000;
#10;x=192200000;
#10;x=192210000;
#10;x=192220000;
#10;x=192230000;
#10;x=192240000;
#10;x=192250000;
#10;x=192260000;
#10;x=192270000;
#10;x=192280000;
#10;x=192290000;
#10;x=192300000;
#10;x=192310000;
#10;x=192320000;
#10;x=192330000;
#10;x=192340000;
#10;x=192350000;
#10;x=192360000;
#10;x=192370000;
#10;x=192380000;
#10;x=192390000;
#10;x=192400000;
#10;x=192410000;
#10;x=192420000;
#10;x=192430000;
#10;x=192440000;
#10;x=192450000;
#10;x=192460000;
#10;x=192470000;
#10;x=192480000;
#10;x=192490000;
#10;x=192500000;
#10;x=192510000;
#10;x=192520000;
#10;x=192530000;
#10;x=192540000;
#10;x=192550000;
#10;x=192560000;
#10;x=192570000;
#10;x=192580000;
#10;x=192590000;
#10;x=192600000;
#10;x=192610000;
#10;x=192620000;
#10;x=192630000;
#10;x=192640000;
#10;x=192650000;
#10;x=192660000;
#10;x=192670000;
#10;x=192680000;
#10;x=192690000;
#10;x=192700000;
#10;x=192710000;
#10;x=192720000;
#10;x=192730000;
#10;x=192740000;
#10;x=192750000;
#10;x=192760000;
#10;x=192770000;
#10;x=192780000;
#10;x=192790000;
#10;x=192800000;
#10;x=192810000;
#10;x=192820000;
#10;x=192830000;
#10;x=192840000;
#10;x=192850000;
#10;x=192860000;
#10;x=192870000;
#10;x=192880000;
#10;x=192890000;
#10;x=192900000;
#10;x=192910000;
#10;x=192920000;
#10;x=192930000;
#10;x=192940000;
#10;x=192950000;
#10;x=192960000;
#10;x=192970000;
#10;x=192980000;
#10;x=192990000;
#10;x=193000000;
#10;x=193010000;
#10;x=193020000;
#10;x=193030000;
#10;x=193040000;
#10;x=193050000;
#10;x=193060000;
#10;x=193070000;
#10;x=193080000;
#10;x=193090000;
#10;x=193100000;
#10;x=193110000;
#10;x=193120000;
#10;x=193130000;
#10;x=193140000;
#10;x=193150000;
#10;x=193160000;
#10;x=193170000;
#10;x=193180000;
#10;x=193190000;
#10;x=193200000;
#10;x=193210000;
#10;x=193220000;
#10;x=193230000;
#10;x=193240000;
#10;x=193250000;
#10;x=193260000;
#10;x=193270000;
#10;x=193280000;
#10;x=193290000;
#10;x=193300000;
#10;x=193310000;
#10;x=193320000;
#10;x=193330000;
#10;x=193340000;
#10;x=193350000;
#10;x=193360000;
#10;x=193370000;
#10;x=193380000;
#10;x=193390000;
#10;x=193400000;
#10;x=193410000;
#10;x=193420000;
#10;x=193430000;
#10;x=193440000;
#10;x=193450000;
#10;x=193460000;
#10;x=193470000;
#10;x=193480000;
#10;x=193490000;
#10;x=193500000;
#10;x=193510000;
#10;x=193520000;
#10;x=193530000;
#10;x=193540000;
#10;x=193550000;
#10;x=193560000;
#10;x=193570000;
#10;x=193580000;
#10;x=193590000;
#10;x=193600000;
#10;x=193610000;
#10;x=193620000;
#10;x=193630000;
#10;x=193640000;
#10;x=193650000;
#10;x=193660000;
#10;x=193670000;
#10;x=193680000;
#10;x=193690000;
#10;x=193700000;
#10;x=193710000;
#10;x=193720000;
#10;x=193730000;
#10;x=193740000;
#10;x=193750000;
#10;x=193760000;
#10;x=193770000;
#10;x=193780000;
#10;x=193790000;
#10;x=193800000;
#10;x=193810000;
#10;x=193820000;
#10;x=193830000;
#10;x=193840000;
#10;x=193850000;
#10;x=193860000;
#10;x=193870000;
#10;x=193880000;
#10;x=193890000;
#10;x=193900000;
#10;x=193910000;
#10;x=193920000;
#10;x=193930000;
#10;x=193940000;
#10;x=193950000;
#10;x=193960000;
#10;x=193970000;
#10;x=193980000;
#10;x=193990000;
#10;x=194000000;
#10;x=194010000;
#10;x=194020000;
#10;x=194030000;
#10;x=194040000;
#10;x=194050000;
#10;x=194060000;
#10;x=194070000;
#10;x=194080000;
#10;x=194090000;
#10;x=194100000;
#10;x=194110000;
#10;x=194120000;
#10;x=194130000;
#10;x=194140000;
#10;x=194150000;
#10;x=194160000;
#10;x=194170000;
#10;x=194180000;
#10;x=194190000;
#10;x=194200000;
#10;x=194210000;
#10;x=194220000;
#10;x=194230000;
#10;x=194240000;
#10;x=194250000;
#10;x=194260000;
#10;x=194270000;
#10;x=194280000;
#10;x=194290000;
#10;x=194300000;
#10;x=194310000;
#10;x=194320000;
#10;x=194330000;
#10;x=194340000;
#10;x=194350000;
#10;x=194360000;
#10;x=194370000;
#10;x=194380000;
#10;x=194390000;
#10;x=194400000;
#10;x=194410000;
#10;x=194420000;
#10;x=194430000;
#10;x=194440000;
#10;x=194450000;
#10;x=194460000;
#10;x=194470000;
#10;x=194480000;
#10;x=194490000;
#10;x=194500000;
#10;x=194510000;
#10;x=194520000;
#10;x=194530000;
#10;x=194540000;
#10;x=194550000;
#10;x=194560000;
#10;x=194570000;
#10;x=194580000;
#10;x=194590000;
#10;x=194600000;
#10;x=194610000;
#10;x=194620000;
#10;x=194630000;
#10;x=194640000;
#10;x=194650000;
#10;x=194660000;
#10;x=194670000;
#10;x=194680000;
#10;x=194690000;
#10;x=194700000;
#10;x=194710000;
#10;x=194720000;
#10;x=194730000;
#10;x=194740000;
#10;x=194750000;
#10;x=194760000;
#10;x=194770000;
#10;x=194780000;
#10;x=194790000;
#10;x=194800000;
#10;x=194810000;
#10;x=194820000;
#10;x=194830000;
#10;x=194840000;
#10;x=194850000;
#10;x=194860000;
#10;x=194870000;
#10;x=194880000;
#10;x=194890000;
#10;x=194900000;
#10;x=194910000;
#10;x=194920000;
#10;x=194930000;
#10;x=194940000;
#10;x=194950000;
#10;x=194960000;
#10;x=194970000;
#10;x=194980000;
#10;x=194990000;
#10;x=195000000;
#10;x=195010000;
#10;x=195020000;
#10;x=195030000;
#10;x=195040000;
#10;x=195050000;
#10;x=195060000;
#10;x=195070000;
#10;x=195080000;
#10;x=195090000;
#10;x=195100000;
#10;x=195110000;
#10;x=195120000;
#10;x=195130000;
#10;x=195140000;
#10;x=195150000;
#10;x=195160000;
#10;x=195170000;
#10;x=195180000;
#10;x=195190000;
#10;x=195200000;
#10;x=195210000;
#10;x=195220000;
#10;x=195230000;
#10;x=195240000;
#10;x=195250000;
#10;x=195260000;
#10;x=195270000;
#10;x=195280000;
#10;x=195290000;
#10;x=195300000;
#10;x=195310000;
#10;x=195320000;
#10;x=195330000;
#10;x=195340000;
#10;x=195350000;
#10;x=195360000;
#10;x=195370000;
#10;x=195380000;
#10;x=195390000;
#10;x=195400000;
#10;x=195410000;
#10;x=195420000;
#10;x=195430000;
#10;x=195440000;
#10;x=195450000;
#10;x=195460000;
#10;x=195470000;
#10;x=195480000;
#10;x=195490000;
#10;x=195500000;
#10;x=195510000;
#10;x=195520000;
#10;x=195530000;
#10;x=195540000;
#10;x=195550000;
#10;x=195560000;
#10;x=195570000;
#10;x=195580000;
#10;x=195590000;
#10;x=195600000;
#10;x=195610000;
#10;x=195620000;
#10;x=195630000;
#10;x=195640000;
#10;x=195650000;
#10;x=195660000;
#10;x=195670000;
#10;x=195680000;
#10;x=195690000;
#10;x=195700000;
#10;x=195710000;
#10;x=195720000;
#10;x=195730000;
#10;x=195740000;
#10;x=195750000;
#10;x=195760000;
#10;x=195770000;
#10;x=195780000;
#10;x=195790000;
#10;x=195800000;
#10;x=195810000;
#10;x=195820000;
#10;x=195830000;
#10;x=195840000;
#10;x=195850000;
#10;x=195860000;
#10;x=195870000;
#10;x=195880000;
#10;x=195890000;
#10;x=195900000;
#10;x=195910000;
#10;x=195920000;
#10;x=195930000;
#10;x=195940000;
#10;x=195950000;
#10;x=195960000;
#10;x=195970000;
#10;x=195980000;
#10;x=195990000;
#10;x=196000000;
#10;x=196010000;
#10;x=196020000;
#10;x=196030000;
#10;x=196040000;
#10;x=196050000;
#10;x=196060000;
#10;x=196070000;
#10;x=196080000;
#10;x=196090000;
#10;x=196100000;
#10;x=196110000;
#10;x=196120000;
#10;x=196130000;
#10;x=196140000;
#10;x=196150000;
#10;x=196160000;
#10;x=196170000;
#10;x=196180000;
#10;x=196190000;
#10;x=196200000;
#10;x=196210000;
#10;x=196220000;
#10;x=196230000;
#10;x=196240000;
#10;x=196250000;
#10;x=196260000;
#10;x=196270000;
#10;x=196280000;
#10;x=196290000;
#10;x=196300000;
#10;x=196310000;
#10;x=196320000;
#10;x=196330000;
#10;x=196340000;
#10;x=196350000;
#10;x=196360000;
#10;x=196370000;
#10;x=196380000;
#10;x=196390000;
#10;x=196400000;
#10;x=196410000;
#10;x=196420000;
#10;x=196430000;
#10;x=196440000;
#10;x=196450000;
#10;x=196460000;
#10;x=196470000;
#10;x=196480000;
#10;x=196490000;
#10;x=196500000;
#10;x=196510000;
#10;x=196520000;
#10;x=196530000;
#10;x=196540000;
#10;x=196550000;
#10;x=196560000;
#10;x=196570000;
#10;x=196580000;
#10;x=196590000;
#10;x=196600000;
#10;x=196610000;
#10;x=196620000;
#10;x=196630000;
#10;x=196640000;
#10;x=196650000;
#10;x=196660000;
#10;x=196670000;
#10;x=196680000;
#10;x=196690000;
#10;x=196700000;
#10;x=196710000;
#10;x=196720000;
#10;x=196730000;
#10;x=196740000;
#10;x=196750000;
#10;x=196760000;
#10;x=196770000;
#10;x=196780000;
#10;x=196790000;
#10;x=196800000;
#10;x=196810000;
#10;x=196820000;
#10;x=196830000;
#10;x=196840000;
#10;x=196850000;
#10;x=196860000;
#10;x=196870000;
#10;x=196880000;
#10;x=196890000;
#10;x=196900000;
#10;x=196910000;
#10;x=196920000;
#10;x=196930000;
#10;x=196940000;
#10;x=196950000;
#10;x=196960000;
#10;x=196970000;
#10;x=196980000;
#10;x=196990000;
#10;x=197000000;
#10;x=197010000;
#10;x=197020000;
#10;x=197030000;
#10;x=197040000;
#10;x=197050000;
#10;x=197060000;
#10;x=197070000;
#10;x=197080000;
#10;x=197090000;
#10;x=197100000;
#10;x=197110000;
#10;x=197120000;
#10;x=197130000;
#10;x=197140000;
#10;x=197150000;
#10;x=197160000;
#10;x=197170000;
#10;x=197180000;
#10;x=197190000;
#10;x=197200000;
#10;x=197210000;
#10;x=197220000;
#10;x=197230000;
#10;x=197240000;
#10;x=197250000;
#10;x=197260000;
#10;x=197270000;
#10;x=197280000;
#10;x=197290000;
#10;x=197300000;
#10;x=197310000;
#10;x=197320000;
#10;x=197330000;
#10;x=197340000;
#10;x=197350000;
#10;x=197360000;
#10;x=197370000;
#10;x=197380000;
#10;x=197390000;
#10;x=197400000;
#10;x=197410000;
#10;x=197420000;
#10;x=197430000;
#10;x=197440000;
#10;x=197450000;
#10;x=197460000;
#10;x=197470000;
#10;x=197480000;
#10;x=197490000;
#10;x=197500000;
#10;x=197510000;
#10;x=197520000;
#10;x=197530000;
#10;x=197540000;
#10;x=197550000;
#10;x=197560000;
#10;x=197570000;
#10;x=197580000;
#10;x=197590000;
#10;x=197600000;
#10;x=197610000;
#10;x=197620000;
#10;x=197630000;
#10;x=197640000;
#10;x=197650000;
#10;x=197660000;
#10;x=197670000;
#10;x=197680000;
#10;x=197690000;
#10;x=197700000;
#10;x=197710000;
#10;x=197720000;
#10;x=197730000;
#10;x=197740000;
#10;x=197750000;
#10;x=197760000;
#10;x=197770000;
#10;x=197780000;
#10;x=197790000;
#10;x=197800000;
#10;x=197810000;
#10;x=197820000;
#10;x=197830000;
#10;x=197840000;
#10;x=197850000;
#10;x=197860000;
#10;x=197870000;
#10;x=197880000;
#10;x=197890000;
#10;x=197900000;
#10;x=197910000;
#10;x=197920000;
#10;x=197930000;
#10;x=197940000;
#10;x=197950000;
#10;x=197960000;
#10;x=197970000;
#10;x=197980000;
#10;x=197990000;
#10;x=198000000;
#10;x=198010000;
#10;x=198020000;
#10;x=198030000;
#10;x=198040000;
#10;x=198050000;
#10;x=198060000;
#10;x=198070000;
#10;x=198080000;
#10;x=198090000;
#10;x=198100000;
#10;x=198110000;
#10;x=198120000;
#10;x=198130000;
#10;x=198140000;
#10;x=198150000;
#10;x=198160000;
#10;x=198170000;
#10;x=198180000;
#10;x=198190000;
#10;x=198200000;
#10;x=198210000;
#10;x=198220000;
#10;x=198230000;
#10;x=198240000;
#10;x=198250000;
#10;x=198260000;
#10;x=198270000;
#10;x=198280000;
#10;x=198290000;
#10;x=198300000;
#10;x=198310000;
#10;x=198320000;
#10;x=198330000;
#10;x=198340000;
#10;x=198350000;
#10;x=198360000;
#10;x=198370000;
#10;x=198380000;
#10;x=198390000;
#10;x=198400000;
#10;x=198410000;
#10;x=198420000;
#10;x=198430000;
#10;x=198440000;
#10;x=198450000;
#10;x=198460000;
#10;x=198470000;
#10;x=198480000;
#10;x=198490000;
#10;x=198500000;
#10;x=198510000;
#10;x=198520000;
#10;x=198530000;
#10;x=198540000;
#10;x=198550000;
#10;x=198560000;
#10;x=198570000;
#10;x=198580000;
#10;x=198590000;
#10;x=198600000;
#10;x=198610000;
#10;x=198620000;
#10;x=198630000;
#10;x=198640000;
#10;x=198650000;
#10;x=198660000;
#10;x=198670000;
#10;x=198680000;
#10;x=198690000;
#10;x=198700000;
#10;x=198710000;
#10;x=198720000;
#10;x=198730000;
#10;x=198740000;
#10;x=198750000;
#10;x=198760000;
#10;x=198770000;
#10;x=198780000;
#10;x=198790000;
#10;x=198800000;
#10;x=198810000;
#10;x=198820000;
#10;x=198830000;
#10;x=198840000;
#10;x=198850000;
#10;x=198860000;
#10;x=198870000;
#10;x=198880000;
#10;x=198890000;
#10;x=198900000;
#10;x=198910000;
#10;x=198920000;
#10;x=198930000;
#10;x=198940000;
#10;x=198950000;
#10;x=198960000;
#10;x=198970000;
#10;x=198980000;
#10;x=198990000;
#10;x=199000000;
#10;x=199010000;
#10;x=199020000;
#10;x=199030000;
#10;x=199040000;
#10;x=199050000;
#10;x=199060000;
#10;x=199070000;
#10;x=199080000;
#10;x=199090000;
#10;x=199100000;
#10;x=199110000;
#10;x=199120000;
#10;x=199130000;
#10;x=199140000;
#10;x=199150000;
#10;x=199160000;
#10;x=199170000;
#10;x=199180000;
#10;x=199190000;
#10;x=199200000;
#10;x=199210000;
#10;x=199220000;
#10;x=199230000;
#10;x=199240000;
#10;x=199250000;
#10;x=199260000;
#10;x=199270000;
#10;x=199280000;
#10;x=199290000;
#10;x=199300000;
#10;x=199310000;
#10;x=199320000;
#10;x=199330000;
#10;x=199340000;
#10;x=199350000;
#10;x=199360000;
#10;x=199370000;
#10;x=199380000;
#10;x=199390000;
#10;x=199400000;
#10;x=199410000;
#10;x=199420000;
#10;x=199430000;
#10;x=199440000;
#10;x=199450000;
#10;x=199460000;
#10;x=199470000;
#10;x=199480000;
#10;x=199490000;
#10;x=199500000;
#10;x=199510000;
#10;x=199520000;
#10;x=199530000;
#10;x=199540000;
#10;x=199550000;
#10;x=199560000;
#10;x=199570000;
#10;x=199580000;
#10;x=199590000;
#10;x=199600000;
#10;x=199610000;
#10;x=199620000;
#10;x=199630000;
#10;x=199640000;
#10;x=199650000;
#10;x=199660000;
#10;x=199670000;
#10;x=199680000;
#10;x=199690000;
#10;x=199700000;
#10;x=199710000;
#10;x=199720000;
#10;x=199730000;
#10;x=199740000;
#10;x=199750000;
#10;x=199760000;
#10;x=199770000;
#10;x=199780000;
#10;x=199790000;
#10;x=199800000;
#10;x=199810000;
#10;x=199820000;
#10;x=199830000;
#10;x=199840000;
#10;x=199850000;
#10;x=199860000;
#10;x=199870000;
#10;x=199880000;
#10;x=199890000;
#10;x=199900000;
#10;x=199910000;
#10;x=199920000;
#10;x=199930000;
#10;x=199940000;
#10;x=199950000;
#10;x=199960000;
#10;x=199970000;
#10;x=199980000;
#10;x=199990000;
#10;x=200000000;
#10;x=200010000;
#10;x=200020000;
#10;x=200030000;
#10;x=200040000;
#10;x=200050000;
#10;x=200060000;
#10;x=200070000;
#10;x=200080000;
#10;x=200090000;
#10;x=200100000;
#10;x=200110000;
#10;x=200120000;
#10;x=200130000;
#10;x=200140000;
#10;x=200150000;
#10;x=200160000;
#10;x=200170000;
#10;x=200180000;
#10;x=200190000;
#10;x=200200000;
#10;x=200210000;
#10;x=200220000;
#10;x=200230000;
#10;x=200240000;
#10;x=200250000;
#10;x=200260000;
#10;x=200270000;
#10;x=200280000;
#10;x=200290000;
#10;x=200300000;
#10;x=200310000;
#10;x=200320000;
#10;x=200330000;
#10;x=200340000;
#10;x=200350000;
#10;x=200360000;
#10;x=200370000;
#10;x=200380000;
#10;x=200390000;
#10;x=200400000;
#10;x=200410000;
#10;x=200420000;
#10;x=200430000;
#10;x=200440000;
#10;x=200450000;
#10;x=200460000;
#10;x=200470000;
#10;x=200480000;
#10;x=200490000;
#10;x=200500000;
#10;x=200510000;
#10;x=200520000;
#10;x=200530000;
#10;x=200540000;
#10;x=200550000;
#10;x=200560000;
#10;x=200570000;
#10;x=200580000;
#10;x=200590000;
#10;x=200600000;
#10;x=200610000;
#10;x=200620000;
#10;x=200630000;
#10;x=200640000;
#10;x=200650000;
#10;x=200660000;
#10;x=200670000;
#10;x=200680000;
#10;x=200690000;
#10;x=200700000;
#10;x=200710000;
#10;x=200720000;
#10;x=200730000;
#10;x=200740000;
#10;x=200750000;
#10;x=200760000;
#10;x=200770000;
#10;x=200780000;
#10;x=200790000;
#10;x=200800000;
#10;x=200810000;
#10;x=200820000;
#10;x=200830000;
#10;x=200840000;
#10;x=200850000;
#10;x=200860000;
#10;x=200870000;
#10;x=200880000;
#10;x=200890000;
#10;x=200900000;
#10;x=200910000;
#10;x=200920000;
#10;x=200930000;
#10;x=200940000;
#10;x=200950000;
#10;x=200960000;
#10;x=200970000;
#10;x=200980000;
#10;x=200990000;
#10;x=201000000;
#10;x=201010000;
#10;x=201020000;
#10;x=201030000;
#10;x=201040000;
#10;x=201050000;
#10;x=201060000;
#10;x=201070000;
#10;x=201080000;
#10;x=201090000;
#10;x=201100000;
#10;x=201110000;
#10;x=201120000;
#10;x=201130000;
#10;x=201140000;
#10;x=201150000;
#10;x=201160000;
#10;x=201170000;
#10;x=201180000;
#10;x=201190000;
#10;x=201200000;
#10;x=201210000;
#10;x=201220000;
#10;x=201230000;
#10;x=201240000;
#10;x=201250000;
#10;x=201260000;
#10;x=201270000;
#10;x=201280000;
#10;x=201290000;
#10;x=201300000;
#10;x=201310000;
#10;x=201320000;
#10;x=201330000;
#10;x=201340000;
#10;x=201350000;
#10;x=201360000;
#10;x=201370000;
#10;x=201380000;
#10;x=201390000;
#10;x=201400000;
#10;x=201410000;
#10;x=201420000;
#10;x=201430000;
#10;x=201440000;
#10;x=201450000;
#10;x=201460000;
#10;x=201470000;
#10;x=201480000;
#10;x=201490000;
#10;x=201500000;
#10;x=201510000;
#10;x=201520000;
#10;x=201530000;
#10;x=201540000;
#10;x=201550000;
#10;x=201560000;
#10;x=201570000;
#10;x=201580000;
#10;x=201590000;
#10;x=201600000;
#10;x=201610000;
#10;x=201620000;
#10;x=201630000;
#10;x=201640000;
#10;x=201650000;
#10;x=201660000;
#10;x=201670000;
#10;x=201680000;
#10;x=201690000;
#10;x=201700000;
#10;x=201710000;
#10;x=201720000;
#10;x=201730000;
#10;x=201740000;
#10;x=201750000;
#10;x=201760000;
#10;x=201770000;
#10;x=201780000;
#10;x=201790000;
#10;x=201800000;
#10;x=201810000;
#10;x=201820000;
#10;x=201830000;
#10;x=201840000;
#10;x=201850000;
#10;x=201860000;
#10;x=201870000;
#10;x=201880000;
#10;x=201890000;
#10;x=201900000;
#10;x=201910000;
#10;x=201920000;
#10;x=201930000;
#10;x=201940000;
#10;x=201950000;
#10;x=201960000;
#10;x=201970000;
#10;x=201980000;
#10;x=201990000;
#10;x=202000000;
#10;x=202010000;
#10;x=202020000;
#10;x=202030000;
#10;x=202040000;
#10;x=202050000;
#10;x=202060000;
#10;x=202070000;
#10;x=202080000;
#10;x=202090000;
#10;x=202100000;
#10;x=202110000;
#10;x=202120000;
#10;x=202130000;
#10;x=202140000;
#10;x=202150000;
#10;x=202160000;
#10;x=202170000;
#10;x=202180000;
#10;x=202190000;
#10;x=202200000;
#10;x=202210000;
#10;x=202220000;
#10;x=202230000;
#10;x=202240000;
#10;x=202250000;
#10;x=202260000;
#10;x=202270000;
#10;x=202280000;
#10;x=202290000;
#10;x=202300000;
#10;x=202310000;
#10;x=202320000;
#10;x=202330000;
#10;x=202340000;
#10;x=202350000;
#10;x=202360000;
#10;x=202370000;
#10;x=202380000;
#10;x=202390000;
#10;x=202400000;
#10;x=202410000;
#10;x=202420000;
#10;x=202430000;
#10;x=202440000;
#10;x=202450000;
#10;x=202460000;
#10;x=202470000;
#10;x=202480000;
#10;x=202490000;
#10;x=202500000;
#10;x=202510000;
#10;x=202520000;
#10;x=202530000;
#10;x=202540000;
#10;x=202550000;
#10;x=202560000;
#10;x=202570000;
#10;x=202580000;
#10;x=202590000;
#10;x=202600000;
#10;x=202610000;
#10;x=202620000;
#10;x=202630000;
#10;x=202640000;
#10;x=202650000;
#10;x=202660000;
#10;x=202670000;
#10;x=202680000;
#10;x=202690000;
#10;x=202700000;
#10;x=202710000;
#10;x=202720000;
#10;x=202730000;
#10;x=202740000;
#10;x=202750000;
#10;x=202760000;
#10;x=202770000;
#10;x=202780000;
#10;x=202790000;
#10;x=202800000;
#10;x=202810000;
#10;x=202820000;
#10;x=202830000;
#10;x=202840000;
#10;x=202850000;
#10;x=202860000;
#10;x=202870000;
#10;x=202880000;
#10;x=202890000;
#10;x=202900000;
#10;x=202910000;
#10;x=202920000;
#10;x=202930000;
#10;x=202940000;
#10;x=202950000;
#10;x=202960000;
#10;x=202970000;
#10;x=202980000;
#10;x=202990000;
#10;x=203000000;
#10;x=203010000;
#10;x=203020000;
#10;x=203030000;
#10;x=203040000;
#10;x=203050000;
#10;x=203060000;
#10;x=203070000;
#10;x=203080000;
#10;x=203090000;
#10;x=203100000;
#10;x=203110000;
#10;x=203120000;
#10;x=203130000;
#10;x=203140000;
#10;x=203150000;
#10;x=203160000;
#10;x=203170000;
#10;x=203180000;
#10;x=203190000;
#10;x=203200000;
#10;x=203210000;
#10;x=203220000;
#10;x=203230000;
#10;x=203240000;
#10;x=203250000;
#10;x=203260000;
#10;x=203270000;
#10;x=203280000;
#10;x=203290000;
#10;x=203300000;
#10;x=203310000;
#10;x=203320000;
#10;x=203330000;
#10;x=203340000;
#10;x=203350000;
#10;x=203360000;
#10;x=203370000;
#10;x=203380000;
#10;x=203390000;
#10;x=203400000;
#10;x=203410000;
#10;x=203420000;
#10;x=203430000;
#10;x=203440000;
#10;x=203450000;
#10;x=203460000;
#10;x=203470000;
#10;x=203480000;
#10;x=203490000;
#10;x=203500000;
#10;x=203510000;
#10;x=203520000;
#10;x=203530000;
#10;x=203540000;
#10;x=203550000;
#10;x=203560000;
#10;x=203570000;
#10;x=203580000;
#10;x=203590000;
#10;x=203600000;
#10;x=203610000;
#10;x=203620000;
#10;x=203630000;
#10;x=203640000;
#10;x=203650000;
#10;x=203660000;
#10;x=203670000;
#10;x=203680000;
#10;x=203690000;
#10;x=203700000;
#10;x=203710000;
#10;x=203720000;
#10;x=203730000;
#10;x=203740000;
#10;x=203750000;
#10;x=203760000;
#10;x=203770000;
#10;x=203780000;
#10;x=203790000;
#10;x=203800000;
#10;x=203810000;
#10;x=203820000;
#10;x=203830000;
#10;x=203840000;
#10;x=203850000;
#10;x=203860000;
#10;x=203870000;
#10;x=203880000;
#10;x=203890000;
#10;x=203900000;
#10;x=203910000;
#10;x=203920000;
#10;x=203930000;
#10;x=203940000;
#10;x=203950000;
#10;x=203960000;
#10;x=203970000;
#10;x=203980000;
#10;x=203990000;
#10;x=204000000;
#10;x=204010000;
#10;x=204020000;
#10;x=204030000;
#10;x=204040000;
#10;x=204050000;
#10;x=204060000;
#10;x=204070000;
#10;x=204080000;
#10;x=204090000;
#10;x=204100000;
#10;x=204110000;
#10;x=204120000;
#10;x=204130000;
#10;x=204140000;
#10;x=204150000;
#10;x=204160000;
#10;x=204170000;
#10;x=204180000;
#10;x=204190000;
#10;x=204200000;
#10;x=204210000;
#10;x=204220000;
#10;x=204230000;
#10;x=204240000;
#10;x=204250000;
#10;x=204260000;
#10;x=204270000;
#10;x=204280000;
#10;x=204290000;
#10;x=204300000;
#10;x=204310000;
#10;x=204320000;
#10;x=204330000;
#10;x=204340000;
#10;x=204350000;
#10;x=204360000;
#10;x=204370000;
#10;x=204380000;
#10;x=204390000;
#10;x=204400000;
#10;x=204410000;
#10;x=204420000;
#10;x=204430000;
#10;x=204440000;
#10;x=204450000;
#10;x=204460000;
#10;x=204470000;
#10;x=204480000;
#10;x=204490000;
#10;x=204500000;
#10;x=204510000;
#10;x=204520000;
#10;x=204530000;
#10;x=204540000;
#10;x=204550000;
#10;x=204560000;
#10;x=204570000;
#10;x=204580000;
#10;x=204590000;
#10;x=204600000;
#10;x=204610000;
#10;x=204620000;
#10;x=204630000;
#10;x=204640000;
#10;x=204650000;
#10;x=204660000;
#10;x=204670000;
#10;x=204680000;
#10;x=204690000;
#10;x=204700000;
#10;x=204710000;
#10;x=204720000;
#10;x=204730000;
#10;x=204740000;
#10;x=204750000;
#10;x=204760000;
#10;x=204770000;
#10;x=204780000;
#10;x=204790000;
#10;x=204800000;
#10;x=204810000;
#10;x=204820000;
#10;x=204830000;
#10;x=204840000;
#10;x=204850000;
#10;x=204860000;
#10;x=204870000;
#10;x=204880000;
#10;x=204890000;
#10;x=204900000;
#10;x=204910000;
#10;x=204920000;
#10;x=204930000;
#10;x=204940000;
#10;x=204950000;
#10;x=204960000;
#10;x=204970000;
#10;x=204980000;
#10;x=204990000;
#10;x=205000000;
#10;x=205010000;
#10;x=205020000;
#10;x=205030000;
#10;x=205040000;
#10;x=205050000;
#10;x=205060000;
#10;x=205070000;
#10;x=205080000;
#10;x=205090000;
#10;x=205100000;
#10;x=205110000;
#10;x=205120000;
#10;x=205130000;
#10;x=205140000;
#10;x=205150000;
#10;x=205160000;
#10;x=205170000;
#10;x=205180000;
#10;x=205190000;
#10;x=205200000;
#10;x=205210000;
#10;x=205220000;
#10;x=205230000;
#10;x=205240000;
#10;x=205250000;
#10;x=205260000;
#10;x=205270000;
#10;x=205280000;
#10;x=205290000;
#10;x=205300000;
#10;x=205310000;
#10;x=205320000;
#10;x=205330000;
#10;x=205340000;
#10;x=205350000;
#10;x=205360000;
#10;x=205370000;
#10;x=205380000;
#10;x=205390000;
#10;x=205400000;
#10;x=205410000;
#10;x=205420000;
#10;x=205430000;
#10;x=205440000;
#10;x=205450000;
#10;x=205460000;
#10;x=205470000;
#10;x=205480000;
#10;x=205490000;
#10;x=205500000;
#10;x=205510000;
#10;x=205520000;
#10;x=205530000;
#10;x=205540000;
#10;x=205550000;
#10;x=205560000;
#10;x=205570000;
#10;x=205580000;
#10;x=205590000;
#10;x=205600000;
#10;x=205610000;
#10;x=205620000;
#10;x=205630000;
#10;x=205640000;
#10;x=205650000;
#10;x=205660000;
#10;x=205670000;
#10;x=205680000;
#10;x=205690000;
#10;x=205700000;
#10;x=205710000;
#10;x=205720000;
#10;x=205730000;
#10;x=205740000;
#10;x=205750000;
#10;x=205760000;
#10;x=205770000;
#10;x=205780000;
#10;x=205790000;
#10;x=205800000;
#10;x=205810000;
#10;x=205820000;
#10;x=205830000;
#10;x=205840000;
#10;x=205850000;
#10;x=205860000;
#10;x=205870000;
#10;x=205880000;
#10;x=205890000;
#10;x=205900000;
#10;x=205910000;
#10;x=205920000;
#10;x=205930000;
#10;x=205940000;
#10;x=205950000;
#10;x=205960000;
#10;x=205970000;
#10;x=205980000;
#10;x=205990000;
#10;x=206000000;
#10;x=206010000;
#10;x=206020000;
#10;x=206030000;
#10;x=206040000;
#10;x=206050000;
#10;x=206060000;
#10;x=206070000;
#10;x=206080000;
#10;x=206090000;
#10;x=206100000;
#10;x=206110000;
#10;x=206120000;
#10;x=206130000;
#10;x=206140000;
#10;x=206150000;
#10;x=206160000;
#10;x=206170000;
#10;x=206180000;
#10;x=206190000;
#10;x=206200000;
#10;x=206210000;
#10;x=206220000;
#10;x=206230000;
#10;x=206240000;
#10;x=206250000;
#10;x=206260000;
#10;x=206270000;
#10;x=206280000;
#10;x=206290000;
#10;x=206300000;
#10;x=206310000;
#10;x=206320000;
#10;x=206330000;
#10;x=206340000;
#10;x=206350000;
#10;x=206360000;
#10;x=206370000;
#10;x=206380000;
#10;x=206390000;
#10;x=206400000;
#10;x=206410000;
#10;x=206420000;
#10;x=206430000;
#10;x=206440000;
#10;x=206450000;
#10;x=206460000;
#10;x=206470000;
#10;x=206480000;
#10;x=206490000;
#10;x=206500000;
#10;x=206510000;
#10;x=206520000;
#10;x=206530000;
#10;x=206540000;
#10;x=206550000;
#10;x=206560000;
#10;x=206570000;
#10;x=206580000;
#10;x=206590000;
#10;x=206600000;
#10;x=206610000;
#10;x=206620000;
#10;x=206630000;
#10;x=206640000;
#10;x=206650000;
#10;x=206660000;
#10;x=206670000;
#10;x=206680000;
#10;x=206690000;
#10;x=206700000;
#10;x=206710000;
#10;x=206720000;
#10;x=206730000;
#10;x=206740000;
#10;x=206750000;
#10;x=206760000;
#10;x=206770000;
#10;x=206780000;
#10;x=206790000;
#10;x=206800000;
#10;x=206810000;
#10;x=206820000;
#10;x=206830000;
#10;x=206840000;
#10;x=206850000;
#10;x=206860000;
#10;x=206870000;
#10;x=206880000;
#10;x=206890000;
#10;x=206900000;
#10;x=206910000;
#10;x=206920000;
#10;x=206930000;
#10;x=206940000;
#10;x=206950000;
#10;x=206960000;
#10;x=206970000;
#10;x=206980000;
#10;x=206990000;
#10;x=207000000;
#10;x=207010000;
#10;x=207020000;
#10;x=207030000;
#10;x=207040000;
#10;x=207050000;
#10;x=207060000;
#10;x=207070000;
#10;x=207080000;
#10;x=207090000;
#10;x=207100000;
#10;x=207110000;
#10;x=207120000;
#10;x=207130000;
#10;x=207140000;
#10;x=207150000;
#10;x=207160000;
#10;x=207170000;
#10;x=207180000;
#10;x=207190000;
#10;x=207200000;
#10;x=207210000;
#10;x=207220000;
#10;x=207230000;
#10;x=207240000;
#10;x=207250000;
#10;x=207260000;
#10;x=207270000;
#10;x=207280000;
#10;x=207290000;
#10;x=207300000;
#10;x=207310000;
#10;x=207320000;
#10;x=207330000;
#10;x=207340000;
#10;x=207350000;
#10;x=207360000;
#10;x=207370000;
#10;x=207380000;
#10;x=207390000;
#10;x=207400000;
#10;x=207410000;
#10;x=207420000;
#10;x=207430000;
#10;x=207440000;
#10;x=207450000;
#10;x=207460000;
#10;x=207470000;
#10;x=207480000;
#10;x=207490000;
#10;x=207500000;
#10;x=207510000;
#10;x=207520000;
#10;x=207530000;
#10;x=207540000;
#10;x=207550000;
#10;x=207560000;
#10;x=207570000;
#10;x=207580000;
#10;x=207590000;
#10;x=207600000;
#10;x=207610000;
#10;x=207620000;
#10;x=207630000;
#10;x=207640000;
#10;x=207650000;
#10;x=207660000;
#10;x=207670000;
#10;x=207680000;
#10;x=207690000;
#10;x=207700000;
#10;x=207710000;
#10;x=207720000;
#10;x=207730000;
#10;x=207740000;
#10;x=207750000;
#10;x=207760000;
#10;x=207770000;
#10;x=207780000;
#10;x=207790000;
#10;x=207800000;
#10;x=207810000;
#10;x=207820000;
#10;x=207830000;
#10;x=207840000;
#10;x=207850000;
#10;x=207860000;
#10;x=207870000;
#10;x=207880000;
#10;x=207890000;
#10;x=207900000;
#10;x=207910000;
#10;x=207920000;
#10;x=207930000;
#10;x=207940000;
#10;x=207950000;
#10;x=207960000;
#10;x=207970000;
#10;x=207980000;
#10;x=207990000;
#10;x=208000000;
#10;x=208010000;
#10;x=208020000;
#10;x=208030000;
#10;x=208040000;
#10;x=208050000;
#10;x=208060000;
#10;x=208070000;
#10;x=208080000;
#10;x=208090000;
#10;x=208100000;
#10;x=208110000;
#10;x=208120000;
#10;x=208130000;
#10;x=208140000;
#10;x=208150000;
#10;x=208160000;
#10;x=208170000;
#10;x=208180000;
#10;x=208190000;
#10;x=208200000;
#10;x=208210000;
#10;x=208220000;
#10;x=208230000;
#10;x=208240000;
#10;x=208250000;
#10;x=208260000;
#10;x=208270000;
#10;x=208280000;
#10;x=208290000;
#10;x=208300000;
#10;x=208310000;
#10;x=208320000;
#10;x=208330000;
#10;x=208340000;
#10;x=208350000;
#10;x=208360000;
#10;x=208370000;
#10;x=208380000;
#10;x=208390000;
#10;x=208400000;
#10;x=208410000;
#10;x=208420000;
#10;x=208430000;
#10;x=208440000;
#10;x=208450000;
#10;x=208460000;
#10;x=208470000;
#10;x=208480000;
#10;x=208490000;
#10;x=208500000;
#10;x=208510000;
#10;x=208520000;
#10;x=208530000;
#10;x=208540000;
#10;x=208550000;
#10;x=208560000;
#10;x=208570000;
#10;x=208580000;
#10;x=208590000;
#10;x=208600000;
#10;x=208610000;
#10;x=208620000;
#10;x=208630000;
#10;x=208640000;
#10;x=208650000;
#10;x=208660000;
#10;x=208670000;
#10;x=208680000;
#10;x=208690000;
#10;x=208700000;
#10;x=208710000;
#10;x=208720000;
#10;x=208730000;
#10;x=208740000;
#10;x=208750000;
#10;x=208760000;
#10;x=208770000;
#10;x=208780000;
#10;x=208790000;
#10;x=208800000;
#10;x=208810000;
#10;x=208820000;
#10;x=208830000;
#10;x=208840000;
#10;x=208850000;
#10;x=208860000;
#10;x=208870000;
#10;x=208880000;
#10;x=208890000;
#10;x=208900000;
#10;x=208910000;
#10;x=208920000;
#10;x=208930000;
#10;x=208940000;
#10;x=208950000;
#10;x=208960000;
#10;x=208970000;
#10;x=208980000;
#10;x=208990000;
#10;x=209000000;
#10;x=209010000;
#10;x=209020000;
#10;x=209030000;
#10;x=209040000;
#10;x=209050000;
#10;x=209060000;
#10;x=209070000;
#10;x=209080000;
#10;x=209090000;
#10;x=209100000;
#10;x=209110000;
#10;x=209120000;
#10;x=209130000;
#10;x=209140000;
#10;x=209150000;
#10;x=209160000;
#10;x=209170000;
#10;x=209180000;
#10;x=209190000;
#10;x=209200000;
#10;x=209210000;
#10;x=209220000;
#10;x=209230000;
#10;x=209240000;
#10;x=209250000;
#10;x=209260000;
#10;x=209270000;
#10;x=209280000;
#10;x=209290000;
#10;x=209300000;
#10;x=209310000;
#10;x=209320000;
#10;x=209330000;
#10;x=209340000;
#10;x=209350000;
#10;x=209360000;
#10;x=209370000;
#10;x=209380000;
#10;x=209390000;
#10;x=209400000;
#10;x=209410000;
#10;x=209420000;
#10;x=209430000;
#10;x=209440000;
#10;x=209450000;
#10;x=209460000;
#10;x=209470000;
#10;x=209480000;
#10;x=209490000;
#10;x=209500000;
#10;x=209510000;
#10;x=209520000;
#10;x=209530000;
#10;x=209540000;
#10;x=209550000;
#10;x=209560000;
#10;x=209570000;
#10;x=209580000;
#10;x=209590000;
#10;x=209600000;
#10;x=209610000;
#10;x=209620000;
#10;x=209630000;
#10;x=209640000;
#10;x=209650000;
#10;x=209660000;
#10;x=209670000;
#10;x=209680000;
#10;x=209690000;
#10;x=209700000;
#10;x=209710000;
#10;x=209720000;
#10;x=209730000;
#10;x=209740000;
#10;x=209750000;
#10;x=209760000;
#10;x=209770000;
#10;x=209780000;
#10;x=209790000;
#10;x=209800000;
#10;x=209810000;
#10;x=209820000;
#10;x=209830000;
#10;x=209840000;
#10;x=209850000;
#10;x=209860000;
#10;x=209870000;
#10;x=209880000;
#10;x=209890000;
#10;x=209900000;
#10;x=209910000;
#10;x=209920000;
#10;x=209930000;
#10;x=209940000;
#10;x=209950000;
#10;x=209960000;
#10;x=209970000;
#10;x=209980000;
#10;x=209990000;
#10;x=210000000;
#10;x=210010000;
#10;x=210020000;
#10;x=210030000;
#10;x=210040000;
#10;x=210050000;
#10;x=210060000;
#10;x=210070000;
#10;x=210080000;
#10;x=210090000;
#10;x=210100000;
#10;x=210110000;
#10;x=210120000;
#10;x=210130000;
#10;x=210140000;
#10;x=210150000;
#10;x=210160000;
#10;x=210170000;
#10;x=210180000;
#10;x=210190000;
#10;x=210200000;
#10;x=210210000;
#10;x=210220000;
#10;x=210230000;
#10;x=210240000;
#10;x=210250000;
#10;x=210260000;
#10;x=210270000;
#10;x=210280000;
#10;x=210290000;
#10;x=210300000;
#10;x=210310000;
#10;x=210320000;
#10;x=210330000;
#10;x=210340000;
#10;x=210350000;
#10;x=210360000;
#10;x=210370000;
#10;x=210380000;
#10;x=210390000;
#10;x=210400000;
#10;x=210410000;
#10;x=210420000;
#10;x=210430000;
#10;x=210440000;
#10;x=210450000;
#10;x=210460000;
#10;x=210470000;
#10;x=210480000;
#10;x=210490000;
#10;x=210500000;
#10;x=210510000;
#10;x=210520000;
#10;x=210530000;
#10;x=210540000;
#10;x=210550000;
#10;x=210560000;
#10;x=210570000;
#10;x=210580000;
#10;x=210590000;
#10;x=210600000;
#10;x=210610000;
#10;x=210620000;
#10;x=210630000;
#10;x=210640000;
#10;x=210650000;
#10;x=210660000;
#10;x=210670000;
#10;x=210680000;
#10;x=210690000;
#10;x=210700000;
#10;x=210710000;
#10;x=210720000;
#10;x=210730000;
#10;x=210740000;
#10;x=210750000;
#10;x=210760000;
#10;x=210770000;
#10;x=210780000;
#10;x=210790000;
#10;x=210800000;
#10;x=210810000;
#10;x=210820000;
#10;x=210830000;
#10;x=210840000;
#10;x=210850000;
#10;x=210860000;
#10;x=210870000;
#10;x=210880000;
#10;x=210890000;
#10;x=210900000;
#10;x=210910000;
#10;x=210920000;
#10;x=210930000;
#10;x=210940000;
#10;x=210950000;
#10;x=210960000;
#10;x=210970000;
#10;x=210980000;
#10;x=210990000;
#10;x=211000000;
#10;x=211010000;
#10;x=211020000;
#10;x=211030000;
#10;x=211040000;
#10;x=211050000;
#10;x=211060000;
#10;x=211070000;
#10;x=211080000;
#10;x=211090000;
#10;x=211100000;
#10;x=211110000;
#10;x=211120000;
#10;x=211130000;
#10;x=211140000;
#10;x=211150000;
#10;x=211160000;
#10;x=211170000;
#10;x=211180000;
#10;x=211190000;
#10;x=211200000;
#10;x=211210000;
#10;x=211220000;
#10;x=211230000;
#10;x=211240000;
#10;x=211250000;
#10;x=211260000;
#10;x=211270000;
#10;x=211280000;
#10;x=211290000;
#10;x=211300000;
#10;x=211310000;
#10;x=211320000;
#10;x=211330000;
#10;x=211340000;
#10;x=211350000;
#10;x=211360000;
#10;x=211370000;
#10;x=211380000;
#10;x=211390000;
#10;x=211400000;
#10;x=211410000;
#10;x=211420000;
#10;x=211430000;
#10;x=211440000;
#10;x=211450000;
#10;x=211460000;
#10;x=211470000;
#10;x=211480000;
#10;x=211490000;
#10;x=211500000;
#10;x=211510000;
#10;x=211520000;
#10;x=211530000;
#10;x=211540000;
#10;x=211550000;
#10;x=211560000;
#10;x=211570000;
#10;x=211580000;
#10;x=211590000;
#10;x=211600000;
#10;x=211610000;
#10;x=211620000;
#10;x=211630000;
#10;x=211640000;
#10;x=211650000;
#10;x=211660000;
#10;x=211670000;
#10;x=211680000;
#10;x=211690000;
#10;x=211700000;
#10;x=211710000;
#10;x=211720000;
#10;x=211730000;
#10;x=211740000;
#10;x=211750000;
#10;x=211760000;
#10;x=211770000;
#10;x=211780000;
#10;x=211790000;
#10;x=211800000;
#10;x=211810000;
#10;x=211820000;
#10;x=211830000;
#10;x=211840000;
#10;x=211850000;
#10;x=211860000;
#10;x=211870000;
#10;x=211880000;
#10;x=211890000;
#10;x=211900000;
#10;x=211910000;
#10;x=211920000;
#10;x=211930000;
#10;x=211940000;
#10;x=211950000;
#10;x=211960000;
#10;x=211970000;
#10;x=211980000;
#10;x=211990000;
#10;x=212000000;
#10;x=212010000;
#10;x=212020000;
#10;x=212030000;
#10;x=212040000;
#10;x=212050000;
#10;x=212060000;
#10;x=212070000;
#10;x=212080000;
#10;x=212090000;
#10;x=212100000;
#10;x=212110000;
#10;x=212120000;
#10;x=212130000;
#10;x=212140000;
#10;x=212150000;
#10;x=212160000;
#10;x=212170000;
#10;x=212180000;
#10;x=212190000;
#10;x=212200000;
#10;x=212210000;
#10;x=212220000;
#10;x=212230000;
#10;x=212240000;
#10;x=212250000;
#10;x=212260000;
#10;x=212270000;
#10;x=212280000;
#10;x=212290000;
#10;x=212300000;
#10;x=212310000;
#10;x=212320000;
#10;x=212330000;
#10;x=212340000;
#10;x=212350000;
#10;x=212360000;
#10;x=212370000;
#10;x=212380000;
#10;x=212390000;
#10;x=212400000;
#10;x=212410000;
#10;x=212420000;
#10;x=212430000;
#10;x=212440000;
#10;x=212450000;
#10;x=212460000;
#10;x=212470000;
#10;x=212480000;
#10;x=212490000;
#10;x=212500000;
#10;x=212510000;
#10;x=212520000;
#10;x=212530000;
#10;x=212540000;
#10;x=212550000;
#10;x=212560000;
#10;x=212570000;
#10;x=212580000;
#10;x=212590000;
#10;x=212600000;
#10;x=212610000;
#10;x=212620000;
#10;x=212630000;
#10;x=212640000;
#10;x=212650000;
#10;x=212660000;
#10;x=212670000;
#10;x=212680000;
#10;x=212690000;
#10;x=212700000;
#10;x=212710000;
#10;x=212720000;
#10;x=212730000;
#10;x=212740000;
#10;x=212750000;
#10;x=212760000;
#10;x=212770000;
#10;x=212780000;
#10;x=212790000;
#10;x=212800000;
#10;x=212810000;
#10;x=212820000;
#10;x=212830000;
#10;x=212840000;
#10;x=212850000;
#10;x=212860000;
#10;x=212870000;
#10;x=212880000;
#10;x=212890000;
#10;x=212900000;
#10;x=212910000;
#10;x=212920000;
#10;x=212930000;
#10;x=212940000;
#10;x=212950000;
#10;x=212960000;
#10;x=212970000;
#10;x=212980000;
#10;x=212990000;
#10;x=213000000;
#10;x=213010000;
#10;x=213020000;
#10;x=213030000;
#10;x=213040000;
#10;x=213050000;
#10;x=213060000;
#10;x=213070000;
#10;x=213080000;
#10;x=213090000;
#10;x=213100000;
#10;x=213110000;
#10;x=213120000;
#10;x=213130000;
#10;x=213140000;
#10;x=213150000;
#10;x=213160000;
#10;x=213170000;
#10;x=213180000;
#10;x=213190000;
#10;x=213200000;
#10;x=213210000;
#10;x=213220000;
#10;x=213230000;
#10;x=213240000;
#10;x=213250000;
#10;x=213260000;
#10;x=213270000;
#10;x=213280000;
#10;x=213290000;
#10;x=213300000;
#10;x=213310000;
#10;x=213320000;
#10;x=213330000;
#10;x=213340000;
#10;x=213350000;
#10;x=213360000;
#10;x=213370000;
#10;x=213380000;
#10;x=213390000;
#10;x=213400000;
#10;x=213410000;
#10;x=213420000;
#10;x=213430000;
#10;x=213440000;
#10;x=213450000;
#10;x=213460000;
#10;x=213470000;
#10;x=213480000;
#10;x=213490000;
#10;x=213500000;
#10;x=213510000;
#10;x=213520000;
#10;x=213530000;
#10;x=213540000;
#10;x=213550000;
#10;x=213560000;
#10;x=213570000;
#10;x=213580000;
#10;x=213590000;
#10;x=213600000;
#10;x=213610000;
#10;x=213620000;
#10;x=213630000;
#10;x=213640000;
#10;x=213650000;
#10;x=213660000;
#10;x=213670000;
#10;x=213680000;
#10;x=213690000;
#10;x=213700000;
#10;x=213710000;
#10;x=213720000;
#10;x=213730000;
#10;x=213740000;
#10;x=213750000;
#10;x=213760000;
#10;x=213770000;
#10;x=213780000;
#10;x=213790000;
#10;x=213800000;
#10;x=213810000;
#10;x=213820000;
#10;x=213830000;
#10;x=213840000;
#10;x=213850000;
#10;x=213860000;
#10;x=213870000;
#10;x=213880000;
#10;x=213890000;
#10;x=213900000;
#10;x=213910000;
#10;x=213920000;
#10;x=213930000;
#10;x=213940000;
#10;x=213950000;
#10;x=213960000;
#10;x=213970000;
#10;x=213980000;
#10;x=213990000;
#10;x=214000000;
#10;x=214010000;
#10;x=214020000;
#10;x=214030000;
#10;x=214040000;
#10;x=214050000;
#10;x=214060000;
#10;x=214070000;
#10;x=214080000;
#10;x=214090000;
#10;x=214100000;
#10;x=214110000;
#10;x=214120000;
#10;x=214130000;
#10;x=214140000;
#10;x=214150000;
#10;x=214160000;
#10;x=214170000;
#10;x=214180000;
#10;x=214190000;
#10;x=214200000;
#10;x=214210000;
#10;x=214220000;
#10;x=214230000;
#10;x=214240000;
#10;x=214250000;
#10;x=214260000;
#10;x=214270000;
#10;x=214280000;
#10;x=214290000;
#10;x=214300000;
#10;x=214310000;
#10;x=214320000;
#10;x=214330000;
#10;x=214340000;
#10;x=214350000;
#10;x=214360000;
#10;x=214370000;
#10;x=214380000;
#10;x=214390000;
#10;x=214400000;
#10;x=214410000;
#10;x=214420000;
#10;x=214430000;
#10;x=214440000;
#10;x=214450000;
#10;x=214460000;
#10;x=214470000;
#10;x=214480000;
#10;x=214490000;
#10;x=214500000;
#10;x=214510000;
#10;x=214520000;
#10;x=214530000;
#10;x=214540000;
#10;x=214550000;
#10;x=214560000;
#10;x=214570000;
#10;x=214580000;
#10;x=214590000;
#10;x=214600000;
#10;x=214610000;
#10;x=214620000;
#10;x=214630000;
#10;x=214640000;
#10;x=214650000;
#10;x=214660000;
#10;x=214670000;
#10;x=214680000;
#10;x=214690000;
#10;x=214700000;
#10;x=214710000;
#10;x=214720000;
#10;x=214730000;
#10;x=214740000;
#10;x=214750000;
#10;x=214760000;
#10;x=214770000;
#10;x=214780000;
#10;x=214790000;
#10;x=214800000;
#10;x=214810000;
#10;x=214820000;
#10;x=214830000;
#10;x=214840000;
#10;x=214850000;
#10;x=214860000;
#10;x=214870000;
#10;x=214880000;
#10;x=214890000;
#10;x=214900000;
#10;x=214910000;
#10;x=214920000;
#10;x=214930000;
#10;x=214940000;
#10;x=214950000;
#10;x=214960000;
#10;x=214970000;
#10;x=214980000;
#10;x=214990000;
#10;x=215000000;
#10;x=215010000;
#10;x=215020000;
#10;x=215030000;
#10;x=215040000;
#10;x=215050000;
#10;x=215060000;
#10;x=215070000;
#10;x=215080000;
#10;x=215090000;
#10;x=215100000;
#10;x=215110000;
#10;x=215120000;
#10;x=215130000;
#10;x=215140000;
#10;x=215150000;
#10;x=215160000;
#10;x=215170000;
#10;x=215180000;
#10;x=215190000;
#10;x=215200000;
#10;x=215210000;
#10;x=215220000;
#10;x=215230000;
#10;x=215240000;
#10;x=215250000;
#10;x=215260000;
#10;x=215270000;
#10;x=215280000;
#10;x=215290000;
#10;x=215300000;
#10;x=215310000;
#10;x=215320000;
#10;x=215330000;
#10;x=215340000;
#10;x=215350000;
#10;x=215360000;
#10;x=215370000;
#10;x=215380000;
#10;x=215390000;
#10;x=215400000;
#10;x=215410000;
#10;x=215420000;
#10;x=215430000;
#10;x=215440000;
#10;x=215450000;
#10;x=215460000;
#10;x=215470000;
#10;x=215480000;
#10;x=215490000;
#10;x=215500000;
#10;x=215510000;
#10;x=215520000;
#10;x=215530000;
#10;x=215540000;
#10;x=215550000;
#10;x=215560000;
#10;x=215570000;
#10;x=215580000;
#10;x=215590000;
#10;x=215600000;
#10;x=215610000;
#10;x=215620000;
#10;x=215630000;
#10;x=215640000;
#10;x=215650000;
#10;x=215660000;
#10;x=215670000;
#10;x=215680000;
#10;x=215690000;
#10;x=215700000;
#10;x=215710000;
#10;x=215720000;
#10;x=215730000;
#10;x=215740000;
#10;x=215750000;
#10;x=215760000;
#10;x=215770000;
#10;x=215780000;
#10;x=215790000;
#10;x=215800000;
#10;x=215810000;
#10;x=215820000;
#10;x=215830000;
#10;x=215840000;
#10;x=215850000;
#10;x=215860000;
#10;x=215870000;
#10;x=215880000;
#10;x=215890000;
#10;x=215900000;
#10;x=215910000;
#10;x=215920000;
#10;x=215930000;
#10;x=215940000;
#10;x=215950000;
#10;x=215960000;
#10;x=215970000;
#10;x=215980000;
#10;x=215990000;
#10;x=216000000;
#10;x=216010000;
#10;x=216020000;
#10;x=216030000;
#10;x=216040000;
#10;x=216050000;
#10;x=216060000;
#10;x=216070000;
#10;x=216080000;
#10;x=216090000;
#10;x=216100000;
#10;x=216110000;
#10;x=216120000;
#10;x=216130000;
#10;x=216140000;
#10;x=216150000;
#10;x=216160000;
#10;x=216170000;
#10;x=216180000;
#10;x=216190000;
#10;x=216200000;
#10;x=216210000;
#10;x=216220000;
#10;x=216230000;
#10;x=216240000;
#10;x=216250000;
#10;x=216260000;
#10;x=216270000;
#10;x=216280000;
#10;x=216290000;
#10;x=216300000;
#10;x=216310000;
#10;x=216320000;
#10;x=216330000;
#10;x=216340000;
#10;x=216350000;
#10;x=216360000;
#10;x=216370000;
#10;x=216380000;
#10;x=216390000;
#10;x=216400000;
#10;x=216410000;
#10;x=216420000;
#10;x=216430000;
#10;x=216440000;
#10;x=216450000;
#10;x=216460000;
#10;x=216470000;
#10;x=216480000;
#10;x=216490000;
#10;x=216500000;
#10;x=216510000;
#10;x=216520000;
#10;x=216530000;
#10;x=216540000;
#10;x=216550000;
#10;x=216560000;
#10;x=216570000;
#10;x=216580000;
#10;x=216590000;
#10;x=216600000;
#10;x=216610000;
#10;x=216620000;
#10;x=216630000;
#10;x=216640000;
#10;x=216650000;
#10;x=216660000;
#10;x=216670000;
#10;x=216680000;
#10;x=216690000;
#10;x=216700000;
#10;x=216710000;
#10;x=216720000;
#10;x=216730000;
#10;x=216740000;
#10;x=216750000;
#10;x=216760000;
#10;x=216770000;
#10;x=216780000;
#10;x=216790000;
#10;x=216800000;
#10;x=216810000;
#10;x=216820000;
#10;x=216830000;
#10;x=216840000;
#10;x=216850000;
#10;x=216860000;
#10;x=216870000;
#10;x=216880000;
#10;x=216890000;
#10;x=216900000;
#10;x=216910000;
#10;x=216920000;
#10;x=216930000;
#10;x=216940000;
#10;x=216950000;
#10;x=216960000;
#10;x=216970000;
#10;x=216980000;
#10;x=216990000;
#10;x=217000000;
#10;x=217010000;
#10;x=217020000;
#10;x=217030000;
#10;x=217040000;
#10;x=217050000;
#10;x=217060000;
#10;x=217070000;
#10;x=217080000;
#10;x=217090000;
#10;x=217100000;
#10;x=217110000;
#10;x=217120000;
#10;x=217130000;
#10;x=217140000;
#10;x=217150000;
#10;x=217160000;
#10;x=217170000;
#10;x=217180000;
#10;x=217190000;
#10;x=217200000;
#10;x=217210000;
#10;x=217220000;
#10;x=217230000;
#10;x=217240000;
#10;x=217250000;
#10;x=217260000;
#10;x=217270000;
#10;x=217280000;
#10;x=217290000;
#10;x=217300000;
#10;x=217310000;
#10;x=217320000;
#10;x=217330000;
#10;x=217340000;
#10;x=217350000;
#10;x=217360000;
#10;x=217370000;
#10;x=217380000;
#10;x=217390000;
#10;x=217400000;
#10;x=217410000;
#10;x=217420000;
#10;x=217430000;
#10;x=217440000;
#10;x=217450000;
#10;x=217460000;
#10;x=217470000;
#10;x=217480000;
#10;x=217490000;
#10;x=217500000;
#10;x=217510000;
#10;x=217520000;
#10;x=217530000;
#10;x=217540000;
#10;x=217550000;
#10;x=217560000;
#10;x=217570000;
#10;x=217580000;
#10;x=217590000;
#10;x=217600000;
#10;x=217610000;
#10;x=217620000;
#10;x=217630000;
#10;x=217640000;
#10;x=217650000;
#10;x=217660000;
#10;x=217670000;
#10;x=217680000;
#10;x=217690000;
#10;x=217700000;
#10;x=217710000;
#10;x=217720000;
#10;x=217730000;
#10;x=217740000;
#10;x=217750000;
#10;x=217760000;
#10;x=217770000;
#10;x=217780000;
#10;x=217790000;
#10;x=217800000;
#10;x=217810000;
#10;x=217820000;
#10;x=217830000;
#10;x=217840000;
#10;x=217850000;
#10;x=217860000;
#10;x=217870000;
#10;x=217880000;
#10;x=217890000;
#10;x=217900000;
#10;x=217910000;
#10;x=217920000;
#10;x=217930000;
#10;x=217940000;
#10;x=217950000;
#10;x=217960000;
#10;x=217970000;
#10;x=217980000;
#10;x=217990000;
#10;x=218000000;
#10;x=218010000;
#10;x=218020000;
#10;x=218030000;
#10;x=218040000;
#10;x=218050000;
#10;x=218060000;
#10;x=218070000;
#10;x=218080000;
#10;x=218090000;
#10;x=218100000;
#10;x=218110000;
#10;x=218120000;
#10;x=218130000;
#10;x=218140000;
#10;x=218150000;
#10;x=218160000;
#10;x=218170000;
#10;x=218180000;
#10;x=218190000;
#10;x=218200000;
#10;x=218210000;
#10;x=218220000;
#10;x=218230000;
#10;x=218240000;
#10;x=218250000;
#10;x=218260000;
#10;x=218270000;
#10;x=218280000;
#10;x=218290000;
#10;x=218300000;
#10;x=218310000;
#10;x=218320000;
#10;x=218330000;
#10;x=218340000;
#10;x=218350000;
#10;x=218360000;
#10;x=218370000;
#10;x=218380000;
#10;x=218390000;
#10;x=218400000;
#10;x=218410000;
#10;x=218420000;
#10;x=218430000;
#10;x=218440000;
#10;x=218450000;
#10;x=218460000;
#10;x=218470000;
#10;x=218480000;
#10;x=218490000;
#10;x=218500000;
#10;x=218510000;
#10;x=218520000;
#10;x=218530000;
#10;x=218540000;
#10;x=218550000;
#10;x=218560000;
#10;x=218570000;
#10;x=218580000;
#10;x=218590000;
#10;x=218600000;
#10;x=218610000;
#10;x=218620000;
#10;x=218630000;
#10;x=218640000;
#10;x=218650000;
#10;x=218660000;
#10;x=218670000;
#10;x=218680000;
#10;x=218690000;
#10;x=218700000;
#10;x=218710000;
#10;x=218720000;
#10;x=218730000;
#10;x=218740000;
#10;x=218750000;
#10;x=218760000;
#10;x=218770000;
#10;x=218780000;
#10;x=218790000;
#10;x=218800000;
#10;x=218810000;
#10;x=218820000;
#10;x=218830000;
#10;x=218840000;
#10;x=218850000;
#10;x=218860000;
#10;x=218870000;
#10;x=218880000;
#10;x=218890000;
#10;x=218900000;
#10;x=218910000;
#10;x=218920000;
#10;x=218930000;
#10;x=218940000;
#10;x=218950000;
#10;x=218960000;
#10;x=218970000;
#10;x=218980000;
#10;x=218990000;
#10;x=219000000;
#10;x=219010000;
#10;x=219020000;
#10;x=219030000;
#10;x=219040000;
#10;x=219050000;
#10;x=219060000;
#10;x=219070000;
#10;x=219080000;
#10;x=219090000;
#10;x=219100000;
#10;x=219110000;
#10;x=219120000;
#10;x=219130000;
#10;x=219140000;
#10;x=219150000;
#10;x=219160000;
#10;x=219170000;
#10;x=219180000;
#10;x=219190000;
#10;x=219200000;
#10;x=219210000;
#10;x=219220000;
#10;x=219230000;
#10;x=219240000;
#10;x=219250000;
#10;x=219260000;
#10;x=219270000;
#10;x=219280000;
#10;x=219290000;
#10;x=219300000;
#10;x=219310000;
#10;x=219320000;
#10;x=219330000;
#10;x=219340000;
#10;x=219350000;
#10;x=219360000;
#10;x=219370000;
#10;x=219380000;
#10;x=219390000;
#10;x=219400000;
#10;x=219410000;
#10;x=219420000;
#10;x=219430000;
#10;x=219440000;
#10;x=219450000;
#10;x=219460000;
#10;x=219470000;
#10;x=219480000;
#10;x=219490000;
#10;x=219500000;
#10;x=219510000;
#10;x=219520000;
#10;x=219530000;
#10;x=219540000;
#10;x=219550000;
#10;x=219560000;
#10;x=219570000;
#10;x=219580000;
#10;x=219590000;
#10;x=219600000;
#10;x=219610000;
#10;x=219620000;
#10;x=219630000;
#10;x=219640000;
#10;x=219650000;
#10;x=219660000;
#10;x=219670000;
#10;x=219680000;
#10;x=219690000;
#10;x=219700000;
#10;x=219710000;
#10;x=219720000;
#10;x=219730000;
#10;x=219740000;
#10;x=219750000;
#10;x=219760000;
#10;x=219770000;
#10;x=219780000;
#10;x=219790000;
#10;x=219800000;
#10;x=219810000;
#10;x=219820000;
#10;x=219830000;
#10;x=219840000;
#10;x=219850000;
#10;x=219860000;
#10;x=219870000;
#10;x=219880000;
#10;x=219890000;
#10;x=219900000;
#10;x=219910000;
#10;x=219920000;
#10;x=219930000;
#10;x=219940000;
#10;x=219950000;
#10;x=219960000;
#10;x=219970000;
#10;x=219980000;
#10;x=219990000;
#10;x=220000000;
#10;x=220010000;
#10;x=220020000;
#10;x=220030000;
#10;x=220040000;
#10;x=220050000;
#10;x=220060000;
#10;x=220070000;
#10;x=220080000;
#10;x=220090000;
#10;x=220100000;
#10;x=220110000;
#10;x=220120000;
#10;x=220130000;
#10;x=220140000;
#10;x=220150000;
#10;x=220160000;
#10;x=220170000;
#10;x=220180000;
#10;x=220190000;
#10;x=220200000;
#10;x=220210000;
#10;x=220220000;
#10;x=220230000;
#10;x=220240000;
#10;x=220250000;
#10;x=220260000;
#10;x=220270000;
#10;x=220280000;
#10;x=220290000;
#10;x=220300000;
#10;x=220310000;
#10;x=220320000;
#10;x=220330000;
#10;x=220340000;
#10;x=220350000;
#10;x=220360000;
#10;x=220370000;
#10;x=220380000;
#10;x=220390000;
#10;x=220400000;
#10;x=220410000;
#10;x=220420000;
#10;x=220430000;
#10;x=220440000;
#10;x=220450000;
#10;x=220460000;
#10;x=220470000;
#10;x=220480000;
#10;x=220490000;
#10;x=220500000;
#10;x=220510000;
#10;x=220520000;
#10;x=220530000;
#10;x=220540000;
#10;x=220550000;
#10;x=220560000;
#10;x=220570000;
#10;x=220580000;
#10;x=220590000;
#10;x=220600000;
#10;x=220610000;
#10;x=220620000;
#10;x=220630000;
#10;x=220640000;
#10;x=220650000;
#10;x=220660000;
#10;x=220670000;
#10;x=220680000;
#10;x=220690000;
#10;x=220700000;
#10;x=220710000;
#10;x=220720000;
#10;x=220730000;
#10;x=220740000;
#10;x=220750000;
#10;x=220760000;
#10;x=220770000;
#10;x=220780000;
#10;x=220790000;
#10;x=220800000;
#10;x=220810000;
#10;x=220820000;
#10;x=220830000;
#10;x=220840000;
#10;x=220850000;
#10;x=220860000;
#10;x=220870000;
#10;x=220880000;
#10;x=220890000;
#10;x=220900000;
#10;x=220910000;
#10;x=220920000;
#10;x=220930000;
#10;x=220940000;
#10;x=220950000;
#10;x=220960000;
#10;x=220970000;
#10;x=220980000;
#10;x=220990000;
#10;x=221000000;
#10;x=221010000;
#10;x=221020000;
#10;x=221030000;
#10;x=221040000;
#10;x=221050000;
#10;x=221060000;
#10;x=221070000;
#10;x=221080000;
#10;x=221090000;
#10;x=221100000;
#10;x=221110000;
#10;x=221120000;
#10;x=221130000;
#10;x=221140000;
#10;x=221150000;
#10;x=221160000;
#10;x=221170000;
#10;x=221180000;
#10;x=221190000;
#10;x=221200000;
#10;x=221210000;
#10;x=221220000;
#10;x=221230000;
#10;x=221240000;
#10;x=221250000;
#10;x=221260000;
#10;x=221270000;
#10;x=221280000;
#10;x=221290000;
#10;x=221300000;
#10;x=221310000;
#10;x=221320000;
#10;x=221330000;
#10;x=221340000;
#10;x=221350000;
#10;x=221360000;
#10;x=221370000;
#10;x=221380000;
#10;x=221390000;
#10;x=221400000;
#10;x=221410000;
#10;x=221420000;
#10;x=221430000;
#10;x=221440000;
#10;x=221450000;
#10;x=221460000;
#10;x=221470000;
#10;x=221480000;
#10;x=221490000;
#10;x=221500000;
#10;x=221510000;
#10;x=221520000;
#10;x=221530000;
#10;x=221540000;
#10;x=221550000;
#10;x=221560000;
#10;x=221570000;
#10;x=221580000;
#10;x=221590000;
#10;x=221600000;
#10;x=221610000;
#10;x=221620000;
#10;x=221630000;
#10;x=221640000;
#10;x=221650000;
#10;x=221660000;
#10;x=221670000;
#10;x=221680000;
#10;x=221690000;
#10;x=221700000;
#10;x=221710000;
#10;x=221720000;
#10;x=221730000;
#10;x=221740000;
#10;x=221750000;
#10;x=221760000;
#10;x=221770000;
#10;x=221780000;
#10;x=221790000;
#10;x=221800000;
#10;x=221810000;
#10;x=221820000;
#10;x=221830000;
#10;x=221840000;
#10;x=221850000;
#10;x=221860000;
#10;x=221870000;
#10;x=221880000;
#10;x=221890000;
#10;x=221900000;
#10;x=221910000;
#10;x=221920000;
#10;x=221930000;
#10;x=221940000;
#10;x=221950000;
#10;x=221960000;
#10;x=221970000;
#10;x=221980000;
#10;x=221990000;
#10;x=222000000;
#10;x=222010000;
#10;x=222020000;
#10;x=222030000;
#10;x=222040000;
#10;x=222050000;
#10;x=222060000;
#10;x=222070000;
#10;x=222080000;
#10;x=222090000;
#10;x=222100000;
#10;x=222110000;
#10;x=222120000;
#10;x=222130000;
#10;x=222140000;
#10;x=222150000;
#10;x=222160000;
#10;x=222170000;
#10;x=222180000;
#10;x=222190000;
#10;x=222200000;
#10;x=222210000;
#10;x=222220000;
#10;x=222230000;
#10;x=222240000;
#10;x=222250000;
#10;x=222260000;
#10;x=222270000;
#10;x=222280000;
#10;x=222290000;
#10;x=222300000;
#10;x=222310000;
#10;x=222320000;
#10;x=222330000;
#10;x=222340000;
#10;x=222350000;
#10;x=222360000;
#10;x=222370000;
#10;x=222380000;
#10;x=222390000;
#10;x=222400000;
#10;x=222410000;
#10;x=222420000;
#10;x=222430000;
#10;x=222440000;
#10;x=222450000;
#10;x=222460000;
#10;x=222470000;
#10;x=222480000;
#10;x=222490000;
#10;x=222500000;
#10;x=222510000;
#10;x=222520000;
#10;x=222530000;
#10;x=222540000;
#10;x=222550000;
#10;x=222560000;
#10;x=222570000;
#10;x=222580000;
#10;x=222590000;
#10;x=222600000;
#10;x=222610000;
#10;x=222620000;
#10;x=222630000;
#10;x=222640000;
#10;x=222650000;
#10;x=222660000;
#10;x=222670000;
#10;x=222680000;
#10;x=222690000;
#10;x=222700000;
#10;x=222710000;
#10;x=222720000;
#10;x=222730000;
#10;x=222740000;
#10;x=222750000;
#10;x=222760000;
#10;x=222770000;
#10;x=222780000;
#10;x=222790000;
#10;x=222800000;
#10;x=222810000;
#10;x=222820000;
#10;x=222830000;
#10;x=222840000;
#10;x=222850000;
#10;x=222860000;
#10;x=222870000;
#10;x=222880000;
#10;x=222890000;
#10;x=222900000;
#10;x=222910000;
#10;x=222920000;
#10;x=222930000;
#10;x=222940000;
#10;x=222950000;
#10;x=222960000;
#10;x=222970000;
#10;x=222980000;
#10;x=222990000;
#10;x=223000000;
#10;x=223010000;
#10;x=223020000;
#10;x=223030000;
#10;x=223040000;
#10;x=223050000;
#10;x=223060000;
#10;x=223070000;
#10;x=223080000;
#10;x=223090000;
#10;x=223100000;
#10;x=223110000;
#10;x=223120000;
#10;x=223130000;
#10;x=223140000;
#10;x=223150000;
#10;x=223160000;
#10;x=223170000;
#10;x=223180000;
#10;x=223190000;
#10;x=223200000;
#10;x=223210000;
#10;x=223220000;
#10;x=223230000;
#10;x=223240000;
#10;x=223250000;
#10;x=223260000;
#10;x=223270000;
#10;x=223280000;
#10;x=223290000;
#10;x=223300000;
#10;x=223310000;
#10;x=223320000;
#10;x=223330000;
#10;x=223340000;
#10;x=223350000;
#10;x=223360000;
#10;x=223370000;
#10;x=223380000;
#10;x=223390000;
#10;x=223400000;
#10;x=223410000;
#10;x=223420000;
#10;x=223430000;
#10;x=223440000;
#10;x=223450000;
#10;x=223460000;
#10;x=223470000;
#10;x=223480000;
#10;x=223490000;
#10;x=223500000;
#10;x=223510000;
#10;x=223520000;
#10;x=223530000;
#10;x=223540000;
#10;x=223550000;
#10;x=223560000;
#10;x=223570000;
#10;x=223580000;
#10;x=223590000;
#10;x=223600000;
#10;x=223610000;
#10;x=223620000;
#10;x=223630000;
#10;x=223640000;
#10;x=223650000;
#10;x=223660000;
#10;x=223670000;
#10;x=223680000;
#10;x=223690000;
#10;x=223700000;
#10;x=223710000;
#10;x=223720000;
#10;x=223730000;
#10;x=223740000;
#10;x=223750000;
#10;x=223760000;
#10;x=223770000;
#10;x=223780000;
#10;x=223790000;
#10;x=223800000;
#10;x=223810000;
#10;x=223820000;
#10;x=223830000;
#10;x=223840000;
#10;x=223850000;
#10;x=223860000;
#10;x=223870000;
#10;x=223880000;
#10;x=223890000;
#10;x=223900000;
#10;x=223910000;
#10;x=223920000;
#10;x=223930000;
#10;x=223940000;
#10;x=223950000;
#10;x=223960000;
#10;x=223970000;
#10;x=223980000;
#10;x=223990000;
#10;x=224000000;
#10;x=224010000;
#10;x=224020000;
#10;x=224030000;
#10;x=224040000;
#10;x=224050000;
#10;x=224060000;
#10;x=224070000;
#10;x=224080000;
#10;x=224090000;
#10;x=224100000;
#10;x=224110000;
#10;x=224120000;
#10;x=224130000;
#10;x=224140000;
#10;x=224150000;
#10;x=224160000;
#10;x=224170000;
#10;x=224180000;
#10;x=224190000;
#10;x=224200000;
#10;x=224210000;
#10;x=224220000;
#10;x=224230000;
#10;x=224240000;
#10;x=224250000;
#10;x=224260000;
#10;x=224270000;
#10;x=224280000;
#10;x=224290000;
#10;x=224300000;
#10;x=224310000;
#10;x=224320000;
#10;x=224330000;
#10;x=224340000;
#10;x=224350000;
#10;x=224360000;
#10;x=224370000;
#10;x=224380000;
#10;x=224390000;
#10;x=224400000;
#10;x=224410000;
#10;x=224420000;
#10;x=224430000;
#10;x=224440000;
#10;x=224450000;
#10;x=224460000;
#10;x=224470000;
#10;x=224480000;
#10;x=224490000;
#10;x=224500000;
#10;x=224510000;
#10;x=224520000;
#10;x=224530000;
#10;x=224540000;
#10;x=224550000;
#10;x=224560000;
#10;x=224570000;
#10;x=224580000;
#10;x=224590000;
#10;x=224600000;
#10;x=224610000;
#10;x=224620000;
#10;x=224630000;
#10;x=224640000;
#10;x=224650000;
#10;x=224660000;
#10;x=224670000;
#10;x=224680000;
#10;x=224690000;
#10;x=224700000;
#10;x=224710000;
#10;x=224720000;
#10;x=224730000;
#10;x=224740000;
#10;x=224750000;
#10;x=224760000;
#10;x=224770000;
#10;x=224780000;
#10;x=224790000;
#10;x=224800000;
#10;x=224810000;
#10;x=224820000;
#10;x=224830000;
#10;x=224840000;
#10;x=224850000;
#10;x=224860000;
#10;x=224870000;
#10;x=224880000;
#10;x=224890000;
#10;x=224900000;
#10;x=224910000;
#10;x=224920000;
#10;x=224930000;
#10;x=224940000;
#10;x=224950000;
#10;x=224960000;
#10;x=224970000;
#10;x=224980000;
#10;x=224990000;
#10;x=225000000;
#10;x=225010000;
#10;x=225020000;
#10;x=225030000;
#10;x=225040000;
#10;x=225050000;
#10;x=225060000;
#10;x=225070000;
#10;x=225080000;
#10;x=225090000;
#10;x=225100000;
#10;x=225110000;
#10;x=225120000;
#10;x=225130000;
#10;x=225140000;
#10;x=225150000;
#10;x=225160000;
#10;x=225170000;
#10;x=225180000;
#10;x=225190000;
#10;x=225200000;
#10;x=225210000;
#10;x=225220000;
#10;x=225230000;
#10;x=225240000;
#10;x=225250000;
#10;x=225260000;
#10;x=225270000;
#10;x=225280000;
#10;x=225290000;
#10;x=225300000;
#10;x=225310000;
#10;x=225320000;
#10;x=225330000;
#10;x=225340000;
#10;x=225350000;
#10;x=225360000;
#10;x=225370000;
#10;x=225380000;
#10;x=225390000;
#10;x=225400000;
#10;x=225410000;
#10;x=225420000;
#10;x=225430000;
#10;x=225440000;
#10;x=225450000;
#10;x=225460000;
#10;x=225470000;
#10;x=225480000;
#10;x=225490000;
#10;x=225500000;
#10;x=225510000;
#10;x=225520000;
#10;x=225530000;
#10;x=225540000;
#10;x=225550000;
#10;x=225560000;
#10;x=225570000;
#10;x=225580000;
#10;x=225590000;
#10;x=225600000;
#10;x=225610000;
#10;x=225620000;
#10;x=225630000;
#10;x=225640000;
#10;x=225650000;
#10;x=225660000;
#10;x=225670000;
#10;x=225680000;
#10;x=225690000;
#10;x=225700000;
#10;x=225710000;
#10;x=225720000;
#10;x=225730000;
#10;x=225740000;
#10;x=225750000;
#10;x=225760000;
#10;x=225770000;
#10;x=225780000;
#10;x=225790000;
#10;x=225800000;
#10;x=225810000;
#10;x=225820000;
#10;x=225830000;
#10;x=225840000;
#10;x=225850000;
#10;x=225860000;
#10;x=225870000;
#10;x=225880000;
#10;x=225890000;
#10;x=225900000;
#10;x=225910000;
#10;x=225920000;
#10;x=225930000;
#10;x=225940000;
#10;x=225950000;
#10;x=225960000;
#10;x=225970000;
#10;x=225980000;
#10;x=225990000;
#10;x=226000000;
#10;x=226010000;
#10;x=226020000;
#10;x=226030000;
#10;x=226040000;
#10;x=226050000;
#10;x=226060000;
#10;x=226070000;
#10;x=226080000;
#10;x=226090000;
#10;x=226100000;
#10;x=226110000;
#10;x=226120000;
#10;x=226130000;
#10;x=226140000;
#10;x=226150000;
#10;x=226160000;
#10;x=226170000;
#10;x=226180000;
#10;x=226190000;
#10;x=226200000;
#10;x=226210000;
#10;x=226220000;
#10;x=226230000;
#10;x=226240000;
#10;x=226250000;
#10;x=226260000;
#10;x=226270000;
#10;x=226280000;
#10;x=226290000;
#10;x=226300000;
#10;x=226310000;
#10;x=226320000;
#10;x=226330000;
#10;x=226340000;
#10;x=226350000;
#10;x=226360000;
#10;x=226370000;
#10;x=226380000;
#10;x=226390000;
#10;x=226400000;
#10;x=226410000;
#10;x=226420000;
#10;x=226430000;
#10;x=226440000;
#10;x=226450000;
#10;x=226460000;
#10;x=226470000;
#10;x=226480000;
#10;x=226490000;
#10;x=226500000;
#10;x=226510000;
#10;x=226520000;
#10;x=226530000;
#10;x=226540000;
#10;x=226550000;
#10;x=226560000;
#10;x=226570000;
#10;x=226580000;
#10;x=226590000;
#10;x=226600000;
#10;x=226610000;
#10;x=226620000;
#10;x=226630000;
#10;x=226640000;
#10;x=226650000;
#10;x=226660000;
#10;x=226670000;
#10;x=226680000;
#10;x=226690000;
#10;x=226700000;
#10;x=226710000;
#10;x=226720000;
#10;x=226730000;
#10;x=226740000;
#10;x=226750000;
#10;x=226760000;
#10;x=226770000;
#10;x=226780000;
#10;x=226790000;
#10;x=226800000;
#10;x=226810000;
#10;x=226820000;
#10;x=226830000;
#10;x=226840000;
#10;x=226850000;
#10;x=226860000;
#10;x=226870000;
#10;x=226880000;
#10;x=226890000;
#10;x=226900000;
#10;x=226910000;
#10;x=226920000;
#10;x=226930000;
#10;x=226940000;
#10;x=226950000;
#10;x=226960000;
#10;x=226970000;
#10;x=226980000;
#10;x=226990000;
#10;x=227000000;
#10;x=227010000;
#10;x=227020000;
#10;x=227030000;
#10;x=227040000;
#10;x=227050000;
#10;x=227060000;
#10;x=227070000;
#10;x=227080000;
#10;x=227090000;
#10;x=227100000;
#10;x=227110000;
#10;x=227120000;
#10;x=227130000;
#10;x=227140000;
#10;x=227150000;
#10;x=227160000;
#10;x=227170000;
#10;x=227180000;
#10;x=227190000;
#10;x=227200000;
#10;x=227210000;
#10;x=227220000;
#10;x=227230000;
#10;x=227240000;
#10;x=227250000;
#10;x=227260000;
#10;x=227270000;
#10;x=227280000;
#10;x=227290000;
#10;x=227300000;
#10;x=227310000;
#10;x=227320000;
#10;x=227330000;
#10;x=227340000;
#10;x=227350000;
#10;x=227360000;
#10;x=227370000;
#10;x=227380000;
#10;x=227390000;
#10;x=227400000;
#10;x=227410000;
#10;x=227420000;
#10;x=227430000;
#10;x=227440000;
#10;x=227450000;
#10;x=227460000;
#10;x=227470000;
#10;x=227480000;
#10;x=227490000;
#10;x=227500000;
#10;x=227510000;
#10;x=227520000;
#10;x=227530000;
#10;x=227540000;
#10;x=227550000;
#10;x=227560000;
#10;x=227570000;
#10;x=227580000;
#10;x=227590000;
#10;x=227600000;
#10;x=227610000;
#10;x=227620000;
#10;x=227630000;
#10;x=227640000;
#10;x=227650000;
#10;x=227660000;
#10;x=227670000;
#10;x=227680000;
#10;x=227690000;
#10;x=227700000;
#10;x=227710000;
#10;x=227720000;
#10;x=227730000;
#10;x=227740000;
#10;x=227750000;
#10;x=227760000;
#10;x=227770000;
#10;x=227780000;
#10;x=227790000;
#10;x=227800000;
#10;x=227810000;
#10;x=227820000;
#10;x=227830000;
#10;x=227840000;
#10;x=227850000;
#10;x=227860000;
#10;x=227870000;
#10;x=227880000;
#10;x=227890000;
#10;x=227900000;
#10;x=227910000;
#10;x=227920000;
#10;x=227930000;
#10;x=227940000;
#10;x=227950000;
#10;x=227960000;
#10;x=227970000;
#10;x=227980000;
#10;x=227990000;
#10;x=228000000;
#10;x=228010000;
#10;x=228020000;
#10;x=228030000;
#10;x=228040000;
#10;x=228050000;
#10;x=228060000;
#10;x=228070000;
#10;x=228080000;
#10;x=228090000;
#10;x=228100000;
#10;x=228110000;
#10;x=228120000;
#10;x=228130000;
#10;x=228140000;
#10;x=228150000;
#10;x=228160000;
#10;x=228170000;
#10;x=228180000;
#10;x=228190000;
#10;x=228200000;
#10;x=228210000;
#10;x=228220000;
#10;x=228230000;
#10;x=228240000;
#10;x=228250000;
#10;x=228260000;
#10;x=228270000;
#10;x=228280000;
#10;x=228290000;
#10;x=228300000;
#10;x=228310000;
#10;x=228320000;
#10;x=228330000;
#10;x=228340000;
#10;x=228350000;
#10;x=228360000;
#10;x=228370000;
#10;x=228380000;
#10;x=228390000;
#10;x=228400000;
#10;x=228410000;
#10;x=228420000;
#10;x=228430000;
#10;x=228440000;
#10;x=228450000;
#10;x=228460000;
#10;x=228470000;
#10;x=228480000;
#10;x=228490000;
#10;x=228500000;
#10;x=228510000;
#10;x=228520000;
#10;x=228530000;
#10;x=228540000;
#10;x=228550000;
#10;x=228560000;
#10;x=228570000;
#10;x=228580000;
#10;x=228590000;
#10;x=228600000;
#10;x=228610000;
#10;x=228620000;
#10;x=228630000;
#10;x=228640000;
#10;x=228650000;
#10;x=228660000;
#10;x=228670000;
#10;x=228680000;
#10;x=228690000;
#10;x=228700000;
#10;x=228710000;
#10;x=228720000;
#10;x=228730000;
#10;x=228740000;
#10;x=228750000;
#10;x=228760000;
#10;x=228770000;
#10;x=228780000;
#10;x=228790000;
#10;x=228800000;
#10;x=228810000;
#10;x=228820000;
#10;x=228830000;
#10;x=228840000;
#10;x=228850000;
#10;x=228860000;
#10;x=228870000;
#10;x=228880000;
#10;x=228890000;
#10;x=228900000;
#10;x=228910000;
#10;x=228920000;
#10;x=228930000;
#10;x=228940000;
#10;x=228950000;
#10;x=228960000;
#10;x=228970000;
#10;x=228980000;
#10;x=228990000;
#10;x=229000000;
#10;x=229010000;
#10;x=229020000;
#10;x=229030000;
#10;x=229040000;
#10;x=229050000;
#10;x=229060000;
#10;x=229070000;
#10;x=229080000;
#10;x=229090000;
#10;x=229100000;
#10;x=229110000;
#10;x=229120000;
#10;x=229130000;
#10;x=229140000;
#10;x=229150000;
#10;x=229160000;
#10;x=229170000;
#10;x=229180000;
#10;x=229190000;
#10;x=229200000;
#10;x=229210000;
#10;x=229220000;
#10;x=229230000;
#10;x=229240000;
#10;x=229250000;
#10;x=229260000;
#10;x=229270000;
#10;x=229280000;
#10;x=229290000;
#10;x=229300000;
#10;x=229310000;
#10;x=229320000;
#10;x=229330000;
#10;x=229340000;
#10;x=229350000;
#10;x=229360000;
#10;x=229370000;
#10;x=229380000;
#10;x=229390000;
#10;x=229400000;
#10;x=229410000;
#10;x=229420000;
#10;x=229430000;
#10;x=229440000;
#10;x=229450000;
#10;x=229460000;
#10;x=229470000;
#10;x=229480000;
#10;x=229490000;
#10;x=229500000;
#10;x=229510000;
#10;x=229520000;
#10;x=229530000;
#10;x=229540000;
#10;x=229550000;
#10;x=229560000;
#10;x=229570000;
#10;x=229580000;
#10;x=229590000;
#10;x=229600000;
#10;x=229610000;
#10;x=229620000;
#10;x=229630000;
#10;x=229640000;
#10;x=229650000;
#10;x=229660000;
#10;x=229670000;
#10;x=229680000;
#10;x=229690000;
#10;x=229700000;
#10;x=229710000;
#10;x=229720000;
#10;x=229730000;
#10;x=229740000;
#10;x=229750000;
#10;x=229760000;
#10;x=229770000;
#10;x=229780000;
#10;x=229790000;
#10;x=229800000;
#10;x=229810000;
#10;x=229820000;
#10;x=229830000;
#10;x=229840000;
#10;x=229850000;
#10;x=229860000;
#10;x=229870000;
#10;x=229880000;
#10;x=229890000;
#10;x=229900000;
#10;x=229910000;
#10;x=229920000;
#10;x=229930000;
#10;x=229940000;
#10;x=229950000;
#10;x=229960000;
#10;x=229970000;
#10;x=229980000;
#10;x=229990000;
#10;x=230000000;
#10;x=230010000;
#10;x=230020000;
#10;x=230030000;
#10;x=230040000;
#10;x=230050000;
#10;x=230060000;
#10;x=230070000;
#10;x=230080000;
#10;x=230090000;
#10;x=230100000;
#10;x=230110000;
#10;x=230120000;
#10;x=230130000;
#10;x=230140000;
#10;x=230150000;
#10;x=230160000;
#10;x=230170000;
#10;x=230180000;
#10;x=230190000;
#10;x=230200000;
#10;x=230210000;
#10;x=230220000;
#10;x=230230000;
#10;x=230240000;
#10;x=230250000;
#10;x=230260000;
#10;x=230270000;
#10;x=230280000;
#10;x=230290000;
#10;x=230300000;
#10;x=230310000;
#10;x=230320000;
#10;x=230330000;
#10;x=230340000;
#10;x=230350000;
#10;x=230360000;
#10;x=230370000;
#10;x=230380000;
#10;x=230390000;
#10;x=230400000;
#10;x=230410000;
#10;x=230420000;
#10;x=230430000;
#10;x=230440000;
#10;x=230450000;
#10;x=230460000;
#10;x=230470000;
#10;x=230480000;
#10;x=230490000;
#10;x=230500000;
#10;x=230510000;
#10;x=230520000;
#10;x=230530000;
#10;x=230540000;
#10;x=230550000;
#10;x=230560000;
#10;x=230570000;
#10;x=230580000;
#10;x=230590000;
#10;x=230600000;
#10;x=230610000;
#10;x=230620000;
#10;x=230630000;
#10;x=230640000;
#10;x=230650000;
#10;x=230660000;
#10;x=230670000;
#10;x=230680000;
#10;x=230690000;
#10;x=230700000;
#10;x=230710000;
#10;x=230720000;
#10;x=230730000;
#10;x=230740000;
#10;x=230750000;
#10;x=230760000;
#10;x=230770000;
#10;x=230780000;
#10;x=230790000;
#10;x=230800000;
#10;x=230810000;
#10;x=230820000;
#10;x=230830000;
#10;x=230840000;
#10;x=230850000;
#10;x=230860000;
#10;x=230870000;
#10;x=230880000;
#10;x=230890000;
#10;x=230900000;
#10;x=230910000;
#10;x=230920000;
#10;x=230930000;
#10;x=230940000;
#10;x=230950000;
#10;x=230960000;
#10;x=230970000;
#10;x=230980000;
#10;x=230990000;
#10;x=231000000;
#10;x=231010000;
#10;x=231020000;
#10;x=231030000;
#10;x=231040000;
#10;x=231050000;
#10;x=231060000;
#10;x=231070000;
#10;x=231080000;
#10;x=231090000;
#10;x=231100000;
#10;x=231110000;
#10;x=231120000;
#10;x=231130000;
#10;x=231140000;
#10;x=231150000;
#10;x=231160000;
#10;x=231170000;
#10;x=231180000;
#10;x=231190000;
#10;x=231200000;
#10;x=231210000;
#10;x=231220000;
#10;x=231230000;
#10;x=231240000;
#10;x=231250000;
#10;x=231260000;
#10;x=231270000;
#10;x=231280000;
#10;x=231290000;
#10;x=231300000;
#10;x=231310000;
#10;x=231320000;
#10;x=231330000;
#10;x=231340000;
#10;x=231350000;
#10;x=231360000;
#10;x=231370000;
#10;x=231380000;
#10;x=231390000;
#10;x=231400000;
#10;x=231410000;
#10;x=231420000;
#10;x=231430000;
#10;x=231440000;
#10;x=231450000;
#10;x=231460000;
#10;x=231470000;
#10;x=231480000;
#10;x=231490000;
#10;x=231500000;
#10;x=231510000;
#10;x=231520000;
#10;x=231530000;
#10;x=231540000;
#10;x=231550000;
#10;x=231560000;
#10;x=231570000;
#10;x=231580000;
#10;x=231590000;
#10;x=231600000;
#10;x=231610000;
#10;x=231620000;
#10;x=231630000;
#10;x=231640000;
#10;x=231650000;
#10;x=231660000;
#10;x=231670000;
#10;x=231680000;
#10;x=231690000;
#10;x=231700000;
#10;x=231710000;
#10;x=231720000;
#10;x=231730000;
#10;x=231740000;
#10;x=231750000;
#10;x=231760000;
#10;x=231770000;
#10;x=231780000;
#10;x=231790000;
#10;x=231800000;
#10;x=231810000;
#10;x=231820000;
#10;x=231830000;
#10;x=231840000;
#10;x=231850000;
#10;x=231860000;
#10;x=231870000;
#10;x=231880000;
#10;x=231890000;
#10;x=231900000;
#10;x=231910000;
#10;x=231920000;
#10;x=231930000;
#10;x=231940000;
#10;x=231950000;
#10;x=231960000;
#10;x=231970000;
#10;x=231980000;
#10;x=231990000;
#10;x=232000000;
#10;x=232010000;
#10;x=232020000;
#10;x=232030000;
#10;x=232040000;
#10;x=232050000;
#10;x=232060000;
#10;x=232070000;
#10;x=232080000;
#10;x=232090000;
#10;x=232100000;
#10;x=232110000;
#10;x=232120000;
#10;x=232130000;
#10;x=232140000;
#10;x=232150000;
#10;x=232160000;
#10;x=232170000;
#10;x=232180000;
#10;x=232190000;
#10;x=232200000;
#10;x=232210000;
#10;x=232220000;
#10;x=232230000;
#10;x=232240000;
#10;x=232250000;
#10;x=232260000;
#10;x=232270000;
#10;x=232280000;
#10;x=232290000;
#10;x=232300000;
#10;x=232310000;
#10;x=232320000;
#10;x=232330000;
#10;x=232340000;
#10;x=232350000;
#10;x=232360000;
#10;x=232370000;
#10;x=232380000;
#10;x=232390000;
#10;x=232400000;
#10;x=232410000;
#10;x=232420000;
#10;x=232430000;
#10;x=232440000;
#10;x=232450000;
#10;x=232460000;
#10;x=232470000;
#10;x=232480000;
#10;x=232490000;
#10;x=232500000;
#10;x=232510000;
#10;x=232520000;
#10;x=232530000;
#10;x=232540000;
#10;x=232550000;
#10;x=232560000;
#10;x=232570000;
#10;x=232580000;
#10;x=232590000;
#10;x=232600000;
#10;x=232610000;
#10;x=232620000;
#10;x=232630000;
#10;x=232640000;
#10;x=232650000;
#10;x=232660000;
#10;x=232670000;
#10;x=232680000;
#10;x=232690000;
#10;x=232700000;
#10;x=232710000;
#10;x=232720000;
#10;x=232730000;
#10;x=232740000;
#10;x=232750000;
#10;x=232760000;
#10;x=232770000;
#10;x=232780000;
#10;x=232790000;
#10;x=232800000;
#10;x=232810000;
#10;x=232820000;
#10;x=232830000;
#10;x=232840000;
#10;x=232850000;
#10;x=232860000;
#10;x=232870000;
#10;x=232880000;
#10;x=232890000;
#10;x=232900000;
#10;x=232910000;
#10;x=232920000;
#10;x=232930000;
#10;x=232940000;
#10;x=232950000;
#10;x=232960000;
#10;x=232970000;
#10;x=232980000;
#10;x=232990000;
#10;x=233000000;
#10;x=233010000;
#10;x=233020000;
#10;x=233030000;
#10;x=233040000;
#10;x=233050000;
#10;x=233060000;
#10;x=233070000;
#10;x=233080000;
#10;x=233090000;
#10;x=233100000;
#10;x=233110000;
#10;x=233120000;
#10;x=233130000;
#10;x=233140000;
#10;x=233150000;
#10;x=233160000;
#10;x=233170000;
#10;x=233180000;
#10;x=233190000;
#10;x=233200000;
#10;x=233210000;
#10;x=233220000;
#10;x=233230000;
#10;x=233240000;
#10;x=233250000;
#10;x=233260000;
#10;x=233270000;
#10;x=233280000;
#10;x=233290000;
#10;x=233300000;
#10;x=233310000;
#10;x=233320000;
#10;x=233330000;
#10;x=233340000;
#10;x=233350000;
#10;x=233360000;
#10;x=233370000;
#10;x=233380000;
#10;x=233390000;
#10;x=233400000;
#10;x=233410000;
#10;x=233420000;
#10;x=233430000;
#10;x=233440000;
#10;x=233450000;
#10;x=233460000;
#10;x=233470000;
#10;x=233480000;
#10;x=233490000;
#10;x=233500000;
#10;x=233510000;
#10;x=233520000;
#10;x=233530000;
#10;x=233540000;
#10;x=233550000;
#10;x=233560000;
#10;x=233570000;
#10;x=233580000;
#10;x=233590000;
#10;x=233600000;
#10;x=233610000;
#10;x=233620000;
#10;x=233630000;
#10;x=233640000;
#10;x=233650000;
#10;x=233660000;
#10;x=233670000;
#10;x=233680000;
#10;x=233690000;
#10;x=233700000;
#10;x=233710000;
#10;x=233720000;
#10;x=233730000;
#10;x=233740000;
#10;x=233750000;
#10;x=233760000;
#10;x=233770000;
#10;x=233780000;
#10;x=233790000;
#10;x=233800000;
#10;x=233810000;
#10;x=233820000;
#10;x=233830000;
#10;x=233840000;
#10;x=233850000;
#10;x=233860000;
#10;x=233870000;
#10;x=233880000;
#10;x=233890000;
#10;x=233900000;
#10;x=233910000;
#10;x=233920000;
#10;x=233930000;
#10;x=233940000;
#10;x=233950000;
#10;x=233960000;
#10;x=233970000;
#10;x=233980000;
#10;x=233990000;
#10;x=234000000;
#10;x=234010000;
#10;x=234020000;
#10;x=234030000;
#10;x=234040000;
#10;x=234050000;
#10;x=234060000;
#10;x=234070000;
#10;x=234080000;
#10;x=234090000;
#10;x=234100000;
#10;x=234110000;
#10;x=234120000;
#10;x=234130000;
#10;x=234140000;
#10;x=234150000;
#10;x=234160000;
#10;x=234170000;
#10;x=234180000;
#10;x=234190000;
#10;x=234200000;
#10;x=234210000;
#10;x=234220000;
#10;x=234230000;
#10;x=234240000;
#10;x=234250000;
#10;x=234260000;
#10;x=234270000;
#10;x=234280000;
#10;x=234290000;
#10;x=234300000;
#10;x=234310000;
#10;x=234320000;
#10;x=234330000;
#10;x=234340000;
#10;x=234350000;
#10;x=234360000;
#10;x=234370000;
#10;x=234380000;
#10;x=234390000;
#10;x=234400000;
#10;x=234410000;
#10;x=234420000;
#10;x=234430000;
#10;x=234440000;
#10;x=234450000;
#10;x=234460000;
#10;x=234470000;
#10;x=234480000;
#10;x=234490000;
#10;x=234500000;
#10;x=234510000;
#10;x=234520000;
#10;x=234530000;
#10;x=234540000;
#10;x=234550000;
#10;x=234560000;
#10;x=234570000;
#10;x=234580000;
#10;x=234590000;
#10;x=234600000;
#10;x=234610000;
#10;x=234620000;
#10;x=234630000;
#10;x=234640000;
#10;x=234650000;
#10;x=234660000;
#10;x=234670000;
#10;x=234680000;
#10;x=234690000;
#10;x=234700000;
#10;x=234710000;
#10;x=234720000;
#10;x=234730000;
#10;x=234740000;
#10;x=234750000;
#10;x=234760000;
#10;x=234770000;
#10;x=234780000;
#10;x=234790000;
#10;x=234800000;
#10;x=234810000;
#10;x=234820000;
#10;x=234830000;
#10;x=234840000;
#10;x=234850000;
#10;x=234860000;
#10;x=234870000;
#10;x=234880000;
#10;x=234890000;
#10;x=234900000;
#10;x=234910000;
#10;x=234920000;
#10;x=234930000;
#10;x=234940000;
#10;x=234950000;
#10;x=234960000;
#10;x=234970000;
#10;x=234980000;
#10;x=234990000;
#10;x=235000000;
#10;x=235010000;
#10;x=235020000;
#10;x=235030000;
#10;x=235040000;
#10;x=235050000;
#10;x=235060000;
#10;x=235070000;
#10;x=235080000;
#10;x=235090000;
#10;x=235100000;
#10;x=235110000;
#10;x=235120000;
#10;x=235130000;
#10;x=235140000;
#10;x=235150000;
#10;x=235160000;
#10;x=235170000;
#10;x=235180000;
#10;x=235190000;
#10;x=235200000;
#10;x=235210000;
#10;x=235220000;
#10;x=235230000;
#10;x=235240000;
#10;x=235250000;
#10;x=235260000;
#10;x=235270000;
#10;x=235280000;
#10;x=235290000;
#10;x=235300000;
#10;x=235310000;
#10;x=235320000;
#10;x=235330000;
#10;x=235340000;
#10;x=235350000;
#10;x=235360000;
#10;x=235370000;
#10;x=235380000;
#10;x=235390000;
#10;x=235400000;
#10;x=235410000;
#10;x=235420000;
#10;x=235430000;
#10;x=235440000;
#10;x=235450000;
#10;x=235460000;
#10;x=235470000;
#10;x=235480000;
#10;x=235490000;
#10;x=235500000;
#10;x=235510000;
#10;x=235520000;
#10;x=235530000;
#10;x=235540000;
#10;x=235550000;
#10;x=235560000;
#10;x=235570000;
#10;x=235580000;
#10;x=235590000;
#10;x=235600000;
#10;x=235610000;
#10;x=235620000;
#10;x=235630000;
#10;x=235640000;
#10;x=235650000;
#10;x=235660000;
#10;x=235670000;
#10;x=235680000;
#10;x=235690000;
#10;x=235700000;
#10;x=235710000;
#10;x=235720000;
#10;x=235730000;
#10;x=235740000;
#10;x=235750000;
#10;x=235760000;
#10;x=235770000;
#10;x=235780000;
#10;x=235790000;
#10;x=235800000;
#10;x=235810000;
#10;x=235820000;
#10;x=235830000;
#10;x=235840000;
#10;x=235850000;
#10;x=235860000;
#10;x=235870000;
#10;x=235880000;
#10;x=235890000;
#10;x=235900000;
#10;x=235910000;
#10;x=235920000;
#10;x=235930000;
#10;x=235940000;
#10;x=235950000;
#10;x=235960000;
#10;x=235970000;
#10;x=235980000;
#10;x=235990000;
#10;x=236000000;
#10;x=236010000;
#10;x=236020000;
#10;x=236030000;
#10;x=236040000;
#10;x=236050000;
#10;x=236060000;
#10;x=236070000;
#10;x=236080000;
#10;x=236090000;
#10;x=236100000;
#10;x=236110000;
#10;x=236120000;
#10;x=236130000;
#10;x=236140000;
#10;x=236150000;
#10;x=236160000;
#10;x=236170000;
#10;x=236180000;
#10;x=236190000;
#10;x=236200000;
#10;x=236210000;
#10;x=236220000;
#10;x=236230000;
#10;x=236240000;
#10;x=236250000;
#10;x=236260000;
#10;x=236270000;
#10;x=236280000;
#10;x=236290000;
#10;x=236300000;
#10;x=236310000;
#10;x=236320000;
#10;x=236330000;
#10;x=236340000;
#10;x=236350000;
#10;x=236360000;
#10;x=236370000;
#10;x=236380000;
#10;x=236390000;
#10;x=236400000;
#10;x=236410000;
#10;x=236420000;
#10;x=236430000;
#10;x=236440000;
#10;x=236450000;
#10;x=236460000;
#10;x=236470000;
#10;x=236480000;
#10;x=236490000;
#10;x=236500000;
#10;x=236510000;
#10;x=236520000;
#10;x=236530000;
#10;x=236540000;
#10;x=236550000;
#10;x=236560000;
#10;x=236570000;
#10;x=236580000;
#10;x=236590000;
#10;x=236600000;
#10;x=236610000;
#10;x=236620000;
#10;x=236630000;
#10;x=236640000;
#10;x=236650000;
#10;x=236660000;
#10;x=236670000;
#10;x=236680000;
#10;x=236690000;
#10;x=236700000;
#10;x=236710000;
#10;x=236720000;
#10;x=236730000;
#10;x=236740000;
#10;x=236750000;
#10;x=236760000;
#10;x=236770000;
#10;x=236780000;
#10;x=236790000;
#10;x=236800000;
#10;x=236810000;
#10;x=236820000;
#10;x=236830000;
#10;x=236840000;
#10;x=236850000;
#10;x=236860000;
#10;x=236870000;
#10;x=236880000;
#10;x=236890000;
#10;x=236900000;
#10;x=236910000;
#10;x=236920000;
#10;x=236930000;
#10;x=236940000;
#10;x=236950000;
#10;x=236960000;
#10;x=236970000;
#10;x=236980000;
#10;x=236990000;
#10;x=237000000;
#10;x=237010000;
#10;x=237020000;
#10;x=237030000;
#10;x=237040000;
#10;x=237050000;
#10;x=237060000;
#10;x=237070000;
#10;x=237080000;
#10;x=237090000;
#10;x=237100000;
#10;x=237110000;
#10;x=237120000;
#10;x=237130000;
#10;x=237140000;
#10;x=237150000;
#10;x=237160000;
#10;x=237170000;
#10;x=237180000;
#10;x=237190000;
#10;x=237200000;
#10;x=237210000;
#10;x=237220000;
#10;x=237230000;
#10;x=237240000;
#10;x=237250000;
#10;x=237260000;
#10;x=237270000;
#10;x=237280000;
#10;x=237290000;
#10;x=237300000;
#10;x=237310000;
#10;x=237320000;
#10;x=237330000;
#10;x=237340000;
#10;x=237350000;
#10;x=237360000;
#10;x=237370000;
#10;x=237380000;
#10;x=237390000;
#10;x=237400000;
#10;x=237410000;
#10;x=237420000;
#10;x=237430000;
#10;x=237440000;
#10;x=237450000;
#10;x=237460000;
#10;x=237470000;
#10;x=237480000;
#10;x=237490000;
#10;x=237500000;
#10;x=237510000;
#10;x=237520000;
#10;x=237530000;
#10;x=237540000;
#10;x=237550000;
#10;x=237560000;
#10;x=237570000;
#10;x=237580000;
#10;x=237590000;
#10;x=237600000;
#10;x=237610000;
#10;x=237620000;
#10;x=237630000;
#10;x=237640000;
#10;x=237650000;
#10;x=237660000;
#10;x=237670000;
#10;x=237680000;
#10;x=237690000;
#10;x=237700000;
#10;x=237710000;
#10;x=237720000;
#10;x=237730000;
#10;x=237740000;
#10;x=237750000;
#10;x=237760000;
#10;x=237770000;
#10;x=237780000;
#10;x=237790000;
#10;x=237800000;
#10;x=237810000;
#10;x=237820000;
#10;x=237830000;
#10;x=237840000;
#10;x=237850000;
#10;x=237860000;
#10;x=237870000;
#10;x=237880000;
#10;x=237890000;
#10;x=237900000;
#10;x=237910000;
#10;x=237920000;
#10;x=237930000;
#10;x=237940000;
#10;x=237950000;
#10;x=237960000;
#10;x=237970000;
#10;x=237980000;
#10;x=237990000;
#10;x=238000000;
#10;x=238010000;
#10;x=238020000;
#10;x=238030000;
#10;x=238040000;
#10;x=238050000;
#10;x=238060000;
#10;x=238070000;
#10;x=238080000;
#10;x=238090000;
#10;x=238100000;
#10;x=238110000;
#10;x=238120000;
#10;x=238130000;
#10;x=238140000;
#10;x=238150000;
#10;x=238160000;
#10;x=238170000;
#10;x=238180000;
#10;x=238190000;
#10;x=238200000;
#10;x=238210000;
#10;x=238220000;
#10;x=238230000;
#10;x=238240000;
#10;x=238250000;
#10;x=238260000;
#10;x=238270000;
#10;x=238280000;
#10;x=238290000;
#10;x=238300000;
#10;x=238310000;
#10;x=238320000;
#10;x=238330000;
#10;x=238340000;
#10;x=238350000;
#10;x=238360000;
#10;x=238370000;
#10;x=238380000;
#10;x=238390000;
#10;x=238400000;
#10;x=238410000;
#10;x=238420000;
#10;x=238430000;
#10;x=238440000;
#10;x=238450000;
#10;x=238460000;
#10;x=238470000;
#10;x=238480000;
#10;x=238490000;
#10;x=238500000;
#10;x=238510000;
#10;x=238520000;
#10;x=238530000;
#10;x=238540000;
#10;x=238550000;
#10;x=238560000;
#10;x=238570000;
#10;x=238580000;
#10;x=238590000;
#10;x=238600000;
#10;x=238610000;
#10;x=238620000;
#10;x=238630000;
#10;x=238640000;
#10;x=238650000;
#10;x=238660000;
#10;x=238670000;
#10;x=238680000;
#10;x=238690000;
#10;x=238700000;
#10;x=238710000;
#10;x=238720000;
#10;x=238730000;
#10;x=238740000;
#10;x=238750000;
#10;x=238760000;
#10;x=238770000;
#10;x=238780000;
#10;x=238790000;
#10;x=238800000;
#10;x=238810000;
#10;x=238820000;
#10;x=238830000;
#10;x=238840000;
#10;x=238850000;
#10;x=238860000;
#10;x=238870000;
#10;x=238880000;
#10;x=238890000;
#10;x=238900000;
#10;x=238910000;
#10;x=238920000;
#10;x=238930000;
#10;x=238940000;
#10;x=238950000;
#10;x=238960000;
#10;x=238970000;
#10;x=238980000;
#10;x=238990000;
#10;x=239000000;
#10;x=239010000;
#10;x=239020000;
#10;x=239030000;
#10;x=239040000;
#10;x=239050000;
#10;x=239060000;
#10;x=239070000;
#10;x=239080000;
#10;x=239090000;
#10;x=239100000;
#10;x=239110000;
#10;x=239120000;
#10;x=239130000;
#10;x=239140000;
#10;x=239150000;
#10;x=239160000;
#10;x=239170000;
#10;x=239180000;
#10;x=239190000;
#10;x=239200000;
#10;x=239210000;
#10;x=239220000;
#10;x=239230000;
#10;x=239240000;
#10;x=239250000;
#10;x=239260000;
#10;x=239270000;
#10;x=239280000;
#10;x=239290000;
#10;x=239300000;
#10;x=239310000;
#10;x=239320000;
#10;x=239330000;
#10;x=239340000;
#10;x=239350000;
#10;x=239360000;
#10;x=239370000;
#10;x=239380000;
#10;x=239390000;
#10;x=239400000;
#10;x=239410000;
#10;x=239420000;
#10;x=239430000;
#10;x=239440000;
#10;x=239450000;
#10;x=239460000;
#10;x=239470000;
#10;x=239480000;
#10;x=239490000;
#10;x=239500000;
#10;x=239510000;
#10;x=239520000;
#10;x=239530000;
#10;x=239540000;
#10;x=239550000;
#10;x=239560000;
#10;x=239570000;
#10;x=239580000;
#10;x=239590000;
#10;x=239600000;
#10;x=239610000;
#10;x=239620000;
#10;x=239630000;
#10;x=239640000;
#10;x=239650000;
#10;x=239660000;
#10;x=239670000;
#10;x=239680000;
#10;x=239690000;
#10;x=239700000;
#10;x=239710000;
#10;x=239720000;
#10;x=239730000;
#10;x=239740000;
#10;x=239750000;
#10;x=239760000;
#10;x=239770000;
#10;x=239780000;
#10;x=239790000;
#10;x=239800000;
#10;x=239810000;
#10;x=239820000;
#10;x=239830000;
#10;x=239840000;
#10;x=239850000;
#10;x=239860000;
#10;x=239870000;
#10;x=239880000;
#10;x=239890000;
#10;x=239900000;
#10;x=239910000;
#10;x=239920000;
#10;x=239930000;
#10;x=239940000;
#10;x=239950000;
#10;x=239960000;
#10;x=239970000;
#10;x=239980000;
#10;x=239990000;
#10;x=240000000;

        #10;
        $finish;
    end
    
    // Monitor
    always @(posedge clk) begin
        $display("%d, %d", x, y);
    end
    
endmodule
