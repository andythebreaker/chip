`include "tanh.sv"
module tanh_tb; reg signed [31:0] x; wire signed [31:0] y; tanh dut (.x(x),
                                                                     .y(y));
    
    // Clock
    reg clk;
    
    // Initialize clock
    initial begin
        clk            = 0;
        forever #5 clk = ~clk;
    end
    
    // Stimulus
    initial begin
        #10;x=-2147483648;
#10;x=-2146483648;
#10;x=-2145483648;
#10;x=-2144483648;
#10;x=-2143483648;
#10;x=-2142483648;
#10;x=-2141483648;
#10;x=-2140483648;
#10;x=-2139483648;
#10;x=-2138483648;
#10;x=-2137483648;
#10;x=-2136483648;
#10;x=-2135483648;
#10;x=-2134483648;
#10;x=-2133483648;
#10;x=-2132483648;
#10;x=-2131483648;
#10;x=-2130483648;
#10;x=-2129483648;
#10;x=-2128483648;
#10;x=-2127483648;
#10;x=-2126483648;
#10;x=-2125483648;
#10;x=-2124483648;
#10;x=-2123483648;
#10;x=-2122483648;
#10;x=-2121483648;
#10;x=-2120483648;
#10;x=-2119483648;
#10;x=-2118483648;
#10;x=-2117483648;
#10;x=-2116483648;
#10;x=-2115483648;
#10;x=-2114483648;
#10;x=-2113483648;
#10;x=-2112483648;
#10;x=-2111483648;
#10;x=-2110483648;
#10;x=-2109483648;
#10;x=-2108483648;
#10;x=-2107483648;
#10;x=-2106483648;
#10;x=-2105483648;
#10;x=-2104483648;
#10;x=-2103483648;
#10;x=-2102483648;
#10;x=-2101483648;
#10;x=-2100483648;
#10;x=-2099483648;
#10;x=-2098483648;
#10;x=-2097483648;
#10;x=-2096483648;
#10;x=-2095483648;
#10;x=-2094483648;
#10;x=-2093483648;
#10;x=-2092483648;
#10;x=-2091483648;
#10;x=-2090483648;
#10;x=-2089483648;
#10;x=-2088483648;
#10;x=-2087483648;
#10;x=-2086483648;
#10;x=-2085483648;
#10;x=-2084483648;
#10;x=-2083483648;
#10;x=-2082483648;
#10;x=-2081483648;
#10;x=-2080483648;
#10;x=-2079483648;
#10;x=-2078483648;
#10;x=-2077483648;
#10;x=-2076483648;
#10;x=-2075483648;
#10;x=-2074483648;
#10;x=-2073483648;
#10;x=-2072483648;
#10;x=-2071483648;
#10;x=-2070483648;
#10;x=-2069483648;
#10;x=-2068483648;
#10;x=-2067483648;
#10;x=-2066483648;
#10;x=-2065483648;
#10;x=-2064483648;
#10;x=-2063483648;
#10;x=-2062483648;
#10;x=-2061483648;
#10;x=-2060483648;
#10;x=-2059483648;
#10;x=-2058483648;
#10;x=-2057483648;
#10;x=-2056483648;
#10;x=-2055483648;
#10;x=-2054483648;
#10;x=-2053483648;
#10;x=-2052483648;
#10;x=-2051483648;
#10;x=-2050483648;
#10;x=-2049483648;
#10;x=-2048483648;
#10;x=-2047483648;
#10;x=-2046483648;
#10;x=-2045483648;
#10;x=-2044483648;
#10;x=-2043483648;
#10;x=-2042483648;
#10;x=-2041483648;
#10;x=-2040483648;
#10;x=-2039483648;
#10;x=-2038483648;
#10;x=-2037483648;
#10;x=-2036483648;
#10;x=-2035483648;
#10;x=-2034483648;
#10;x=-2033483648;
#10;x=-2032483648;
#10;x=-2031483648;
#10;x=-2030483648;
#10;x=-2029483648;
#10;x=-2028483648;
#10;x=-2027483648;
#10;x=-2026483648;
#10;x=-2025483648;
#10;x=-2024483648;
#10;x=-2023483648;
#10;x=-2022483648;
#10;x=-2021483648;
#10;x=-2020483648;
#10;x=-2019483648;
#10;x=-2018483648;
#10;x=-2017483648;
#10;x=-2016483648;
#10;x=-2015483648;
#10;x=-2014483648;
#10;x=-2013483648;
#10;x=-2012483648;
#10;x=-2011483648;
#10;x=-2010483648;
#10;x=-2009483648;
#10;x=-2008483648;
#10;x=-2007483648;
#10;x=-2006483648;
#10;x=-2005483648;
#10;x=-2004483648;
#10;x=-2003483648;
#10;x=-2002483648;
#10;x=-2001483648;
#10;x=-2000483648;
#10;x=-1999483648;
#10;x=-1998483648;
#10;x=-1997483648;
#10;x=-1996483648;
#10;x=-1995483648;
#10;x=-1994483648;
#10;x=-1993483648;
#10;x=-1992483648;
#10;x=-1991483648;
#10;x=-1990483648;
#10;x=-1989483648;
#10;x=-1988483648;
#10;x=-1987483648;
#10;x=-1986483648;
#10;x=-1985483648;
#10;x=-1984483648;
#10;x=-1983483648;
#10;x=-1982483648;
#10;x=-1981483648;
#10;x=-1980483648;
#10;x=-1979483648;
#10;x=-1978483648;
#10;x=-1977483648;
#10;x=-1976483648;
#10;x=-1975483648;
#10;x=-1974483648;
#10;x=-1973483648;
#10;x=-1972483648;
#10;x=-1971483648;
#10;x=-1970483648;
#10;x=-1969483648;
#10;x=-1968483648;
#10;x=-1967483648;
#10;x=-1966483648;
#10;x=-1965483648;
#10;x=-1964483648;
#10;x=-1963483648;
#10;x=-1962483648;
#10;x=-1961483648;
#10;x=-1960483648;
#10;x=-1959483648;
#10;x=-1958483648;
#10;x=-1957483648;
#10;x=-1956483648;
#10;x=-1955483648;
#10;x=-1954483648;
#10;x=-1953483648;
#10;x=-1952483648;
#10;x=-1951483648;
#10;x=-1950483648;
#10;x=-1949483648;
#10;x=-1948483648;
#10;x=-1947483648;
#10;x=-1946483648;
#10;x=-1945483648;
#10;x=-1944483648;
#10;x=-1943483648;
#10;x=-1942483648;
#10;x=-1941483648;
#10;x=-1940483648;
#10;x=-1939483648;
#10;x=-1938483648;
#10;x=-1937483648;
#10;x=-1936483648;
#10;x=-1935483648;
#10;x=-1934483648;
#10;x=-1933483648;
#10;x=-1932483648;
#10;x=-1931483648;
#10;x=-1930483648;
#10;x=-1929483648;
#10;x=-1928483648;
#10;x=-1927483648;
#10;x=-1926483648;
#10;x=-1925483648;
#10;x=-1924483648;
#10;x=-1923483648;
#10;x=-1922483648;
#10;x=-1921483648;
#10;x=-1920483648;
#10;x=-1919483648;
#10;x=-1918483648;
#10;x=-1917483648;
#10;x=-1916483648;
#10;x=-1915483648;
#10;x=-1914483648;
#10;x=-1913483648;
#10;x=-1912483648;
#10;x=-1911483648;
#10;x=-1910483648;
#10;x=-1909483648;
#10;x=-1908483648;
#10;x=-1907483648;
#10;x=-1906483648;
#10;x=-1905483648;
#10;x=-1904483648;
#10;x=-1903483648;
#10;x=-1902483648;
#10;x=-1901483648;
#10;x=-1900483648;
#10;x=-1899483648;
#10;x=-1898483648;
#10;x=-1897483648;
#10;x=-1896483648;
#10;x=-1895483648;
#10;x=-1894483648;
#10;x=-1893483648;
#10;x=-1892483648;
#10;x=-1891483648;
#10;x=-1890483648;
#10;x=-1889483648;
#10;x=-1888483648;
#10;x=-1887483648;
#10;x=-1886483648;
#10;x=-1885483648;
#10;x=-1884483648;
#10;x=-1883483648;
#10;x=-1882483648;
#10;x=-1881483648;
#10;x=-1880483648;
#10;x=-1879483648;
#10;x=-1878483648;
#10;x=-1877483648;
#10;x=-1876483648;
#10;x=-1875483648;
#10;x=-1874483648;
#10;x=-1873483648;
#10;x=-1872483648;
#10;x=-1871483648;
#10;x=-1870483648;
#10;x=-1869483648;
#10;x=-1868483648;
#10;x=-1867483648;
#10;x=-1866483648;
#10;x=-1865483648;
#10;x=-1864483648;
#10;x=-1863483648;
#10;x=-1862483648;
#10;x=-1861483648;
#10;x=-1860483648;
#10;x=-1859483648;
#10;x=-1858483648;
#10;x=-1857483648;
#10;x=-1856483648;
#10;x=-1855483648;
#10;x=-1854483648;
#10;x=-1853483648;
#10;x=-1852483648;
#10;x=-1851483648;
#10;x=-1850483648;
#10;x=-1849483648;
#10;x=-1848483648;
#10;x=-1847483648;
#10;x=-1846483648;
#10;x=-1845483648;
#10;x=-1844483648;
#10;x=-1843483648;
#10;x=-1842483648;
#10;x=-1841483648;
#10;x=-1840483648;
#10;x=-1839483648;
#10;x=-1838483648;
#10;x=-1837483648;
#10;x=-1836483648;
#10;x=-1835483648;
#10;x=-1834483648;
#10;x=-1833483648;
#10;x=-1832483648;
#10;x=-1831483648;
#10;x=-1830483648;
#10;x=-1829483648;
#10;x=-1828483648;
#10;x=-1827483648;
#10;x=-1826483648;
#10;x=-1825483648;
#10;x=-1824483648;
#10;x=-1823483648;
#10;x=-1822483648;
#10;x=-1821483648;
#10;x=-1820483648;
#10;x=-1819483648;
#10;x=-1818483648;
#10;x=-1817483648;
#10;x=-1816483648;
#10;x=-1815483648;
#10;x=-1814483648;
#10;x=-1813483648;
#10;x=-1812483648;
#10;x=-1811483648;
#10;x=-1810483648;
#10;x=-1809483648;
#10;x=-1808483648;
#10;x=-1807483648;
#10;x=-1806483648;
#10;x=-1805483648;
#10;x=-1804483648;
#10;x=-1803483648;
#10;x=-1802483648;
#10;x=-1801483648;
#10;x=-1800483648;
#10;x=-1799483648;
#10;x=-1798483648;
#10;x=-1797483648;
#10;x=-1796483648;
#10;x=-1795483648;
#10;x=-1794483648;
#10;x=-1793483648;
#10;x=-1792483648;
#10;x=-1791483648;
#10;x=-1790483648;
#10;x=-1789483648;
#10;x=-1788483648;
#10;x=-1787483648;
#10;x=-1786483648;
#10;x=-1785483648;
#10;x=-1784483648;
#10;x=-1783483648;
#10;x=-1782483648;
#10;x=-1781483648;
#10;x=-1780483648;
#10;x=-1779483648;
#10;x=-1778483648;
#10;x=-1777483648;
#10;x=-1776483648;
#10;x=-1775483648;
#10;x=-1774483648;
#10;x=-1773483648;
#10;x=-1772483648;
#10;x=-1771483648;
#10;x=-1770483648;
#10;x=-1769483648;
#10;x=-1768483648;
#10;x=-1767483648;
#10;x=-1766483648;
#10;x=-1765483648;
#10;x=-1764483648;
#10;x=-1763483648;
#10;x=-1762483648;
#10;x=-1761483648;
#10;x=-1760483648;
#10;x=-1759483648;
#10;x=-1758483648;
#10;x=-1757483648;
#10;x=-1756483648;
#10;x=-1755483648;
#10;x=-1754483648;
#10;x=-1753483648;
#10;x=-1752483648;
#10;x=-1751483648;
#10;x=-1750483648;
#10;x=-1749483648;
#10;x=-1748483648;
#10;x=-1747483648;
#10;x=-1746483648;
#10;x=-1745483648;
#10;x=-1744483648;
#10;x=-1743483648;
#10;x=-1742483648;
#10;x=-1741483648;
#10;x=-1740483648;
#10;x=-1739483648;
#10;x=-1738483648;
#10;x=-1737483648;
#10;x=-1736483648;
#10;x=-1735483648;
#10;x=-1734483648;
#10;x=-1733483648;
#10;x=-1732483648;
#10;x=-1731483648;
#10;x=-1730483648;
#10;x=-1729483648;
#10;x=-1728483648;
#10;x=-1727483648;
#10;x=-1726483648;
#10;x=-1725483648;
#10;x=-1724483648;
#10;x=-1723483648;
#10;x=-1722483648;
#10;x=-1721483648;
#10;x=-1720483648;
#10;x=-1719483648;
#10;x=-1718483648;
#10;x=-1717483648;
#10;x=-1716483648;
#10;x=-1715483648;
#10;x=-1714483648;
#10;x=-1713483648;
#10;x=-1712483648;
#10;x=-1711483648;
#10;x=-1710483648;
#10;x=-1709483648;
#10;x=-1708483648;
#10;x=-1707483648;
#10;x=-1706483648;
#10;x=-1705483648;
#10;x=-1704483648;
#10;x=-1703483648;
#10;x=-1702483648;
#10;x=-1701483648;
#10;x=-1700483648;
#10;x=-1699483648;
#10;x=-1698483648;
#10;x=-1697483648;
#10;x=-1696483648;
#10;x=-1695483648;
#10;x=-1694483648;
#10;x=-1693483648;
#10;x=-1692483648;
#10;x=-1691483648;
#10;x=-1690483648;
#10;x=-1689483648;
#10;x=-1688483648;
#10;x=-1687483648;
#10;x=-1686483648;
#10;x=-1685483648;
#10;x=-1684483648;
#10;x=-1683483648;
#10;x=-1682483648;
#10;x=-1681483648;
#10;x=-1680483648;
#10;x=-1679483648;
#10;x=-1678483648;
#10;x=-1677483648;
#10;x=-1676483648;
#10;x=-1675483648;
#10;x=-1674483648;
#10;x=-1673483648;
#10;x=-1672483648;
#10;x=-1671483648;
#10;x=-1670483648;
#10;x=-1669483648;
#10;x=-1668483648;
#10;x=-1667483648;
#10;x=-1666483648;
#10;x=-1665483648;
#10;x=-1664483648;
#10;x=-1663483648;
#10;x=-1662483648;
#10;x=-1661483648;
#10;x=-1660483648;
#10;x=-1659483648;
#10;x=-1658483648;
#10;x=-1657483648;
#10;x=-1656483648;
#10;x=-1655483648;
#10;x=-1654483648;
#10;x=-1653483648;
#10;x=-1652483648;
#10;x=-1651483648;
#10;x=-1650483648;
#10;x=-1649483648;
#10;x=-1648483648;
#10;x=-1647483648;
#10;x=-1646483648;
#10;x=-1645483648;
#10;x=-1644483648;
#10;x=-1643483648;
#10;x=-1642483648;
#10;x=-1641483648;
#10;x=-1640483648;
#10;x=-1639483648;
#10;x=-1638483648;
#10;x=-1637483648;
#10;x=-1636483648;
#10;x=-1635483648;
#10;x=-1634483648;
#10;x=-1633483648;
#10;x=-1632483648;
#10;x=-1631483648;
#10;x=-1630483648;
#10;x=-1629483648;
#10;x=-1628483648;
#10;x=-1627483648;
#10;x=-1626483648;
#10;x=-1625483648;
#10;x=-1624483648;
#10;x=-1623483648;
#10;x=-1622483648;
#10;x=-1621483648;
#10;x=-1620483648;
#10;x=-1619483648;
#10;x=-1618483648;
#10;x=-1617483648;
#10;x=-1616483648;
#10;x=-1615483648;
#10;x=-1614483648;
#10;x=-1613483648;
#10;x=-1612483648;
#10;x=-1611483648;
#10;x=-1610483648;
#10;x=-1609483648;
#10;x=-1608483648;
#10;x=-1607483648;
#10;x=-1606483648;
#10;x=-1605483648;
#10;x=-1604483648;
#10;x=-1603483648;
#10;x=-1602483648;
#10;x=-1601483648;
#10;x=-1600483648;
#10;x=-1599483648;
#10;x=-1598483648;
#10;x=-1597483648;
#10;x=-1596483648;
#10;x=-1595483648;
#10;x=-1594483648;
#10;x=-1593483648;
#10;x=-1592483648;
#10;x=-1591483648;
#10;x=-1590483648;
#10;x=-1589483648;
#10;x=-1588483648;
#10;x=-1587483648;
#10;x=-1586483648;
#10;x=-1585483648;
#10;x=-1584483648;
#10;x=-1583483648;
#10;x=-1582483648;
#10;x=-1581483648;
#10;x=-1580483648;
#10;x=-1579483648;
#10;x=-1578483648;
#10;x=-1577483648;
#10;x=-1576483648;
#10;x=-1575483648;
#10;x=-1574483648;
#10;x=-1573483648;
#10;x=-1572483648;
#10;x=-1571483648;
#10;x=-1570483648;
#10;x=-1569483648;
#10;x=-1568483648;
#10;x=-1567483648;
#10;x=-1566483648;
#10;x=-1565483648;
#10;x=-1564483648;
#10;x=-1563483648;
#10;x=-1562483648;
#10;x=-1561483648;
#10;x=-1560483648;
#10;x=-1559483648;
#10;x=-1558483648;
#10;x=-1557483648;
#10;x=-1556483648;
#10;x=-1555483648;
#10;x=-1554483648;
#10;x=-1553483648;
#10;x=-1552483648;
#10;x=-1551483648;
#10;x=-1550483648;
#10;x=-1549483648;
#10;x=-1548483648;
#10;x=-1547483648;
#10;x=-1546483648;
#10;x=-1545483648;
#10;x=-1544483648;
#10;x=-1543483648;
#10;x=-1542483648;
#10;x=-1541483648;
#10;x=-1540483648;
#10;x=-1539483648;
#10;x=-1538483648;
#10;x=-1537483648;
#10;x=-1536483648;
#10;x=-1535483648;
#10;x=-1534483648;
#10;x=-1533483648;
#10;x=-1532483648;
#10;x=-1531483648;
#10;x=-1530483648;
#10;x=-1529483648;
#10;x=-1528483648;
#10;x=-1527483648;
#10;x=-1526483648;
#10;x=-1525483648;
#10;x=-1524483648;
#10;x=-1523483648;
#10;x=-1522483648;
#10;x=-1521483648;
#10;x=-1520483648;
#10;x=-1519483648;
#10;x=-1518483648;
#10;x=-1517483648;
#10;x=-1516483648;
#10;x=-1515483648;
#10;x=-1514483648;
#10;x=-1513483648;
#10;x=-1512483648;
#10;x=-1511483648;
#10;x=-1510483648;
#10;x=-1509483648;
#10;x=-1508483648;
#10;x=-1507483648;
#10;x=-1506483648;
#10;x=-1505483648;
#10;x=-1504483648;
#10;x=-1503483648;
#10;x=-1502483648;
#10;x=-1501483648;
#10;x=-1500483648;
#10;x=-1499483648;
#10;x=-1498483648;
#10;x=-1497483648;
#10;x=-1496483648;
#10;x=-1495483648;
#10;x=-1494483648;
#10;x=-1493483648;
#10;x=-1492483648;
#10;x=-1491483648;
#10;x=-1490483648;
#10;x=-1489483648;
#10;x=-1488483648;
#10;x=-1487483648;
#10;x=-1486483648;
#10;x=-1485483648;
#10;x=-1484483648;
#10;x=-1483483648;
#10;x=-1482483648;
#10;x=-1481483648;
#10;x=-1480483648;
#10;x=-1479483648;
#10;x=-1478483648;
#10;x=-1477483648;
#10;x=-1476483648;
#10;x=-1475483648;
#10;x=-1474483648;
#10;x=-1473483648;
#10;x=-1472483648;
#10;x=-1471483648;
#10;x=-1470483648;
#10;x=-1469483648;
#10;x=-1468483648;
#10;x=-1467483648;
#10;x=-1466483648;
#10;x=-1465483648;
#10;x=-1464483648;
#10;x=-1463483648;
#10;x=-1462483648;
#10;x=-1461483648;
#10;x=-1460483648;
#10;x=-1459483648;
#10;x=-1458483648;
#10;x=-1457483648;
#10;x=-1456483648;
#10;x=-1455483648;
#10;x=-1454483648;
#10;x=-1453483648;
#10;x=-1452483648;
#10;x=-1451483648;
#10;x=-1450483648;
#10;x=-1449483648;
#10;x=-1448483648;
#10;x=-1447483648;
#10;x=-1446483648;
#10;x=-1445483648;
#10;x=-1444483648;
#10;x=-1443483648;
#10;x=-1442483648;
#10;x=-1441483648;
#10;x=-1440483648;
#10;x=-1439483648;
#10;x=-1438483648;
#10;x=-1437483648;
#10;x=-1436483648;
#10;x=-1435483648;
#10;x=-1434483648;
#10;x=-1433483648;
#10;x=-1432483648;
#10;x=-1431483648;
#10;x=-1430483648;
#10;x=-1429483648;
#10;x=-1428483648;
#10;x=-1427483648;
#10;x=-1426483648;
#10;x=-1425483648;
#10;x=-1424483648;
#10;x=-1423483648;
#10;x=-1422483648;
#10;x=-1421483648;
#10;x=-1420483648;
#10;x=-1419483648;
#10;x=-1418483648;
#10;x=-1417483648;
#10;x=-1416483648;
#10;x=-1415483648;
#10;x=-1414483648;
#10;x=-1413483648;
#10;x=-1412483648;
#10;x=-1411483648;
#10;x=-1410483648;
#10;x=-1409483648;
#10;x=-1408483648;
#10;x=-1407483648;
#10;x=-1406483648;
#10;x=-1405483648;
#10;x=-1404483648;
#10;x=-1403483648;
#10;x=-1402483648;
#10;x=-1401483648;
#10;x=-1400483648;
#10;x=-1399483648;
#10;x=-1398483648;
#10;x=-1397483648;
#10;x=-1396483648;
#10;x=-1395483648;
#10;x=-1394483648;
#10;x=-1393483648;
#10;x=-1392483648;
#10;x=-1391483648;
#10;x=-1390483648;
#10;x=-1389483648;
#10;x=-1388483648;
#10;x=-1387483648;
#10;x=-1386483648;
#10;x=-1385483648;
#10;x=-1384483648;
#10;x=-1383483648;
#10;x=-1382483648;
#10;x=-1381483648;
#10;x=-1380483648;
#10;x=-1379483648;
#10;x=-1378483648;
#10;x=-1377483648;
#10;x=-1376483648;
#10;x=-1375483648;
#10;x=-1374483648;
#10;x=-1373483648;
#10;x=-1372483648;
#10;x=-1371483648;
#10;x=-1370483648;
#10;x=-1369483648;
#10;x=-1368483648;
#10;x=-1367483648;
#10;x=-1366483648;
#10;x=-1365483648;
#10;x=-1364483648;
#10;x=-1363483648;
#10;x=-1362483648;
#10;x=-1361483648;
#10;x=-1360483648;
#10;x=-1359483648;
#10;x=-1358483648;
#10;x=-1357483648;
#10;x=-1356483648;
#10;x=-1355483648;
#10;x=-1354483648;
#10;x=-1353483648;
#10;x=-1352483648;
#10;x=-1351483648;
#10;x=-1350483648;
#10;x=-1349483648;
#10;x=-1348483648;
#10;x=-1347483648;
#10;x=-1346483648;
#10;x=-1345483648;
#10;x=-1344483648;
#10;x=-1343483648;
#10;x=-1342483648;
#10;x=-1341483648;
#10;x=-1340483648;
#10;x=-1339483648;
#10;x=-1338483648;
#10;x=-1337483648;
#10;x=-1336483648;
#10;x=-1335483648;
#10;x=-1334483648;
#10;x=-1333483648;
#10;x=-1332483648;
#10;x=-1331483648;
#10;x=-1330483648;
#10;x=-1329483648;
#10;x=-1328483648;
#10;x=-1327483648;
#10;x=-1326483648;
#10;x=-1325483648;
#10;x=-1324483648;
#10;x=-1323483648;
#10;x=-1322483648;
#10;x=-1321483648;
#10;x=-1320483648;
#10;x=-1319483648;
#10;x=-1318483648;
#10;x=-1317483648;
#10;x=-1316483648;
#10;x=-1315483648;
#10;x=-1314483648;
#10;x=-1313483648;
#10;x=-1312483648;
#10;x=-1311483648;
#10;x=-1310483648;
#10;x=-1309483648;
#10;x=-1308483648;
#10;x=-1307483648;
#10;x=-1306483648;
#10;x=-1305483648;
#10;x=-1304483648;
#10;x=-1303483648;
#10;x=-1302483648;
#10;x=-1301483648;
#10;x=-1300483648;
#10;x=-1299483648;
#10;x=-1298483648;
#10;x=-1297483648;
#10;x=-1296483648;
#10;x=-1295483648;
#10;x=-1294483648;
#10;x=-1293483648;
#10;x=-1292483648;
#10;x=-1291483648;
#10;x=-1290483648;
#10;x=-1289483648;
#10;x=-1288483648;
#10;x=-1287483648;
#10;x=-1286483648;
#10;x=-1285483648;
#10;x=-1284483648;
#10;x=-1283483648;
#10;x=-1282483648;
#10;x=-1281483648;
#10;x=-1280483648;
#10;x=-1279483648;
#10;x=-1278483648;
#10;x=-1277483648;
#10;x=-1276483648;
#10;x=-1275483648;
#10;x=-1274483648;
#10;x=-1273483648;
#10;x=-1272483648;
#10;x=-1271483648;
#10;x=-1270483648;
#10;x=-1269483648;
#10;x=-1268483648;
#10;x=-1267483648;
#10;x=-1266483648;
#10;x=-1265483648;
#10;x=-1264483648;
#10;x=-1263483648;
#10;x=-1262483648;
#10;x=-1261483648;
#10;x=-1260483648;
#10;x=-1259483648;
#10;x=-1258483648;
#10;x=-1257483648;
#10;x=-1256483648;
#10;x=-1255483648;
#10;x=-1254483648;
#10;x=-1253483648;
#10;x=-1252483648;
#10;x=-1251483648;
#10;x=-1250483648;
#10;x=-1249483648;
#10;x=-1248483648;
#10;x=-1247483648;
#10;x=-1246483648;
#10;x=-1245483648;
#10;x=-1244483648;
#10;x=-1243483648;
#10;x=-1242483648;
#10;x=-1241483648;
#10;x=-1240483648;
#10;x=-1239483648;
#10;x=-1238483648;
#10;x=-1237483648;
#10;x=-1236483648;
#10;x=-1235483648;
#10;x=-1234483648;
#10;x=-1233483648;
#10;x=-1232483648;
#10;x=-1231483648;
#10;x=-1230483648;
#10;x=-1229483648;
#10;x=-1228483648;
#10;x=-1227483648;
#10;x=-1226483648;
#10;x=-1225483648;
#10;x=-1224483648;
#10;x=-1223483648;
#10;x=-1222483648;
#10;x=-1221483648;
#10;x=-1220483648;
#10;x=-1219483648;
#10;x=-1218483648;
#10;x=-1217483648;
#10;x=-1216483648;
#10;x=-1215483648;
#10;x=-1214483648;
#10;x=-1213483648;
#10;x=-1212483648;
#10;x=-1211483648;
#10;x=-1210483648;
#10;x=-1209483648;
#10;x=-1208483648;
#10;x=-1207483648;
#10;x=-1206483648;
#10;x=-1205483648;
#10;x=-1204483648;
#10;x=-1203483648;
#10;x=-1202483648;
#10;x=-1201483648;
#10;x=-1200483648;
#10;x=-1199483648;
#10;x=-1198483648;
#10;x=-1197483648;
#10;x=-1196483648;
#10;x=-1195483648;
#10;x=-1194483648;
#10;x=-1193483648;
#10;x=-1192483648;
#10;x=-1191483648;
#10;x=-1190483648;
#10;x=-1189483648;
#10;x=-1188483648;
#10;x=-1187483648;
#10;x=-1186483648;
#10;x=-1185483648;
#10;x=-1184483648;
#10;x=-1183483648;
#10;x=-1182483648;
#10;x=-1181483648;
#10;x=-1180483648;
#10;x=-1179483648;
#10;x=-1178483648;
#10;x=-1177483648;
#10;x=-1176483648;
#10;x=-1175483648;
#10;x=-1174483648;
#10;x=-1173483648;
#10;x=-1172483648;
#10;x=-1171483648;
#10;x=-1170483648;
#10;x=-1169483648;
#10;x=-1168483648;
#10;x=-1167483648;
#10;x=-1166483648;
#10;x=-1165483648;
#10;x=-1164483648;
#10;x=-1163483648;
#10;x=-1162483648;
#10;x=-1161483648;
#10;x=-1160483648;
#10;x=-1159483648;
#10;x=-1158483648;
#10;x=-1157483648;
#10;x=-1156483648;
#10;x=-1155483648;
#10;x=-1154483648;
#10;x=-1153483648;
#10;x=-1152483648;
#10;x=-1151483648;
#10;x=-1150483648;
#10;x=-1149483648;
#10;x=-1148483648;
#10;x=-1147483648;
#10;x=-1146483648;
#10;x=-1145483648;
#10;x=-1144483648;
#10;x=-1143483648;
#10;x=-1142483648;
#10;x=-1141483648;
#10;x=-1140483648;
#10;x=-1139483648;
#10;x=-1138483648;
#10;x=-1137483648;
#10;x=-1136483648;
#10;x=-1135483648;
#10;x=-1134483648;
#10;x=-1133483648;
#10;x=-1132483648;
#10;x=-1131483648;
#10;x=-1130483648;
#10;x=-1129483648;
#10;x=-1128483648;
#10;x=-1127483648;
#10;x=-1126483648;
#10;x=-1125483648;
#10;x=-1124483648;
#10;x=-1123483648;
#10;x=-1122483648;
#10;x=-1121483648;
#10;x=-1120483648;
#10;x=-1119483648;
#10;x=-1118483648;
#10;x=-1117483648;
#10;x=-1116483648;
#10;x=-1115483648;
#10;x=-1114483648;
#10;x=-1113483648;
#10;x=-1112483648;
#10;x=-1111483648;
#10;x=-1110483648;
#10;x=-1109483648;
#10;x=-1108483648;
#10;x=-1107483648;
#10;x=-1106483648;
#10;x=-1105483648;
#10;x=-1104483648;
#10;x=-1103483648;
#10;x=-1102483648;
#10;x=-1101483648;
#10;x=-1100483648;
#10;x=-1099483648;
#10;x=-1098483648;
#10;x=-1097483648;
#10;x=-1096483648;
#10;x=-1095483648;
#10;x=-1094483648;
#10;x=-1093483648;
#10;x=-1092483648;
#10;x=-1091483648;
#10;x=-1090483648;
#10;x=-1089483648;
#10;x=-1088483648;
#10;x=-1087483648;
#10;x=-1086483648;
#10;x=-1085483648;
#10;x=-1084483648;
#10;x=-1083483648;
#10;x=-1082483648;
#10;x=-1081483648;
#10;x=-1080483648;
#10;x=-1079483648;
#10;x=-1078483648;
#10;x=-1077483648;
#10;x=-1076483648;
#10;x=-1075483648;
#10;x=-1074483648;
#10;x=-1073483648;
#10;x=-1072483648;
#10;x=-1071483648;
#10;x=-1070483648;
#10;x=-1069483648;
#10;x=-1068483648;
#10;x=-1067483648;
#10;x=-1066483648;
#10;x=-1065483648;
#10;x=-1064483648;
#10;x=-1063483648;
#10;x=-1062483648;
#10;x=-1061483648;
#10;x=-1060483648;
#10;x=-1059483648;
#10;x=-1058483648;
#10;x=-1057483648;
#10;x=-1056483648;
#10;x=-1055483648;
#10;x=-1054483648;
#10;x=-1053483648;
#10;x=-1052483648;
#10;x=-1051483648;
#10;x=-1050483648;
#10;x=-1049483648;
#10;x=-1048483648;
#10;x=-1047483648;
#10;x=-1046483648;
#10;x=-1045483648;
#10;x=-1044483648;
#10;x=-1043483648;
#10;x=-1042483648;
#10;x=-1041483648;
#10;x=-1040483648;
#10;x=-1039483648;
#10;x=-1038483648;
#10;x=-1037483648;
#10;x=-1036483648;
#10;x=-1035483648;
#10;x=-1034483648;
#10;x=-1033483648;
#10;x=-1032483648;
#10;x=-1031483648;
#10;x=-1030483648;
#10;x=-1029483648;
#10;x=-1028483648;
#10;x=-1027483648;
#10;x=-1026483648;
#10;x=-1025483648;
#10;x=-1024483648;
#10;x=-1023483648;
#10;x=-1022483648;
#10;x=-1021483648;
#10;x=-1020483648;
#10;x=-1019483648;
#10;x=-1018483648;
#10;x=-1017483648;
#10;x=-1016483648;
#10;x=-1015483648;
#10;x=-1014483648;
#10;x=-1013483648;
#10;x=-1012483648;
#10;x=-1011483648;
#10;x=-1010483648;
#10;x=-1009483648;
#10;x=-1008483648;
#10;x=-1007483648;
#10;x=-1006483648;
#10;x=-1005483648;
#10;x=-1004483648;
#10;x=-1003483648;
#10;x=-1002483648;
#10;x=-1001483648;
#10;x=-1000483648;
#10;x=-999483648;
#10;x=-999383648;
#10;x=-999283648;
#10;x=-999183648;
#10;x=-999083648;
#10;x=-998983648;
#10;x=-998883648;
#10;x=-998783648;
#10;x=-998683648;
#10;x=-998583648;
#10;x=-998483648;
#10;x=-998383648;
#10;x=-998283648;
#10;x=-998183648;
#10;x=-998083648;
#10;x=-997983648;
#10;x=-997883648;
#10;x=-997783648;
#10;x=-997683648;
#10;x=-997583648;
#10;x=-997483648;
#10;x=-997383648;
#10;x=-997283648;
#10;x=-997183648;
#10;x=-997083648;
#10;x=-996983648;
#10;x=-996883648;
#10;x=-996783648;
#10;x=-996683648;
#10;x=-996583648;
#10;x=-996483648;
#10;x=-996383648;
#10;x=-996283648;
#10;x=-996183648;
#10;x=-996083648;
#10;x=-995983648;
#10;x=-995883648;
#10;x=-995783648;
#10;x=-995683648;
#10;x=-995583648;
#10;x=-995483648;
#10;x=-995383648;
#10;x=-995283648;
#10;x=-995183648;
#10;x=-995083648;
#10;x=-994983648;
#10;x=-994883648;
#10;x=-994783648;
#10;x=-994683648;
#10;x=-994583648;
#10;x=-994483648;
#10;x=-994383648;
#10;x=-994283648;
#10;x=-994183648;
#10;x=-994083648;
#10;x=-993983648;
#10;x=-993883648;
#10;x=-993783648;
#10;x=-993683648;
#10;x=-993583648;
#10;x=-993483648;
#10;x=-993383648;
#10;x=-993283648;
#10;x=-993183648;
#10;x=-993083648;
#10;x=-992983648;
#10;x=-992883648;
#10;x=-992783648;
#10;x=-992683648;
#10;x=-992583648;
#10;x=-992483648;
#10;x=-992383648;
#10;x=-992283648;
#10;x=-992183648;
#10;x=-992083648;
#10;x=-991983648;
#10;x=-991883648;
#10;x=-991783648;
#10;x=-991683648;
#10;x=-991583648;
#10;x=-991483648;
#10;x=-991383648;
#10;x=-991283648;
#10;x=-991183648;
#10;x=-991083648;
#10;x=-990983648;
#10;x=-990883648;
#10;x=-990783648;
#10;x=-990683648;
#10;x=-990583648;
#10;x=-990483648;
#10;x=-990383648;
#10;x=-990283648;
#10;x=-990183648;
#10;x=-990083648;
#10;x=-989983648;
#10;x=-989883648;
#10;x=-989783648;
#10;x=-989683648;
#10;x=-989583648;
#10;x=-989483648;
#10;x=-989383648;
#10;x=-989283648;
#10;x=-989183648;
#10;x=-989083648;
#10;x=-988983648;
#10;x=-988883648;
#10;x=-988783648;
#10;x=-988683648;
#10;x=-988583648;
#10;x=-988483648;
#10;x=-988383648;
#10;x=-988283648;
#10;x=-988183648;
#10;x=-988083648;
#10;x=-987983648;
#10;x=-987883648;
#10;x=-987783648;
#10;x=-987683648;
#10;x=-987583648;
#10;x=-987483648;
#10;x=-987383648;
#10;x=-987283648;
#10;x=-987183648;
#10;x=-987083648;
#10;x=-986983648;
#10;x=-986883648;
#10;x=-986783648;
#10;x=-986683648;
#10;x=-986583648;
#10;x=-986483648;
#10;x=-986383648;
#10;x=-986283648;
#10;x=-986183648;
#10;x=-986083648;
#10;x=-985983648;
#10;x=-985883648;
#10;x=-985783648;
#10;x=-985683648;
#10;x=-985583648;
#10;x=-985483648;
#10;x=-985383648;
#10;x=-985283648;
#10;x=-985183648;
#10;x=-985083648;
#10;x=-984983648;
#10;x=-984883648;
#10;x=-984783648;
#10;x=-984683648;
#10;x=-984583648;
#10;x=-984483648;
#10;x=-984383648;
#10;x=-984283648;
#10;x=-984183648;
#10;x=-984083648;
#10;x=-983983648;
#10;x=-983883648;
#10;x=-983783648;
#10;x=-983683648;
#10;x=-983583648;
#10;x=-983483648;
#10;x=-983383648;
#10;x=-983283648;
#10;x=-983183648;
#10;x=-983083648;
#10;x=-982983648;
#10;x=-982883648;
#10;x=-982783648;
#10;x=-982683648;
#10;x=-982583648;
#10;x=-982483648;
#10;x=-982383648;
#10;x=-982283648;
#10;x=-982183648;
#10;x=-982083648;
#10;x=-981983648;
#10;x=-981883648;
#10;x=-981783648;
#10;x=-981683648;
#10;x=-981583648;
#10;x=-981483648;
#10;x=-981383648;
#10;x=-981283648;
#10;x=-981183648;
#10;x=-981083648;
#10;x=-980983648;
#10;x=-980883648;
#10;x=-980783648;
#10;x=-980683648;
#10;x=-980583648;
#10;x=-980483648;
#10;x=-980383648;
#10;x=-980283648;
#10;x=-980183648;
#10;x=-980083648;
#10;x=-979983648;
#10;x=-979883648;
#10;x=-979783648;
#10;x=-979683648;
#10;x=-979583648;
#10;x=-979483648;
#10;x=-979383648;
#10;x=-979283648;
#10;x=-979183648;
#10;x=-979083648;
#10;x=-978983648;
#10;x=-978883648;
#10;x=-978783648;
#10;x=-978683648;
#10;x=-978583648;
#10;x=-978483648;
#10;x=-978383648;
#10;x=-978283648;
#10;x=-978183648;
#10;x=-978083648;
#10;x=-977983648;
#10;x=-977883648;
#10;x=-977783648;
#10;x=-977683648;
#10;x=-977583648;
#10;x=-977483648;
#10;x=-977383648;
#10;x=-977283648;
#10;x=-977183648;
#10;x=-977083648;
#10;x=-976983648;
#10;x=-976883648;
#10;x=-976783648;
#10;x=-976683648;
#10;x=-976583648;
#10;x=-976483648;
#10;x=-976383648;
#10;x=-976283648;
#10;x=-976183648;
#10;x=-976083648;
#10;x=-975983648;
#10;x=-975883648;
#10;x=-975783648;
#10;x=-975683648;
#10;x=-975583648;
#10;x=-975483648;
#10;x=-975383648;
#10;x=-975283648;
#10;x=-975183648;
#10;x=-975083648;
#10;x=-974983648;
#10;x=-974883648;
#10;x=-974783648;
#10;x=-974683648;
#10;x=-974583648;
#10;x=-974483648;
#10;x=-974383648;
#10;x=-974283648;
#10;x=-974183648;
#10;x=-974083648;
#10;x=-973983648;
#10;x=-973883648;
#10;x=-973783648;
#10;x=-973683648;
#10;x=-973583648;
#10;x=-973483648;
#10;x=-973383648;
#10;x=-973283648;
#10;x=-973183648;
#10;x=-973083648;
#10;x=-972983648;
#10;x=-972883648;
#10;x=-972783648;
#10;x=-972683648;
#10;x=-972583648;
#10;x=-972483648;
#10;x=-972383648;
#10;x=-972283648;
#10;x=-972183648;
#10;x=-972083648;
#10;x=-971983648;
#10;x=-971883648;
#10;x=-971783648;
#10;x=-971683648;
#10;x=-971583648;
#10;x=-971483648;
#10;x=-971383648;
#10;x=-971283648;
#10;x=-971183648;
#10;x=-971083648;
#10;x=-970983648;
#10;x=-970883648;
#10;x=-970783648;
#10;x=-970683648;
#10;x=-970583648;
#10;x=-970483648;
#10;x=-970383648;
#10;x=-970283648;
#10;x=-970183648;
#10;x=-970083648;
#10;x=-969983648;
#10;x=-969883648;
#10;x=-969783648;
#10;x=-969683648;
#10;x=-969583648;
#10;x=-969483648;
#10;x=-969383648;
#10;x=-969283648;
#10;x=-969183648;
#10;x=-969083648;
#10;x=-968983648;
#10;x=-968883648;
#10;x=-968783648;
#10;x=-968683648;
#10;x=-968583648;
#10;x=-968483648;
#10;x=-968383648;
#10;x=-968283648;
#10;x=-968183648;
#10;x=-968083648;
#10;x=-967983648;
#10;x=-967883648;
#10;x=-967783648;
#10;x=-967683648;
#10;x=-967583648;
#10;x=-967483648;
#10;x=-967383648;
#10;x=-967283648;
#10;x=-967183648;
#10;x=-967083648;
#10;x=-966983648;
#10;x=-966883648;
#10;x=-966783648;
#10;x=-966683648;
#10;x=-966583648;
#10;x=-966483648;
#10;x=-966383648;
#10;x=-966283648;
#10;x=-966183648;
#10;x=-966083648;
#10;x=-965983648;
#10;x=-965883648;
#10;x=-965783648;
#10;x=-965683648;
#10;x=-965583648;
#10;x=-965483648;
#10;x=-965383648;
#10;x=-965283648;
#10;x=-965183648;
#10;x=-965083648;
#10;x=-964983648;
#10;x=-964883648;
#10;x=-964783648;
#10;x=-964683648;
#10;x=-964583648;
#10;x=-964483648;
#10;x=-964383648;
#10;x=-964283648;
#10;x=-964183648;
#10;x=-964083648;
#10;x=-963983648;
#10;x=-963883648;
#10;x=-963783648;
#10;x=-963683648;
#10;x=-963583648;
#10;x=-963483648;
#10;x=-963383648;
#10;x=-963283648;
#10;x=-963183648;
#10;x=-963083648;
#10;x=-962983648;
#10;x=-962883648;
#10;x=-962783648;
#10;x=-962683648;
#10;x=-962583648;
#10;x=-962483648;
#10;x=-962383648;
#10;x=-962283648;
#10;x=-962183648;
#10;x=-962083648;
#10;x=-961983648;
#10;x=-961883648;
#10;x=-961783648;
#10;x=-961683648;
#10;x=-961583648;
#10;x=-961483648;
#10;x=-961383648;
#10;x=-961283648;
#10;x=-961183648;
#10;x=-961083648;
#10;x=-960983648;
#10;x=-960883648;
#10;x=-960783648;
#10;x=-960683648;
#10;x=-960583648;
#10;x=-960483648;
#10;x=-960383648;
#10;x=-960283648;
#10;x=-960183648;
#10;x=-960083648;
#10;x=-959983648;
#10;x=-959883648;
#10;x=-959783648;
#10;x=-959683648;
#10;x=-959583648;
#10;x=-959483648;
#10;x=-959383648;
#10;x=-959283648;
#10;x=-959183648;
#10;x=-959083648;
#10;x=-958983648;
#10;x=-958883648;
#10;x=-958783648;
#10;x=-958683648;
#10;x=-958583648;
#10;x=-958483648;
#10;x=-958383648;
#10;x=-958283648;
#10;x=-958183648;
#10;x=-958083648;
#10;x=-957983648;
#10;x=-957883648;
#10;x=-957783648;
#10;x=-957683648;
#10;x=-957583648;
#10;x=-957483648;
#10;x=-957383648;
#10;x=-957283648;
#10;x=-957183648;
#10;x=-957083648;
#10;x=-956983648;
#10;x=-956883648;
#10;x=-956783648;
#10;x=-956683648;
#10;x=-956583648;
#10;x=-956483648;
#10;x=-956383648;
#10;x=-956283648;
#10;x=-956183648;
#10;x=-956083648;
#10;x=-955983648;
#10;x=-955883648;
#10;x=-955783648;
#10;x=-955683648;
#10;x=-955583648;
#10;x=-955483648;
#10;x=-955383648;
#10;x=-955283648;
#10;x=-955183648;
#10;x=-955083648;
#10;x=-954983648;
#10;x=-954883648;
#10;x=-954783648;
#10;x=-954683648;
#10;x=-954583648;
#10;x=-954483648;
#10;x=-954383648;
#10;x=-954283648;
#10;x=-954183648;
#10;x=-954083648;
#10;x=-953983648;
#10;x=-953883648;
#10;x=-953783648;
#10;x=-953683648;
#10;x=-953583648;
#10;x=-953483648;
#10;x=-953383648;
#10;x=-953283648;
#10;x=-953183648;
#10;x=-953083648;
#10;x=-952983648;
#10;x=-952883648;
#10;x=-952783648;
#10;x=-952683648;
#10;x=-952583648;
#10;x=-952483648;
#10;x=-952383648;
#10;x=-952283648;
#10;x=-952183648;
#10;x=-952083648;
#10;x=-951983648;
#10;x=-951883648;
#10;x=-951783648;
#10;x=-951683648;
#10;x=-951583648;
#10;x=-951483648;
#10;x=-951383648;
#10;x=-951283648;
#10;x=-951183648;
#10;x=-951083648;
#10;x=-950983648;
#10;x=-950883648;
#10;x=-950783648;
#10;x=-950683648;
#10;x=-950583648;
#10;x=-950483648;
#10;x=-950383648;
#10;x=-950283648;
#10;x=-950183648;
#10;x=-950083648;
#10;x=-949983648;
#10;x=-949883648;
#10;x=-949783648;
#10;x=-949683648;
#10;x=-949583648;
#10;x=-949483648;
#10;x=-949383648;
#10;x=-949283648;
#10;x=-949183648;
#10;x=-949083648;
#10;x=-948983648;
#10;x=-948883648;
#10;x=-948783648;
#10;x=-948683648;
#10;x=-948583648;
#10;x=-948483648;
#10;x=-948383648;
#10;x=-948283648;
#10;x=-948183648;
#10;x=-948083648;
#10;x=-947983648;
#10;x=-947883648;
#10;x=-947783648;
#10;x=-947683648;
#10;x=-947583648;
#10;x=-947483648;
#10;x=-947383648;
#10;x=-947283648;
#10;x=-947183648;
#10;x=-947083648;
#10;x=-946983648;
#10;x=-946883648;
#10;x=-946783648;
#10;x=-946683648;
#10;x=-946583648;
#10;x=-946483648;
#10;x=-946383648;
#10;x=-946283648;
#10;x=-946183648;
#10;x=-946083648;
#10;x=-945983648;
#10;x=-945883648;
#10;x=-945783648;
#10;x=-945683648;
#10;x=-945583648;
#10;x=-945483648;
#10;x=-945383648;
#10;x=-945283648;
#10;x=-945183648;
#10;x=-945083648;
#10;x=-944983648;
#10;x=-944883648;
#10;x=-944783648;
#10;x=-944683648;
#10;x=-944583648;
#10;x=-944483648;
#10;x=-944383648;
#10;x=-944283648;
#10;x=-944183648;
#10;x=-944083648;
#10;x=-943983648;
#10;x=-943883648;
#10;x=-943783648;
#10;x=-943683648;
#10;x=-943583648;
#10;x=-943483648;
#10;x=-943383648;
#10;x=-943283648;
#10;x=-943183648;
#10;x=-943083648;
#10;x=-942983648;
#10;x=-942883648;
#10;x=-942783648;
#10;x=-942683648;
#10;x=-942583648;
#10;x=-942483648;
#10;x=-942383648;
#10;x=-942283648;
#10;x=-942183648;
#10;x=-942083648;
#10;x=-941983648;
#10;x=-941883648;
#10;x=-941783648;
#10;x=-941683648;
#10;x=-941583648;
#10;x=-941483648;
#10;x=-941383648;
#10;x=-941283648;
#10;x=-941183648;
#10;x=-941083648;
#10;x=-940983648;
#10;x=-940883648;
#10;x=-940783648;
#10;x=-940683648;
#10;x=-940583648;
#10;x=-940483648;
#10;x=-940383648;
#10;x=-940283648;
#10;x=-940183648;
#10;x=-940083648;
#10;x=-939983648;
#10;x=-939883648;
#10;x=-939783648;
#10;x=-939683648;
#10;x=-939583648;
#10;x=-939483648;
#10;x=-939383648;
#10;x=-939283648;
#10;x=-939183648;
#10;x=-939083648;
#10;x=-938983648;
#10;x=-938883648;
#10;x=-938783648;
#10;x=-938683648;
#10;x=-938583648;
#10;x=-938483648;
#10;x=-938383648;
#10;x=-938283648;
#10;x=-938183648;
#10;x=-938083648;
#10;x=-937983648;
#10;x=-937883648;
#10;x=-937783648;
#10;x=-937683648;
#10;x=-937583648;
#10;x=-937483648;
#10;x=-937383648;
#10;x=-937283648;
#10;x=-937183648;
#10;x=-937083648;
#10;x=-936983648;
#10;x=-936883648;
#10;x=-936783648;
#10;x=-936683648;
#10;x=-936583648;
#10;x=-936483648;
#10;x=-936383648;
#10;x=-936283648;
#10;x=-936183648;
#10;x=-936083648;
#10;x=-935983648;
#10;x=-935883648;
#10;x=-935783648;
#10;x=-935683648;
#10;x=-935583648;
#10;x=-935483648;
#10;x=-935383648;
#10;x=-935283648;
#10;x=-935183648;
#10;x=-935083648;
#10;x=-934983648;
#10;x=-934883648;
#10;x=-934783648;
#10;x=-934683648;
#10;x=-934583648;
#10;x=-934483648;
#10;x=-934383648;
#10;x=-934283648;
#10;x=-934183648;
#10;x=-934083648;
#10;x=-933983648;
#10;x=-933883648;
#10;x=-933783648;
#10;x=-933683648;
#10;x=-933583648;
#10;x=-933483648;
#10;x=-933383648;
#10;x=-933283648;
#10;x=-933183648;
#10;x=-933083648;
#10;x=-932983648;
#10;x=-932883648;
#10;x=-932783648;
#10;x=-932683648;
#10;x=-932583648;
#10;x=-932483648;
#10;x=-932383648;
#10;x=-932283648;
#10;x=-932183648;
#10;x=-932083648;
#10;x=-931983648;
#10;x=-931883648;
#10;x=-931783648;
#10;x=-931683648;
#10;x=-931583648;
#10;x=-931483648;
#10;x=-931383648;
#10;x=-931283648;
#10;x=-931183648;
#10;x=-931083648;
#10;x=-930983648;
#10;x=-930883648;
#10;x=-930783648;
#10;x=-930683648;
#10;x=-930583648;
#10;x=-930483648;
#10;x=-930383648;
#10;x=-930283648;
#10;x=-930183648;
#10;x=-930083648;
#10;x=-929983648;
#10;x=-929883648;
#10;x=-929783648;
#10;x=-929683648;
#10;x=-929583648;
#10;x=-929483648;
#10;x=-929383648;
#10;x=-929283648;
#10;x=-929183648;
#10;x=-929083648;
#10;x=-928983648;
#10;x=-928883648;
#10;x=-928783648;
#10;x=-928683648;
#10;x=-928583648;
#10;x=-928483648;
#10;x=-928383648;
#10;x=-928283648;
#10;x=-928183648;
#10;x=-928083648;
#10;x=-927983648;
#10;x=-927883648;
#10;x=-927783648;
#10;x=-927683648;
#10;x=-927583648;
#10;x=-927483648;
#10;x=-927383648;
#10;x=-927283648;
#10;x=-927183648;
#10;x=-927083648;
#10;x=-926983648;
#10;x=-926883648;
#10;x=-926783648;
#10;x=-926683648;
#10;x=-926583648;
#10;x=-926483648;
#10;x=-926383648;
#10;x=-926283648;
#10;x=-926183648;
#10;x=-926083648;
#10;x=-925983648;
#10;x=-925883648;
#10;x=-925783648;
#10;x=-925683648;
#10;x=-925583648;
#10;x=-925483648;
#10;x=-925383648;
#10;x=-925283648;
#10;x=-925183648;
#10;x=-925083648;
#10;x=-924983648;
#10;x=-924883648;
#10;x=-924783648;
#10;x=-924683648;
#10;x=-924583648;
#10;x=-924483648;
#10;x=-924383648;
#10;x=-924283648;
#10;x=-924183648;
#10;x=-924083648;
#10;x=-923983648;
#10;x=-923883648;
#10;x=-923783648;
#10;x=-923683648;
#10;x=-923583648;
#10;x=-923483648;
#10;x=-923383648;
#10;x=-923283648;
#10;x=-923183648;
#10;x=-923083648;
#10;x=-922983648;
#10;x=-922883648;
#10;x=-922783648;
#10;x=-922683648;
#10;x=-922583648;
#10;x=-922483648;
#10;x=-922383648;
#10;x=-922283648;
#10;x=-922183648;
#10;x=-922083648;
#10;x=-921983648;
#10;x=-921883648;
#10;x=-921783648;
#10;x=-921683648;
#10;x=-921583648;
#10;x=-921483648;
#10;x=-921383648;
#10;x=-921283648;
#10;x=-921183648;
#10;x=-921083648;
#10;x=-920983648;
#10;x=-920883648;
#10;x=-920783648;
#10;x=-920683648;
#10;x=-920583648;
#10;x=-920483648;
#10;x=-920383648;
#10;x=-920283648;
#10;x=-920183648;
#10;x=-920083648;
#10;x=-919983648;
#10;x=-919883648;
#10;x=-919783648;
#10;x=-919683648;
#10;x=-919583648;
#10;x=-919483648;
#10;x=-919383648;
#10;x=-919283648;
#10;x=-919183648;
#10;x=-919083648;
#10;x=-918983648;
#10;x=-918883648;
#10;x=-918783648;
#10;x=-918683648;
#10;x=-918583648;
#10;x=-918483648;
#10;x=-918383648;
#10;x=-918283648;
#10;x=-918183648;
#10;x=-918083648;
#10;x=-917983648;
#10;x=-917883648;
#10;x=-917783648;
#10;x=-917683648;
#10;x=-917583648;
#10;x=-917483648;
#10;x=-917383648;
#10;x=-917283648;
#10;x=-917183648;
#10;x=-917083648;
#10;x=-916983648;
#10;x=-916883648;
#10;x=-916783648;
#10;x=-916683648;
#10;x=-916583648;
#10;x=-916483648;
#10;x=-916383648;
#10;x=-916283648;
#10;x=-916183648;
#10;x=-916083648;
#10;x=-915983648;
#10;x=-915883648;
#10;x=-915783648;
#10;x=-915683648;
#10;x=-915583648;
#10;x=-915483648;
#10;x=-915383648;
#10;x=-915283648;
#10;x=-915183648;
#10;x=-915083648;
#10;x=-914983648;
#10;x=-914883648;
#10;x=-914783648;
#10;x=-914683648;
#10;x=-914583648;
#10;x=-914483648;
#10;x=-914383648;
#10;x=-914283648;
#10;x=-914183648;
#10;x=-914083648;
#10;x=-913983648;
#10;x=-913883648;
#10;x=-913783648;
#10;x=-913683648;
#10;x=-913583648;
#10;x=-913483648;
#10;x=-913383648;
#10;x=-913283648;
#10;x=-913183648;
#10;x=-913083648;
#10;x=-912983648;
#10;x=-912883648;
#10;x=-912783648;
#10;x=-912683648;
#10;x=-912583648;
#10;x=-912483648;
#10;x=-912383648;
#10;x=-912283648;
#10;x=-912183648;
#10;x=-912083648;
#10;x=-911983648;
#10;x=-911883648;
#10;x=-911783648;
#10;x=-911683648;
#10;x=-911583648;
#10;x=-911483648;
#10;x=-911383648;
#10;x=-911283648;
#10;x=-911183648;
#10;x=-911083648;
#10;x=-910983648;
#10;x=-910883648;
#10;x=-910783648;
#10;x=-910683648;
#10;x=-910583648;
#10;x=-910483648;
#10;x=-910383648;
#10;x=-910283648;
#10;x=-910183648;
#10;x=-910083648;
#10;x=-909983648;
#10;x=-909883648;
#10;x=-909783648;
#10;x=-909683648;
#10;x=-909583648;
#10;x=-909483648;
#10;x=-909383648;
#10;x=-909283648;
#10;x=-909183648;
#10;x=-909083648;
#10;x=-908983648;
#10;x=-908883648;
#10;x=-908783648;
#10;x=-908683648;
#10;x=-908583648;
#10;x=-908483648;
#10;x=-908383648;
#10;x=-908283648;
#10;x=-908183648;
#10;x=-908083648;
#10;x=-907983648;
#10;x=-907883648;
#10;x=-907783648;
#10;x=-907683648;
#10;x=-907583648;
#10;x=-907483648;
#10;x=-907383648;
#10;x=-907283648;
#10;x=-907183648;
#10;x=-907083648;
#10;x=-906983648;
#10;x=-906883648;
#10;x=-906783648;
#10;x=-906683648;
#10;x=-906583648;
#10;x=-906483648;
#10;x=-906383648;
#10;x=-906283648;
#10;x=-906183648;
#10;x=-906083648;
#10;x=-905983648;
#10;x=-905883648;
#10;x=-905783648;
#10;x=-905683648;
#10;x=-905583648;
#10;x=-905483648;
#10;x=-905383648;
#10;x=-905283648;
#10;x=-905183648;
#10;x=-905083648;
#10;x=-904983648;
#10;x=-904883648;
#10;x=-904783648;
#10;x=-904683648;
#10;x=-904583648;
#10;x=-904483648;
#10;x=-904383648;
#10;x=-904283648;
#10;x=-904183648;
#10;x=-904083648;
#10;x=-903983648;
#10;x=-903883648;
#10;x=-903783648;
#10;x=-903683648;
#10;x=-903583648;
#10;x=-903483648;
#10;x=-903383648;
#10;x=-903283648;
#10;x=-903183648;
#10;x=-903083648;
#10;x=-902983648;
#10;x=-902883648;
#10;x=-902783648;
#10;x=-902683648;
#10;x=-902583648;
#10;x=-902483648;
#10;x=-902383648;
#10;x=-902283648;
#10;x=-902183648;
#10;x=-902083648;
#10;x=-901983648;
#10;x=-901883648;
#10;x=-901783648;
#10;x=-901683648;
#10;x=-901583648;
#10;x=-901483648;
#10;x=-901383648;
#10;x=-901283648;
#10;x=-901183648;
#10;x=-901083648;
#10;x=-900983648;
#10;x=-900883648;
#10;x=-900783648;
#10;x=-900683648;
#10;x=-900583648;
#10;x=-900483648;
#10;x=-900383648;
#10;x=-900283648;
#10;x=-900183648;
#10;x=-900083648;
#10;x=-899983648;
#10;x=-899883648;
#10;x=-899783648;
#10;x=-899683648;
#10;x=-899583648;
#10;x=-899483648;
#10;x=-899383648;
#10;x=-899283648;
#10;x=-899183648;
#10;x=-899083648;
#10;x=-898983648;
#10;x=-898883648;
#10;x=-898783648;
#10;x=-898683648;
#10;x=-898583648;
#10;x=-898483648;
#10;x=-898383648;
#10;x=-898283648;
#10;x=-898183648;
#10;x=-898083648;
#10;x=-897983648;
#10;x=-897883648;
#10;x=-897783648;
#10;x=-897683648;
#10;x=-897583648;
#10;x=-897483648;
#10;x=-897383648;
#10;x=-897283648;
#10;x=-897183648;
#10;x=-897083648;
#10;x=-896983648;
#10;x=-896883648;
#10;x=-896783648;
#10;x=-896683648;
#10;x=-896583648;
#10;x=-896483648;
#10;x=-896383648;
#10;x=-896283648;
#10;x=-896183648;
#10;x=-896083648;
#10;x=-895983648;
#10;x=-895883648;
#10;x=-895783648;
#10;x=-895683648;
#10;x=-895583648;
#10;x=-895483648;
#10;x=-895383648;
#10;x=-895283648;
#10;x=-895183648;
#10;x=-895083648;
#10;x=-894983648;
#10;x=-894883648;
#10;x=-894783648;
#10;x=-894683648;
#10;x=-894583648;
#10;x=-894483648;
#10;x=-894383648;
#10;x=-894283648;
#10;x=-894183648;
#10;x=-894083648;
#10;x=-893983648;
#10;x=-893883648;
#10;x=-893783648;
#10;x=-893683648;
#10;x=-893583648;
#10;x=-893483648;
#10;x=-893383648;
#10;x=-893283648;
#10;x=-893183648;
#10;x=-893083648;
#10;x=-892983648;
#10;x=-892883648;
#10;x=-892783648;
#10;x=-892683648;
#10;x=-892583648;
#10;x=-892483648;
#10;x=-892383648;
#10;x=-892283648;
#10;x=-892183648;
#10;x=-892083648;
#10;x=-891983648;
#10;x=-891883648;
#10;x=-891783648;
#10;x=-891683648;
#10;x=-891583648;
#10;x=-891483648;
#10;x=-891383648;
#10;x=-891283648;
#10;x=-891183648;
#10;x=-891083648;
#10;x=-890983648;
#10;x=-890883648;
#10;x=-890783648;
#10;x=-890683648;
#10;x=-890583648;
#10;x=-890483648;
#10;x=-890383648;
#10;x=-890283648;
#10;x=-890183648;
#10;x=-890083648;
#10;x=-889983648;
#10;x=-889883648;
#10;x=-889783648;
#10;x=-889683648;
#10;x=-889583648;
#10;x=-889483648;
#10;x=-889383648;
#10;x=-889283648;
#10;x=-889183648;
#10;x=-889083648;
#10;x=-888983648;
#10;x=-888883648;
#10;x=-888783648;
#10;x=-888683648;
#10;x=-888583648;
#10;x=-888483648;
#10;x=-888383648;
#10;x=-888283648;
#10;x=-888183648;
#10;x=-888083648;
#10;x=-887983648;
#10;x=-887883648;
#10;x=-887783648;
#10;x=-887683648;
#10;x=-887583648;
#10;x=-887483648;
#10;x=-887383648;
#10;x=-887283648;
#10;x=-887183648;
#10;x=-887083648;
#10;x=-886983648;
#10;x=-886883648;
#10;x=-886783648;
#10;x=-886683648;
#10;x=-886583648;
#10;x=-886483648;
#10;x=-886383648;
#10;x=-886283648;
#10;x=-886183648;
#10;x=-886083648;
#10;x=-885983648;
#10;x=-885883648;
#10;x=-885783648;
#10;x=-885683648;
#10;x=-885583648;
#10;x=-885483648;
#10;x=-885383648;
#10;x=-885283648;
#10;x=-885183648;
#10;x=-885083648;
#10;x=-884983648;
#10;x=-884883648;
#10;x=-884783648;
#10;x=-884683648;
#10;x=-884583648;
#10;x=-884483648;
#10;x=-884383648;
#10;x=-884283648;
#10;x=-884183648;
#10;x=-884083648;
#10;x=-883983648;
#10;x=-883883648;
#10;x=-883783648;
#10;x=-883683648;
#10;x=-883583648;
#10;x=-883483648;
#10;x=-883383648;
#10;x=-883283648;
#10;x=-883183648;
#10;x=-883083648;
#10;x=-882983648;
#10;x=-882883648;
#10;x=-882783648;
#10;x=-882683648;
#10;x=-882583648;
#10;x=-882483648;
#10;x=-882383648;
#10;x=-882283648;
#10;x=-882183648;
#10;x=-882083648;
#10;x=-881983648;
#10;x=-881883648;
#10;x=-881783648;
#10;x=-881683648;
#10;x=-881583648;
#10;x=-881483648;
#10;x=-881383648;
#10;x=-881283648;
#10;x=-881183648;
#10;x=-881083648;
#10;x=-880983648;
#10;x=-880883648;
#10;x=-880783648;
#10;x=-880683648;
#10;x=-880583648;
#10;x=-880483648;
#10;x=-880383648;
#10;x=-880283648;
#10;x=-880183648;
#10;x=-880083648;
#10;x=-879983648;
#10;x=-879883648;
#10;x=-879783648;
#10;x=-879683648;
#10;x=-879583648;
#10;x=-879483648;
#10;x=-879383648;
#10;x=-879283648;
#10;x=-879183648;
#10;x=-879083648;
#10;x=-878983648;
#10;x=-878883648;
#10;x=-878783648;
#10;x=-878683648;
#10;x=-878583648;
#10;x=-878483648;
#10;x=-878383648;
#10;x=-878283648;
#10;x=-878183648;
#10;x=-878083648;
#10;x=-877983648;
#10;x=-877883648;
#10;x=-877783648;
#10;x=-877683648;
#10;x=-877583648;
#10;x=-877483648;
#10;x=-877383648;
#10;x=-877283648;
#10;x=-877183648;
#10;x=-877083648;
#10;x=-876983648;
#10;x=-876883648;
#10;x=-876783648;
#10;x=-876683648;
#10;x=-876583648;
#10;x=-876483648;
#10;x=-876383648;
#10;x=-876283648;
#10;x=-876183648;
#10;x=-876083648;
#10;x=-875983648;
#10;x=-875883648;
#10;x=-875783648;
#10;x=-875683648;
#10;x=-875583648;
#10;x=-875483648;
#10;x=-875383648;
#10;x=-875283648;
#10;x=-875183648;
#10;x=-875083648;
#10;x=-874983648;
#10;x=-874883648;
#10;x=-874783648;
#10;x=-874683648;
#10;x=-874583648;
#10;x=-874483648;
#10;x=-874383648;
#10;x=-874283648;
#10;x=-874183648;
#10;x=-874083648;
#10;x=-873983648;
#10;x=-873883648;
#10;x=-873783648;
#10;x=-873683648;
#10;x=-873583648;
#10;x=-873483648;
#10;x=-873383648;
#10;x=-873283648;
#10;x=-873183648;
#10;x=-873083648;
#10;x=-872983648;
#10;x=-872883648;
#10;x=-872783648;
#10;x=-872683648;
#10;x=-872583648;
#10;x=-872483648;
#10;x=-872383648;
#10;x=-872283648;
#10;x=-872183648;
#10;x=-872083648;
#10;x=-871983648;
#10;x=-871883648;
#10;x=-871783648;
#10;x=-871683648;
#10;x=-871583648;
#10;x=-871483648;
#10;x=-871383648;
#10;x=-871283648;
#10;x=-871183648;
#10;x=-871083648;
#10;x=-870983648;
#10;x=-870883648;
#10;x=-870783648;
#10;x=-870683648;
#10;x=-870583648;
#10;x=-870483648;
#10;x=-870383648;
#10;x=-870283648;
#10;x=-870183648;
#10;x=-870083648;
#10;x=-869983648;
#10;x=-869883648;
#10;x=-869783648;
#10;x=-869683648;
#10;x=-869583648;
#10;x=-869483648;
#10;x=-869383648;
#10;x=-869283648;
#10;x=-869183648;
#10;x=-869083648;
#10;x=-868983648;
#10;x=-868883648;
#10;x=-868783648;
#10;x=-868683648;
#10;x=-868583648;
#10;x=-868483648;
#10;x=-868383648;
#10;x=-868283648;
#10;x=-868183648;
#10;x=-868083648;
#10;x=-867983648;
#10;x=-867883648;
#10;x=-867783648;
#10;x=-867683648;
#10;x=-867583648;
#10;x=-867483648;
#10;x=-867383648;
#10;x=-867283648;
#10;x=-867183648;
#10;x=-867083648;
#10;x=-866983648;
#10;x=-866883648;
#10;x=-866783648;
#10;x=-866683648;
#10;x=-866583648;
#10;x=-866483648;
#10;x=-866383648;
#10;x=-866283648;
#10;x=-866183648;
#10;x=-866083648;
#10;x=-865983648;
#10;x=-865883648;
#10;x=-865783648;
#10;x=-865683648;
#10;x=-865583648;
#10;x=-865483648;
#10;x=-865383648;
#10;x=-865283648;
#10;x=-865183648;
#10;x=-865083648;
#10;x=-864983648;
#10;x=-864883648;
#10;x=-864783648;
#10;x=-864683648;
#10;x=-864583648;
#10;x=-864483648;
#10;x=-864383648;
#10;x=-864283648;
#10;x=-864183648;
#10;x=-864083648;
#10;x=-863983648;
#10;x=-863883648;
#10;x=-863783648;
#10;x=-863683648;
#10;x=-863583648;
#10;x=-863483648;
#10;x=-863383648;
#10;x=-863283648;
#10;x=-863183648;
#10;x=-863083648;
#10;x=-862983648;
#10;x=-862883648;
#10;x=-862783648;
#10;x=-862683648;
#10;x=-862583648;
#10;x=-862483648;
#10;x=-862383648;
#10;x=-862283648;
#10;x=-862183648;
#10;x=-862083648;
#10;x=-861983648;
#10;x=-861883648;
#10;x=-861783648;
#10;x=-861683648;
#10;x=-861583648;
#10;x=-861483648;
#10;x=-861383648;
#10;x=-861283648;
#10;x=-861183648;
#10;x=-861083648;
#10;x=-860983648;
#10;x=-860883648;
#10;x=-860783648;
#10;x=-860683648;
#10;x=-860583648;
#10;x=-860483648;
#10;x=-860383648;
#10;x=-860283648;
#10;x=-860183648;
#10;x=-860083648;
#10;x=-859983648;
#10;x=-859883648;
#10;x=-859783648;
#10;x=-859683648;
#10;x=-859583648;
#10;x=-859483648;
#10;x=-859383648;
#10;x=-859283648;
#10;x=-859183648;
#10;x=-859083648;
#10;x=-858983648;
#10;x=-858883648;
#10;x=-858783648;
#10;x=-858683648;
#10;x=-858583648;
#10;x=-858483648;
#10;x=-858383648;
#10;x=-858283648;
#10;x=-858183648;
#10;x=-858083648;
#10;x=-857983648;
#10;x=-857883648;
#10;x=-857783648;
#10;x=-857683648;
#10;x=-857583648;
#10;x=-857483648;
#10;x=-857383648;
#10;x=-857283648;
#10;x=-857183648;
#10;x=-857083648;
#10;x=-856983648;
#10;x=-856883648;
#10;x=-856783648;
#10;x=-856683648;
#10;x=-856583648;
#10;x=-856483648;
#10;x=-856383648;
#10;x=-856283648;
#10;x=-856183648;
#10;x=-856083648;
#10;x=-855983648;
#10;x=-855883648;
#10;x=-855783648;
#10;x=-855683648;
#10;x=-855583648;
#10;x=-855483648;
#10;x=-855383648;
#10;x=-855283648;
#10;x=-855183648;
#10;x=-855083648;
#10;x=-854983648;
#10;x=-854883648;
#10;x=-854783648;
#10;x=-854683648;
#10;x=-854583648;
#10;x=-854483648;
#10;x=-854383648;
#10;x=-854283648;
#10;x=-854183648;
#10;x=-854083648;
#10;x=-853983648;
#10;x=-853883648;
#10;x=-853783648;
#10;x=-853683648;
#10;x=-853583648;
#10;x=-853483648;
#10;x=-853383648;
#10;x=-853283648;
#10;x=-853183648;
#10;x=-853083648;
#10;x=-852983648;
#10;x=-852883648;
#10;x=-852783648;
#10;x=-852683648;
#10;x=-852583648;
#10;x=-852483648;
#10;x=-852383648;
#10;x=-852283648;
#10;x=-852183648;
#10;x=-852083648;
#10;x=-851983648;
#10;x=-851883648;
#10;x=-851783648;
#10;x=-851683648;
#10;x=-851583648;
#10;x=-851483648;
#10;x=-851383648;
#10;x=-851283648;
#10;x=-851183648;
#10;x=-851083648;
#10;x=-850983648;
#10;x=-850883648;
#10;x=-850783648;
#10;x=-850683648;
#10;x=-850583648;
#10;x=-850483648;
#10;x=-850383648;
#10;x=-850283648;
#10;x=-850183648;
#10;x=-850083648;
#10;x=-849983648;
#10;x=-849883648;
#10;x=-849783648;
#10;x=-849683648;
#10;x=-849583648;
#10;x=-849483648;
#10;x=-849383648;
#10;x=-849283648;
#10;x=-849183648;
#10;x=-849083648;
#10;x=-848983648;
#10;x=-848883648;
#10;x=-848783648;
#10;x=-848683648;
#10;x=-848583648;
#10;x=-848483648;
#10;x=-848383648;
#10;x=-848283648;
#10;x=-848183648;
#10;x=-848083648;
#10;x=-847983648;
#10;x=-847883648;
#10;x=-847783648;
#10;x=-847683648;
#10;x=-847583648;
#10;x=-847483648;
#10;x=-847383648;
#10;x=-847283648;
#10;x=-847183648;
#10;x=-847083648;
#10;x=-846983648;
#10;x=-846883648;
#10;x=-846783648;
#10;x=-846683648;
#10;x=-846583648;
#10;x=-846483648;
#10;x=-846383648;
#10;x=-846283648;
#10;x=-846183648;
#10;x=-846083648;
#10;x=-845983648;
#10;x=-845883648;
#10;x=-845783648;
#10;x=-845683648;
#10;x=-845583648;
#10;x=-845483648;
#10;x=-845383648;
#10;x=-845283648;
#10;x=-845183648;
#10;x=-845083648;
#10;x=-844983648;
#10;x=-844883648;
#10;x=-844783648;
#10;x=-844683648;
#10;x=-844583648;
#10;x=-844483648;
#10;x=-844383648;
#10;x=-844283648;
#10;x=-844183648;
#10;x=-844083648;
#10;x=-843983648;
#10;x=-843883648;
#10;x=-843783648;
#10;x=-843683648;
#10;x=-843583648;
#10;x=-843483648;
#10;x=-843383648;
#10;x=-843283648;
#10;x=-843183648;
#10;x=-843083648;
#10;x=-842983648;
#10;x=-842883648;
#10;x=-842783648;
#10;x=-842683648;
#10;x=-842583648;
#10;x=-842483648;
#10;x=-842383648;
#10;x=-842283648;
#10;x=-842183648;
#10;x=-842083648;
#10;x=-841983648;
#10;x=-841883648;
#10;x=-841783648;
#10;x=-841683648;
#10;x=-841583648;
#10;x=-841483648;
#10;x=-841383648;
#10;x=-841283648;
#10;x=-841183648;
#10;x=-841083648;
#10;x=-840983648;
#10;x=-840883648;
#10;x=-840783648;
#10;x=-840683648;
#10;x=-840583648;
#10;x=-840483648;
#10;x=-840383648;
#10;x=-840283648;
#10;x=-840183648;
#10;x=-840083648;
#10;x=-839983648;
#10;x=-839883648;
#10;x=-839783648;
#10;x=-839683648;
#10;x=-839583648;
#10;x=-839483648;
#10;x=-839383648;
#10;x=-839283648;
#10;x=-839183648;
#10;x=-839083648;
#10;x=-838983648;
#10;x=-838883648;
#10;x=-838783648;
#10;x=-838683648;
#10;x=-838583648;
#10;x=-838483648;
#10;x=-838383648;
#10;x=-838283648;
#10;x=-838183648;
#10;x=-838083648;
#10;x=-837983648;
#10;x=-837883648;
#10;x=-837783648;
#10;x=-837683648;
#10;x=-837583648;
#10;x=-837483648;
#10;x=-837383648;
#10;x=-837283648;
#10;x=-837183648;
#10;x=-837083648;
#10;x=-836983648;
#10;x=-836883648;
#10;x=-836783648;
#10;x=-836683648;
#10;x=-836583648;
#10;x=-836483648;
#10;x=-836383648;
#10;x=-836283648;
#10;x=-836183648;
#10;x=-836083648;
#10;x=-835983648;
#10;x=-835883648;
#10;x=-835783648;
#10;x=-835683648;
#10;x=-835583648;
#10;x=-835483648;
#10;x=-835383648;
#10;x=-835283648;
#10;x=-835183648;
#10;x=-835083648;
#10;x=-834983648;
#10;x=-834883648;
#10;x=-834783648;
#10;x=-834683648;
#10;x=-834583648;
#10;x=-834483648;
#10;x=-834383648;
#10;x=-834283648;
#10;x=-834183648;
#10;x=-834083648;
#10;x=-833983648;
#10;x=-833883648;
#10;x=-833783648;
#10;x=-833683648;
#10;x=-833583648;
#10;x=-833483648;
#10;x=-833383648;
#10;x=-833283648;
#10;x=-833183648;
#10;x=-833083648;
#10;x=-832983648;
#10;x=-832883648;
#10;x=-832783648;
#10;x=-832683648;
#10;x=-832583648;
#10;x=-832483648;
#10;x=-832383648;
#10;x=-832283648;
#10;x=-832183648;
#10;x=-832083648;
#10;x=-831983648;
#10;x=-831883648;
#10;x=-831783648;
#10;x=-831683648;
#10;x=-831583648;
#10;x=-831483648;
#10;x=-831383648;
#10;x=-831283648;
#10;x=-831183648;
#10;x=-831083648;
#10;x=-830983648;
#10;x=-830883648;
#10;x=-830783648;
#10;x=-830683648;
#10;x=-830583648;
#10;x=-830483648;
#10;x=-830383648;
#10;x=-830283648;
#10;x=-830183648;
#10;x=-830083648;
#10;x=-829983648;
#10;x=-829883648;
#10;x=-829783648;
#10;x=-829683648;
#10;x=-829583648;
#10;x=-829483648;
#10;x=-829383648;
#10;x=-829283648;
#10;x=-829183648;
#10;x=-829083648;
#10;x=-828983648;
#10;x=-828883648;
#10;x=-828783648;
#10;x=-828683648;
#10;x=-828583648;
#10;x=-828483648;
#10;x=-828383648;
#10;x=-828283648;
#10;x=-828183648;
#10;x=-828083648;
#10;x=-827983648;
#10;x=-827883648;
#10;x=-827783648;
#10;x=-827683648;
#10;x=-827583648;
#10;x=-827483648;
#10;x=-827383648;
#10;x=-827283648;
#10;x=-827183648;
#10;x=-827083648;
#10;x=-826983648;
#10;x=-826883648;
#10;x=-826783648;
#10;x=-826683648;
#10;x=-826583648;
#10;x=-826483648;
#10;x=-826383648;
#10;x=-826283648;
#10;x=-826183648;
#10;x=-826083648;
#10;x=-825983648;
#10;x=-825883648;
#10;x=-825783648;
#10;x=-825683648;
#10;x=-825583648;
#10;x=-825483648;
#10;x=-825383648;
#10;x=-825283648;
#10;x=-825183648;
#10;x=-825083648;
#10;x=-824983648;
#10;x=-824883648;
#10;x=-824783648;
#10;x=-824683648;
#10;x=-824583648;
#10;x=-824483648;
#10;x=-824383648;
#10;x=-824283648;
#10;x=-824183648;
#10;x=-824083648;
#10;x=-823983648;
#10;x=-823883648;
#10;x=-823783648;
#10;x=-823683648;
#10;x=-823583648;
#10;x=-823483648;
#10;x=-823383648;
#10;x=-823283648;
#10;x=-823183648;
#10;x=-823083648;
#10;x=-822983648;
#10;x=-822883648;
#10;x=-822783648;
#10;x=-822683648;
#10;x=-822583648;
#10;x=-822483648;
#10;x=-822383648;
#10;x=-822283648;
#10;x=-822183648;
#10;x=-822083648;
#10;x=-821983648;
#10;x=-821883648;
#10;x=-821783648;
#10;x=-821683648;
#10;x=-821583648;
#10;x=-821483648;
#10;x=-821383648;
#10;x=-821283648;
#10;x=-821183648;
#10;x=-821083648;
#10;x=-820983648;
#10;x=-820883648;
#10;x=-820783648;
#10;x=-820683648;
#10;x=-820583648;
#10;x=-820483648;
#10;x=-820383648;
#10;x=-820283648;
#10;x=-820183648;
#10;x=-820083648;
#10;x=-819983648;
#10;x=-819883648;
#10;x=-819783648;
#10;x=-819683648;
#10;x=-819583648;
#10;x=-819483648;
#10;x=-819383648;
#10;x=-819283648;
#10;x=-819183648;
#10;x=-819083648;
#10;x=-818983648;
#10;x=-818883648;
#10;x=-818783648;
#10;x=-818683648;
#10;x=-818583648;
#10;x=-818483648;
#10;x=-818383648;
#10;x=-818283648;
#10;x=-818183648;
#10;x=-818083648;
#10;x=-817983648;
#10;x=-817883648;
#10;x=-817783648;
#10;x=-817683648;
#10;x=-817583648;
#10;x=-817483648;
#10;x=-817383648;
#10;x=-817283648;
#10;x=-817183648;
#10;x=-817083648;
#10;x=-816983648;
#10;x=-816883648;
#10;x=-816783648;
#10;x=-816683648;
#10;x=-816583648;
#10;x=-816483648;
#10;x=-816383648;
#10;x=-816283648;
#10;x=-816183648;
#10;x=-816083648;
#10;x=-815983648;
#10;x=-815883648;
#10;x=-815783648;
#10;x=-815683648;
#10;x=-815583648;
#10;x=-815483648;
#10;x=-815383648;
#10;x=-815283648;
#10;x=-815183648;
#10;x=-815083648;
#10;x=-814983648;
#10;x=-814883648;
#10;x=-814783648;
#10;x=-814683648;
#10;x=-814583648;
#10;x=-814483648;
#10;x=-814383648;
#10;x=-814283648;
#10;x=-814183648;
#10;x=-814083648;
#10;x=-813983648;
#10;x=-813883648;
#10;x=-813783648;
#10;x=-813683648;
#10;x=-813583648;
#10;x=-813483648;
#10;x=-813383648;
#10;x=-813283648;
#10;x=-813183648;
#10;x=-813083648;
#10;x=-812983648;
#10;x=-812883648;
#10;x=-812783648;
#10;x=-812683648;
#10;x=-812583648;
#10;x=-812483648;
#10;x=-812383648;
#10;x=-812283648;
#10;x=-812183648;
#10;x=-812083648;
#10;x=-811983648;
#10;x=-811883648;
#10;x=-811783648;
#10;x=-811683648;
#10;x=-811583648;
#10;x=-811483648;
#10;x=-811383648;
#10;x=-811283648;
#10;x=-811183648;
#10;x=-811083648;
#10;x=-810983648;
#10;x=-810883648;
#10;x=-810783648;
#10;x=-810683648;
#10;x=-810583648;
#10;x=-810483648;
#10;x=-810383648;
#10;x=-810283648;
#10;x=-810183648;
#10;x=-810083648;
#10;x=-809983648;
#10;x=-809883648;
#10;x=-809783648;
#10;x=-809683648;
#10;x=-809583648;
#10;x=-809483648;
#10;x=-809383648;
#10;x=-809283648;
#10;x=-809183648;
#10;x=-809083648;
#10;x=-808983648;
#10;x=-808883648;
#10;x=-808783648;
#10;x=-808683648;
#10;x=-808583648;
#10;x=-808483648;
#10;x=-808383648;
#10;x=-808283648;
#10;x=-808183648;
#10;x=-808083648;
#10;x=-807983648;
#10;x=-807883648;
#10;x=-807783648;
#10;x=-807683648;
#10;x=-807583648;
#10;x=-807483648;
#10;x=-807383648;
#10;x=-807283648;
#10;x=-807183648;
#10;x=-807083648;
#10;x=-806983648;
#10;x=-806883648;
#10;x=-806783648;
#10;x=-806683648;
#10;x=-806583648;
#10;x=-806483648;
#10;x=-806383648;
#10;x=-806283648;
#10;x=-806183648;
#10;x=-806083648;
#10;x=-805983648;
#10;x=-805883648;
#10;x=-805783648;
#10;x=-805683648;
#10;x=-805583648;
#10;x=-805483648;
#10;x=-805383648;
#10;x=-805283648;
#10;x=-805183648;
#10;x=-805083648;
#10;x=-804983648;
#10;x=-804883648;
#10;x=-804783648;
#10;x=-804683648;
#10;x=-804583648;
#10;x=-804483648;
#10;x=-804383648;
#10;x=-804283648;
#10;x=-804183648;
#10;x=-804083648;
#10;x=-803983648;
#10;x=-803883648;
#10;x=-803783648;
#10;x=-803683648;
#10;x=-803583648;
#10;x=-803483648;
#10;x=-803383648;
#10;x=-803283648;
#10;x=-803183648;
#10;x=-803083648;
#10;x=-802983648;
#10;x=-802883648;
#10;x=-802783648;
#10;x=-802683648;
#10;x=-802583648;
#10;x=-802483648;
#10;x=-802383648;
#10;x=-802283648;
#10;x=-802183648;
#10;x=-802083648;
#10;x=-801983648;
#10;x=-801883648;
#10;x=-801783648;
#10;x=-801683648;
#10;x=-801583648;
#10;x=-801483648;
#10;x=-801383648;
#10;x=-801283648;
#10;x=-801183648;
#10;x=-801083648;
#10;x=-800983648;
#10;x=-800883648;
#10;x=-800783648;
#10;x=-800683648;
#10;x=-800583648;
#10;x=-800483648;
#10;x=-800383648;
#10;x=-800283648;
#10;x=-800183648;
#10;x=-800083648;
#10;x=-799983648;
#10;x=-799883648;
#10;x=-799783648;
#10;x=-799683648;
#10;x=-799583648;
#10;x=-799483648;
#10;x=-799383648;
#10;x=-799283648;
#10;x=-799183648;
#10;x=-799083648;
#10;x=-798983648;
#10;x=-798883648;
#10;x=-798783648;
#10;x=-798683648;
#10;x=-798583648;
#10;x=-798483648;
#10;x=-798383648;
#10;x=-798283648;
#10;x=-798183648;
#10;x=-798083648;
#10;x=-797983648;
#10;x=-797883648;
#10;x=-797783648;
#10;x=-797683648;
#10;x=-797583648;
#10;x=-797483648;
#10;x=-797383648;
#10;x=-797283648;
#10;x=-797183648;
#10;x=-797083648;
#10;x=-796983648;
#10;x=-796883648;
#10;x=-796783648;
#10;x=-796683648;
#10;x=-796583648;
#10;x=-796483648;
#10;x=-796383648;
#10;x=-796283648;
#10;x=-796183648;
#10;x=-796083648;
#10;x=-795983648;
#10;x=-795883648;
#10;x=-795783648;
#10;x=-795683648;
#10;x=-795583648;
#10;x=-795483648;
#10;x=-795383648;
#10;x=-795283648;
#10;x=-795183648;
#10;x=-795083648;
#10;x=-794983648;
#10;x=-794883648;
#10;x=-794783648;
#10;x=-794683648;
#10;x=-794583648;
#10;x=-794483648;
#10;x=-794383648;
#10;x=-794283648;
#10;x=-794183648;
#10;x=-794083648;
#10;x=-793983648;
#10;x=-793883648;
#10;x=-793783648;
#10;x=-793683648;
#10;x=-793583648;
#10;x=-793483648;
#10;x=-793383648;
#10;x=-793283648;
#10;x=-793183648;
#10;x=-793083648;
#10;x=-792983648;
#10;x=-792883648;
#10;x=-792783648;
#10;x=-792683648;
#10;x=-792583648;
#10;x=-792483648;
#10;x=-792383648;
#10;x=-792283648;
#10;x=-792183648;
#10;x=-792083648;
#10;x=-791983648;
#10;x=-791883648;
#10;x=-791783648;
#10;x=-791683648;
#10;x=-791583648;
#10;x=-791483648;
#10;x=-791383648;
#10;x=-791283648;
#10;x=-791183648;
#10;x=-791083648;
#10;x=-790983648;
#10;x=-790883648;
#10;x=-790783648;
#10;x=-790683648;
#10;x=-790583648;
#10;x=-790483648;
#10;x=-790383648;
#10;x=-790283648;
#10;x=-790183648;
#10;x=-790083648;
#10;x=-789983648;
#10;x=-789883648;
#10;x=-789783648;
#10;x=-789683648;
#10;x=-789583648;
#10;x=-789483648;
#10;x=-789383648;
#10;x=-789283648;
#10;x=-789183648;
#10;x=-789083648;
#10;x=-788983648;
#10;x=-788883648;
#10;x=-788783648;
#10;x=-788683648;
#10;x=-788583648;
#10;x=-788483648;
#10;x=-788383648;
#10;x=-788283648;
#10;x=-788183648;
#10;x=-788083648;
#10;x=-787983648;
#10;x=-787883648;
#10;x=-787783648;
#10;x=-787683648;
#10;x=-787583648;
#10;x=-787483648;
#10;x=-787383648;
#10;x=-787283648;
#10;x=-787183648;
#10;x=-787083648;
#10;x=-786983648;
#10;x=-786883648;
#10;x=-786783648;
#10;x=-786683648;
#10;x=-786583648;
#10;x=-786483648;
#10;x=-786383648;
#10;x=-786283648;
#10;x=-786183648;
#10;x=-786083648;
#10;x=-785983648;
#10;x=-785883648;
#10;x=-785783648;
#10;x=-785683648;
#10;x=-785583648;
#10;x=-785483648;
#10;x=-785383648;
#10;x=-785283648;
#10;x=-785183648;
#10;x=-785083648;
#10;x=-784983648;
#10;x=-784883648;
#10;x=-784783648;
#10;x=-784683648;
#10;x=-784583648;
#10;x=-784483648;
#10;x=-784383648;
#10;x=-784283648;
#10;x=-784183648;
#10;x=-784083648;
#10;x=-783983648;
#10;x=-783883648;
#10;x=-783783648;
#10;x=-783683648;
#10;x=-783583648;
#10;x=-783483648;
#10;x=-783383648;
#10;x=-783283648;
#10;x=-783183648;
#10;x=-783083648;
#10;x=-782983648;
#10;x=-782883648;
#10;x=-782783648;
#10;x=-782683648;
#10;x=-782583648;
#10;x=-782483648;
#10;x=-782383648;
#10;x=-782283648;
#10;x=-782183648;
#10;x=-782083648;
#10;x=-781983648;
#10;x=-781883648;
#10;x=-781783648;
#10;x=-781683648;
#10;x=-781583648;
#10;x=-781483648;
#10;x=-781383648;
#10;x=-781283648;
#10;x=-781183648;
#10;x=-781083648;
#10;x=-780983648;
#10;x=-780883648;
#10;x=-780783648;
#10;x=-780683648;
#10;x=-780583648;
#10;x=-780483648;
#10;x=-780383648;
#10;x=-780283648;
#10;x=-780183648;
#10;x=-780083648;
#10;x=-779983648;
#10;x=-779883648;
#10;x=-779783648;
#10;x=-779683648;
#10;x=-779583648;
#10;x=-779483648;
#10;x=-779383648;
#10;x=-779283648;
#10;x=-779183648;
#10;x=-779083648;
#10;x=-778983648;
#10;x=-778883648;
#10;x=-778783648;
#10;x=-778683648;
#10;x=-778583648;
#10;x=-778483648;
#10;x=-778383648;
#10;x=-778283648;
#10;x=-778183648;
#10;x=-778083648;
#10;x=-777983648;
#10;x=-777883648;
#10;x=-777783648;
#10;x=-777683648;
#10;x=-777583648;
#10;x=-777483648;
#10;x=-777383648;
#10;x=-777283648;
#10;x=-777183648;
#10;x=-777083648;
#10;x=-776983648;
#10;x=-776883648;
#10;x=-776783648;
#10;x=-776683648;
#10;x=-776583648;
#10;x=-776483648;
#10;x=-776383648;
#10;x=-776283648;
#10;x=-776183648;
#10;x=-776083648;
#10;x=-775983648;
#10;x=-775883648;
#10;x=-775783648;
#10;x=-775683648;
#10;x=-775583648;
#10;x=-775483648;
#10;x=-775383648;
#10;x=-775283648;
#10;x=-775183648;
#10;x=-775083648;
#10;x=-774983648;
#10;x=-774883648;
#10;x=-774783648;
#10;x=-774683648;
#10;x=-774583648;
#10;x=-774483648;
#10;x=-774383648;
#10;x=-774283648;
#10;x=-774183648;
#10;x=-774083648;
#10;x=-773983648;
#10;x=-773883648;
#10;x=-773783648;
#10;x=-773683648;
#10;x=-773583648;
#10;x=-773483648;
#10;x=-773383648;
#10;x=-773283648;
#10;x=-773183648;
#10;x=-773083648;
#10;x=-772983648;
#10;x=-772883648;
#10;x=-772783648;
#10;x=-772683648;
#10;x=-772583648;
#10;x=-772483648;
#10;x=-772383648;
#10;x=-772283648;
#10;x=-772183648;
#10;x=-772083648;
#10;x=-771983648;
#10;x=-771883648;
#10;x=-771783648;
#10;x=-771683648;
#10;x=-771583648;
#10;x=-771483648;
#10;x=-771383648;
#10;x=-771283648;
#10;x=-771183648;
#10;x=-771083648;
#10;x=-770983648;
#10;x=-770883648;
#10;x=-770783648;
#10;x=-770683648;
#10;x=-770583648;
#10;x=-770483648;
#10;x=-770383648;
#10;x=-770283648;
#10;x=-770183648;
#10;x=-770083648;
#10;x=-769983648;
#10;x=-769883648;
#10;x=-769783648;
#10;x=-769683648;
#10;x=-769583648;
#10;x=-769483648;
#10;x=-769383648;
#10;x=-769283648;
#10;x=-769183648;
#10;x=-769083648;
#10;x=-768983648;
#10;x=-768883648;
#10;x=-768783648;
#10;x=-768683648;
#10;x=-768583648;
#10;x=-768483648;
#10;x=-768383648;
#10;x=-768283648;
#10;x=-768183648;
#10;x=-768083648;
#10;x=-767983648;
#10;x=-767883648;
#10;x=-767783648;
#10;x=-767683648;
#10;x=-767583648;
#10;x=-767483648;
#10;x=-767383648;
#10;x=-767283648;
#10;x=-767183648;
#10;x=-767083648;
#10;x=-766983648;
#10;x=-766883648;
#10;x=-766783648;
#10;x=-766683648;
#10;x=-766583648;
#10;x=-766483648;
#10;x=-766383648;
#10;x=-766283648;
#10;x=-766183648;
#10;x=-766083648;
#10;x=-765983648;
#10;x=-765883648;
#10;x=-765783648;
#10;x=-765683648;
#10;x=-765583648;
#10;x=-765483648;
#10;x=-765383648;
#10;x=-765283648;
#10;x=-765183648;
#10;x=-765083648;
#10;x=-764983648;
#10;x=-764883648;
#10;x=-764783648;
#10;x=-764683648;
#10;x=-764583648;
#10;x=-764483648;
#10;x=-764383648;
#10;x=-764283648;
#10;x=-764183648;
#10;x=-764083648;
#10;x=-763983648;
#10;x=-763883648;
#10;x=-763783648;
#10;x=-763683648;
#10;x=-763583648;
#10;x=-763483648;
#10;x=-763383648;
#10;x=-763283648;
#10;x=-763183648;
#10;x=-763083648;
#10;x=-762983648;
#10;x=-762883648;
#10;x=-762783648;
#10;x=-762683648;
#10;x=-762583648;
#10;x=-762483648;
#10;x=-762383648;
#10;x=-762283648;
#10;x=-762183648;
#10;x=-762083648;
#10;x=-761983648;
#10;x=-761883648;
#10;x=-761783648;
#10;x=-761683648;
#10;x=-761583648;
#10;x=-761483648;
#10;x=-761383648;
#10;x=-761283648;
#10;x=-761183648;
#10;x=-761083648;
#10;x=-760983648;
#10;x=-760883648;
#10;x=-760783648;
#10;x=-760683648;
#10;x=-760583648;
#10;x=-760483648;
#10;x=-760383648;
#10;x=-760283648;
#10;x=-760183648;
#10;x=-760083648;
#10;x=-759983648;
#10;x=-759883648;
#10;x=-759783648;
#10;x=-759683648;
#10;x=-759583648;
#10;x=-759483648;
#10;x=-759383648;
#10;x=-759283648;
#10;x=-759183648;
#10;x=-759083648;
#10;x=-758983648;
#10;x=-758883648;
#10;x=-758783648;
#10;x=-758683648;
#10;x=-758583648;
#10;x=-758483648;
#10;x=-758383648;
#10;x=-758283648;
#10;x=-758183648;
#10;x=-758083648;
#10;x=-757983648;
#10;x=-757883648;
#10;x=-757783648;
#10;x=-757683648;
#10;x=-757583648;
#10;x=-757483648;
#10;x=-757383648;
#10;x=-757283648;
#10;x=-757183648;
#10;x=-757083648;
#10;x=-756983648;
#10;x=-756883648;
#10;x=-756783648;
#10;x=-756683648;
#10;x=-756583648;
#10;x=-756483648;
#10;x=-756383648;
#10;x=-756283648;
#10;x=-756183648;
#10;x=-756083648;
#10;x=-755983648;
#10;x=-755883648;
#10;x=-755783648;
#10;x=-755683648;
#10;x=-755583648;
#10;x=-755483648;
#10;x=-755383648;
#10;x=-755283648;
#10;x=-755183648;
#10;x=-755083648;
#10;x=-754983648;
#10;x=-754883648;
#10;x=-754783648;
#10;x=-754683648;
#10;x=-754583648;
#10;x=-754483648;
#10;x=-754383648;
#10;x=-754283648;
#10;x=-754183648;
#10;x=-754083648;
#10;x=-753983648;
#10;x=-753883648;
#10;x=-753783648;
#10;x=-753683648;
#10;x=-753583648;
#10;x=-753483648;
#10;x=-753383648;
#10;x=-753283648;
#10;x=-753183648;
#10;x=-753083648;
#10;x=-752983648;
#10;x=-752883648;
#10;x=-752783648;
#10;x=-752683648;
#10;x=-752583648;
#10;x=-752483648;
#10;x=-752383648;
#10;x=-752283648;
#10;x=-752183648;
#10;x=-752083648;
#10;x=-751983648;
#10;x=-751883648;
#10;x=-751783648;
#10;x=-751683648;
#10;x=-751583648;
#10;x=-751483648;
#10;x=-751383648;
#10;x=-751283648;
#10;x=-751183648;
#10;x=-751083648;
#10;x=-750983648;
#10;x=-750883648;
#10;x=-750783648;
#10;x=-750683648;
#10;x=-750583648;
#10;x=-750483648;
#10;x=-750383648;
#10;x=-750283648;
#10;x=-750183648;
#10;x=-750083648;
#10;x=-749983648;
#10;x=-749883648;
#10;x=-749783648;
#10;x=-749683648;
#10;x=-749583648;
#10;x=-749483648;
#10;x=-749383648;
#10;x=-749283648;
#10;x=-749183648;
#10;x=-749083648;
#10;x=-748983648;
#10;x=-748883648;
#10;x=-748783648;
#10;x=-748683648;
#10;x=-748583648;
#10;x=-748483648;
#10;x=-748383648;
#10;x=-748283648;
#10;x=-748183648;
#10;x=-748083648;
#10;x=-747983648;
#10;x=-747883648;
#10;x=-747783648;
#10;x=-747683648;
#10;x=-747583648;
#10;x=-747483648;
#10;x=-747383648;
#10;x=-747283648;
#10;x=-747183648;
#10;x=-747083648;
#10;x=-746983648;
#10;x=-746883648;
#10;x=-746783648;
#10;x=-746683648;
#10;x=-746583648;
#10;x=-746483648;
#10;x=-746383648;
#10;x=-746283648;
#10;x=-746183648;
#10;x=-746083648;
#10;x=-745983648;
#10;x=-745883648;
#10;x=-745783648;
#10;x=-745683648;
#10;x=-745583648;
#10;x=-745483648;
#10;x=-745383648;
#10;x=-745283648;
#10;x=-745183648;
#10;x=-745083648;
#10;x=-744983648;
#10;x=-744883648;
#10;x=-744783648;
#10;x=-744683648;
#10;x=-744583648;
#10;x=-744483648;
#10;x=-744383648;
#10;x=-744283648;
#10;x=-744183648;
#10;x=-744083648;
#10;x=-743983648;
#10;x=-743883648;
#10;x=-743783648;
#10;x=-743683648;
#10;x=-743583648;
#10;x=-743483648;
#10;x=-743383648;
#10;x=-743283648;
#10;x=-743183648;
#10;x=-743083648;
#10;x=-742983648;
#10;x=-742883648;
#10;x=-742783648;
#10;x=-742683648;
#10;x=-742583648;
#10;x=-742483648;
#10;x=-742383648;
#10;x=-742283648;
#10;x=-742183648;
#10;x=-742083648;
#10;x=-741983648;
#10;x=-741883648;
#10;x=-741783648;
#10;x=-741683648;
#10;x=-741583648;
#10;x=-741483648;
#10;x=-741383648;
#10;x=-741283648;
#10;x=-741183648;
#10;x=-741083648;
#10;x=-740983648;
#10;x=-740883648;
#10;x=-740783648;
#10;x=-740683648;
#10;x=-740583648;
#10;x=-740483648;
#10;x=-740383648;
#10;x=-740283648;
#10;x=-740183648;
#10;x=-740083648;
#10;x=-739983648;
#10;x=-739883648;
#10;x=-739783648;
#10;x=-739683648;
#10;x=-739583648;
#10;x=-739483648;
#10;x=-739383648;
#10;x=-739283648;
#10;x=-739183648;
#10;x=-739083648;
#10;x=-738983648;
#10;x=-738883648;
#10;x=-738783648;
#10;x=-738683648;
#10;x=-738583648;
#10;x=-738483648;
#10;x=-738383648;
#10;x=-738283648;
#10;x=-738183648;
#10;x=-738083648;
#10;x=-737983648;
#10;x=-737883648;
#10;x=-737783648;
#10;x=-737683648;
#10;x=-737583648;
#10;x=-737483648;
#10;x=-737383648;
#10;x=-737283648;
#10;x=-737183648;
#10;x=-737083648;
#10;x=-736983648;
#10;x=-736883648;
#10;x=-736783648;
#10;x=-736683648;
#10;x=-736583648;
#10;x=-736483648;
#10;x=-736383648;
#10;x=-736283648;
#10;x=-736183648;
#10;x=-736083648;
#10;x=-735983648;
#10;x=-735883648;
#10;x=-735783648;
#10;x=-735683648;
#10;x=-735583648;
#10;x=-735483648;
#10;x=-735383648;
#10;x=-735283648;
#10;x=-735183648;
#10;x=-735083648;
#10;x=-734983648;
#10;x=-734883648;
#10;x=-734783648;
#10;x=-734683648;
#10;x=-734583648;
#10;x=-734483648;
#10;x=-734383648;
#10;x=-734283648;
#10;x=-734183648;
#10;x=-734083648;
#10;x=-733983648;
#10;x=-733883648;
#10;x=-733783648;
#10;x=-733683648;
#10;x=-733583648;
#10;x=-733483648;
#10;x=-733383648;
#10;x=-733283648;
#10;x=-733183648;
#10;x=-733083648;
#10;x=-732983648;
#10;x=-732883648;
#10;x=-732783648;
#10;x=-732683648;
#10;x=-732583648;
#10;x=-732483648;
#10;x=-732383648;
#10;x=-732283648;
#10;x=-732183648;
#10;x=-732083648;
#10;x=-731983648;
#10;x=-731883648;
#10;x=-731783648;
#10;x=-731683648;
#10;x=-731583648;
#10;x=-731483648;
#10;x=-731383648;
#10;x=-731283648;
#10;x=-731183648;
#10;x=-731083648;
#10;x=-730983648;
#10;x=-730883648;
#10;x=-730783648;
#10;x=-730683648;
#10;x=-730583648;
#10;x=-730483648;
#10;x=-730383648;
#10;x=-730283648;
#10;x=-730183648;
#10;x=-730083648;
#10;x=-729983648;
#10;x=-729883648;
#10;x=-729783648;
#10;x=-729683648;
#10;x=-729583648;
#10;x=-729483648;
#10;x=-729383648;
#10;x=-729283648;
#10;x=-729183648;
#10;x=-729083648;
#10;x=-728983648;
#10;x=-728883648;
#10;x=-728783648;
#10;x=-728683648;
#10;x=-728583648;
#10;x=-728483648;
#10;x=-728383648;
#10;x=-728283648;
#10;x=-728183648;
#10;x=-728083648;
#10;x=-727983648;
#10;x=-727883648;
#10;x=-727783648;
#10;x=-727683648;
#10;x=-727583648;
#10;x=-727483648;
#10;x=-727383648;
#10;x=-727283648;
#10;x=-727183648;
#10;x=-727083648;
#10;x=-726983648;
#10;x=-726883648;
#10;x=-726783648;
#10;x=-726683648;
#10;x=-726583648;
#10;x=-726483648;
#10;x=-726383648;
#10;x=-726283648;
#10;x=-726183648;
#10;x=-726083648;
#10;x=-725983648;
#10;x=-725883648;
#10;x=-725783648;
#10;x=-725683648;
#10;x=-725583648;
#10;x=-725483648;
#10;x=-725383648;
#10;x=-725283648;
#10;x=-725183648;
#10;x=-725083648;
#10;x=-724983648;
#10;x=-724883648;
#10;x=-724783648;
#10;x=-724683648;
#10;x=-724583648;
#10;x=-724483648;
#10;x=-724383648;
#10;x=-724283648;
#10;x=-724183648;
#10;x=-724083648;
#10;x=-723983648;
#10;x=-723883648;
#10;x=-723783648;
#10;x=-723683648;
#10;x=-723583648;
#10;x=-723483648;
#10;x=-723383648;
#10;x=-723283648;
#10;x=-723183648;
#10;x=-723083648;
#10;x=-722983648;
#10;x=-722883648;
#10;x=-722783648;
#10;x=-722683648;
#10;x=-722583648;
#10;x=-722483648;
#10;x=-722383648;
#10;x=-722283648;
#10;x=-722183648;
#10;x=-722083648;
#10;x=-721983648;
#10;x=-721883648;
#10;x=-721783648;
#10;x=-721683648;
#10;x=-721583648;
#10;x=-721483648;
#10;x=-721383648;
#10;x=-721283648;
#10;x=-721183648;
#10;x=-721083648;
#10;x=-720983648;
#10;x=-720883648;
#10;x=-720783648;
#10;x=-720683648;
#10;x=-720583648;
#10;x=-720483648;
#10;x=-720383648;
#10;x=-720283648;
#10;x=-720183648;
#10;x=-720083648;
#10;x=-719983648;
#10;x=-719883648;
#10;x=-719783648;
#10;x=-719683648;
#10;x=-719583648;
#10;x=-719483648;
#10;x=-719383648;
#10;x=-719283648;
#10;x=-719183648;
#10;x=-719083648;
#10;x=-718983648;
#10;x=-718883648;
#10;x=-718783648;
#10;x=-718683648;
#10;x=-718583648;
#10;x=-718483648;
#10;x=-718383648;
#10;x=-718283648;
#10;x=-718183648;
#10;x=-718083648;
#10;x=-717983648;
#10;x=-717883648;
#10;x=-717783648;
#10;x=-717683648;
#10;x=-717583648;
#10;x=-717483648;
#10;x=-717383648;
#10;x=-717283648;
#10;x=-717183648;
#10;x=-717083648;
#10;x=-716983648;
#10;x=-716883648;
#10;x=-716783648;
#10;x=-716683648;
#10;x=-716583648;
#10;x=-716483648;
#10;x=-716383648;
#10;x=-716283648;
#10;x=-716183648;
#10;x=-716083648;
#10;x=-715983648;
#10;x=-715883648;
#10;x=-715783648;
#10;x=-715683648;
#10;x=-715583648;
#10;x=-715483648;
#10;x=-715383648;
#10;x=-715283648;
#10;x=-715183648;
#10;x=-715083648;
#10;x=-714983648;
#10;x=-714883648;
#10;x=-714783648;
#10;x=-714683648;
#10;x=-714583648;
#10;x=-714483648;
#10;x=-714383648;
#10;x=-714283648;
#10;x=-714183648;
#10;x=-714083648;
#10;x=-713983648;
#10;x=-713883648;
#10;x=-713783648;
#10;x=-713683648;
#10;x=-713583648;
#10;x=-713483648;
#10;x=-713383648;
#10;x=-713283648;
#10;x=-713183648;
#10;x=-713083648;
#10;x=-712983648;
#10;x=-712883648;
#10;x=-712783648;
#10;x=-712683648;
#10;x=-712583648;
#10;x=-712483648;
#10;x=-712383648;
#10;x=-712283648;
#10;x=-712183648;
#10;x=-712083648;
#10;x=-711983648;
#10;x=-711883648;
#10;x=-711783648;
#10;x=-711683648;
#10;x=-711583648;
#10;x=-711483648;
#10;x=-711383648;
#10;x=-711283648;
#10;x=-711183648;
#10;x=-711083648;
#10;x=-710983648;
#10;x=-710883648;
#10;x=-710783648;
#10;x=-710683648;
#10;x=-710583648;
#10;x=-710483648;
#10;x=-710383648;
#10;x=-710283648;
#10;x=-710183648;
#10;x=-710083648;
#10;x=-709983648;
#10;x=-709883648;
#10;x=-709783648;
#10;x=-709683648;
#10;x=-709583648;
#10;x=-709483648;
#10;x=-709383648;
#10;x=-709283648;
#10;x=-709183648;
#10;x=-709083648;
#10;x=-708983648;
#10;x=-708883648;
#10;x=-708783648;
#10;x=-708683648;
#10;x=-708583648;
#10;x=-708483648;
#10;x=-708383648;
#10;x=-708283648;
#10;x=-708183648;
#10;x=-708083648;
#10;x=-707983648;
#10;x=-707883648;
#10;x=-707783648;
#10;x=-707683648;
#10;x=-707583648;
#10;x=-707483648;
#10;x=-707383648;
#10;x=-707283648;
#10;x=-707183648;
#10;x=-707083648;
#10;x=-706983648;
#10;x=-706883648;
#10;x=-706783648;
#10;x=-706683648;
#10;x=-706583648;
#10;x=-706483648;
#10;x=-706383648;
#10;x=-706283648;
#10;x=-706183648;
#10;x=-706083648;
#10;x=-705983648;
#10;x=-705883648;
#10;x=-705783648;
#10;x=-705683648;
#10;x=-705583648;
#10;x=-705483648;
#10;x=-705383648;
#10;x=-705283648;
#10;x=-705183648;
#10;x=-705083648;
#10;x=-704983648;
#10;x=-704883648;
#10;x=-704783648;
#10;x=-704683648;
#10;x=-704583648;
#10;x=-704483648;
#10;x=-704383648;
#10;x=-704283648;
#10;x=-704183648;
#10;x=-704083648;
#10;x=-703983648;
#10;x=-703883648;
#10;x=-703783648;
#10;x=-703683648;
#10;x=-703583648;
#10;x=-703483648;
#10;x=-703383648;
#10;x=-703283648;
#10;x=-703183648;
#10;x=-703083648;
#10;x=-702983648;
#10;x=-702883648;
#10;x=-702783648;
#10;x=-702683648;
#10;x=-702583648;
#10;x=-702483648;
#10;x=-702383648;
#10;x=-702283648;
#10;x=-702183648;
#10;x=-702083648;
#10;x=-701983648;
#10;x=-701883648;
#10;x=-701783648;
#10;x=-701683648;
#10;x=-701583648;
#10;x=-701483648;
#10;x=-701383648;
#10;x=-701283648;
#10;x=-701183648;
#10;x=-701083648;
#10;x=-700983648;
#10;x=-700883648;
#10;x=-700783648;
#10;x=-700683648;
#10;x=-700583648;
#10;x=-700483648;
#10;x=-700383648;
#10;x=-700283648;
#10;x=-700183648;
#10;x=-700083648;
#10;x=-699983648;
#10;x=-699883648;
#10;x=-699783648;
#10;x=-699683648;
#10;x=-699583648;
#10;x=-699483648;
#10;x=-699383648;
#10;x=-699283648;
#10;x=-699183648;
#10;x=-699083648;
#10;x=-698983648;
#10;x=-698883648;
#10;x=-698783648;
#10;x=-698683648;
#10;x=-698583648;
#10;x=-698483648;
#10;x=-698383648;
#10;x=-698283648;
#10;x=-698183648;
#10;x=-698083648;
#10;x=-697983648;
#10;x=-697883648;
#10;x=-697783648;
#10;x=-697683648;
#10;x=-697583648;
#10;x=-697483648;
#10;x=-697383648;
#10;x=-697283648;
#10;x=-697183648;
#10;x=-697083648;
#10;x=-696983648;
#10;x=-696883648;
#10;x=-696783648;
#10;x=-696683648;
#10;x=-696583648;
#10;x=-696483648;
#10;x=-696383648;
#10;x=-696283648;
#10;x=-696183648;
#10;x=-696083648;
#10;x=-695983648;
#10;x=-695883648;
#10;x=-695783648;
#10;x=-695683648;
#10;x=-695583648;
#10;x=-695483648;
#10;x=-695383648;
#10;x=-695283648;
#10;x=-695183648;
#10;x=-695083648;
#10;x=-694983648;
#10;x=-694883648;
#10;x=-694783648;
#10;x=-694683648;
#10;x=-694583648;
#10;x=-694483648;
#10;x=-694383648;
#10;x=-694283648;
#10;x=-694183648;
#10;x=-694083648;
#10;x=-693983648;
#10;x=-693883648;
#10;x=-693783648;
#10;x=-693683648;
#10;x=-693583648;
#10;x=-693483648;
#10;x=-693383648;
#10;x=-693283648;
#10;x=-693183648;
#10;x=-693083648;
#10;x=-692983648;
#10;x=-692883648;
#10;x=-692783648;
#10;x=-692683648;
#10;x=-692583648;
#10;x=-692483648;
#10;x=-692383648;
#10;x=-692283648;
#10;x=-692183648;
#10;x=-692083648;
#10;x=-691983648;
#10;x=-691883648;
#10;x=-691783648;
#10;x=-691683648;
#10;x=-691583648;
#10;x=-691483648;
#10;x=-691383648;
#10;x=-691283648;
#10;x=-691183648;
#10;x=-691083648;
#10;x=-690983648;
#10;x=-690883648;
#10;x=-690783648;
#10;x=-690683648;
#10;x=-690583648;
#10;x=-690483648;
#10;x=-690383648;
#10;x=-690283648;
#10;x=-690183648;
#10;x=-690083648;
#10;x=-689983648;
#10;x=-689883648;
#10;x=-689783648;
#10;x=-689683648;
#10;x=-689583648;
#10;x=-689483648;
#10;x=-689383648;
#10;x=-689283648;
#10;x=-689183648;
#10;x=-689083648;
#10;x=-688983648;
#10;x=-688883648;
#10;x=-688783648;
#10;x=-688683648;
#10;x=-688583648;
#10;x=-688483648;
#10;x=-688383648;
#10;x=-688283648;
#10;x=-688183648;
#10;x=-688083648;
#10;x=-687983648;
#10;x=-687883648;
#10;x=-687783648;
#10;x=-687683648;
#10;x=-687583648;
#10;x=-687483648;
#10;x=-687383648;
#10;x=-687283648;
#10;x=-687183648;
#10;x=-687083648;
#10;x=-686983648;
#10;x=-686883648;
#10;x=-686783648;
#10;x=-686683648;
#10;x=-686583648;
#10;x=-686483648;
#10;x=-686383648;
#10;x=-686283648;
#10;x=-686183648;
#10;x=-686083648;
#10;x=-685983648;
#10;x=-685883648;
#10;x=-685783648;
#10;x=-685683648;
#10;x=-685583648;
#10;x=-685483648;
#10;x=-685383648;
#10;x=-685283648;
#10;x=-685183648;
#10;x=-685083648;
#10;x=-684983648;
#10;x=-684883648;
#10;x=-684783648;
#10;x=-684683648;
#10;x=-684583648;
#10;x=-684483648;
#10;x=-684383648;
#10;x=-684283648;
#10;x=-684183648;
#10;x=-684083648;
#10;x=-683983648;
#10;x=-683883648;
#10;x=-683783648;
#10;x=-683683648;
#10;x=-683583648;
#10;x=-683483648;
#10;x=-683383648;
#10;x=-683283648;
#10;x=-683183648;
#10;x=-683083648;
#10;x=-682983648;
#10;x=-682883648;
#10;x=-682783648;
#10;x=-682683648;
#10;x=-682583648;
#10;x=-682483648;
#10;x=-682383648;
#10;x=-682283648;
#10;x=-682183648;
#10;x=-682083648;
#10;x=-681983648;
#10;x=-681883648;
#10;x=-681783648;
#10;x=-681683648;
#10;x=-681583648;
#10;x=-681483648;
#10;x=-681383648;
#10;x=-681283648;
#10;x=-681183648;
#10;x=-681083648;
#10;x=-680983648;
#10;x=-680883648;
#10;x=-680783648;
#10;x=-680683648;
#10;x=-680583648;
#10;x=-680483648;
#10;x=-680383648;
#10;x=-680283648;
#10;x=-680183648;
#10;x=-680083648;
#10;x=-679983648;
#10;x=-679883648;
#10;x=-679783648;
#10;x=-679683648;
#10;x=-679583648;
#10;x=-679483648;
#10;x=-679383648;
#10;x=-679283648;
#10;x=-679183648;
#10;x=-679083648;
#10;x=-678983648;
#10;x=-678883648;
#10;x=-678783648;
#10;x=-678683648;
#10;x=-678583648;
#10;x=-678483648;
#10;x=-678383648;
#10;x=-678283648;
#10;x=-678183648;
#10;x=-678083648;
#10;x=-677983648;
#10;x=-677883648;
#10;x=-677783648;
#10;x=-677683648;
#10;x=-677583648;
#10;x=-677483648;
#10;x=-677383648;
#10;x=-677283648;
#10;x=-677183648;
#10;x=-677083648;
#10;x=-676983648;
#10;x=-676883648;
#10;x=-676783648;
#10;x=-676683648;
#10;x=-676583648;
#10;x=-676483648;
#10;x=-676383648;
#10;x=-676283648;
#10;x=-676183648;
#10;x=-676083648;
#10;x=-675983648;
#10;x=-675883648;
#10;x=-675783648;
#10;x=-675683648;
#10;x=-675583648;
#10;x=-675483648;
#10;x=-675383648;
#10;x=-675283648;
#10;x=-675183648;
#10;x=-675083648;
#10;x=-674983648;
#10;x=-674883648;
#10;x=-674783648;
#10;x=-674683648;
#10;x=-674583648;
#10;x=-674483648;
#10;x=-674383648;
#10;x=-674283648;
#10;x=-674183648;
#10;x=-674083648;
#10;x=-673983648;
#10;x=-673883648;
#10;x=-673783648;
#10;x=-673683648;
#10;x=-673583648;
#10;x=-673483648;
#10;x=-673383648;
#10;x=-673283648;
#10;x=-673183648;
#10;x=-673083648;
#10;x=-672983648;
#10;x=-672883648;
#10;x=-672783648;
#10;x=-672683648;
#10;x=-672583648;
#10;x=-672483648;
#10;x=-672383648;
#10;x=-672283648;
#10;x=-672183648;
#10;x=-672083648;
#10;x=-671983648;
#10;x=-671883648;
#10;x=-671783648;
#10;x=-671683648;
#10;x=-671583648;
#10;x=-671483648;
#10;x=-671383648;
#10;x=-671283648;
#10;x=-671183648;
#10;x=-671083648;
#10;x=-670983648;
#10;x=-670883648;
#10;x=-670783648;
#10;x=-670683648;
#10;x=-670583648;
#10;x=-670483648;
#10;x=-670383648;
#10;x=-670283648;
#10;x=-670183648;
#10;x=-670083648;
#10;x=-669983648;
#10;x=-669883648;
#10;x=-669783648;
#10;x=-669683648;
#10;x=-669583648;
#10;x=-669483648;
#10;x=-669383648;
#10;x=-669283648;
#10;x=-669183648;
#10;x=-669083648;
#10;x=-668983648;
#10;x=-668883648;
#10;x=-668783648;
#10;x=-668683648;
#10;x=-668583648;
#10;x=-668483648;
#10;x=-668383648;
#10;x=-668283648;
#10;x=-668183648;
#10;x=-668083648;
#10;x=-667983648;
#10;x=-667883648;
#10;x=-667783648;
#10;x=-667683648;
#10;x=-667583648;
#10;x=-667483648;
#10;x=-667383648;
#10;x=-667283648;
#10;x=-667183648;
#10;x=-667083648;
#10;x=-666983648;
#10;x=-666883648;
#10;x=-666783648;
#10;x=-666683648;
#10;x=-666583648;
#10;x=-666483648;
#10;x=-666383648;
#10;x=-666283648;
#10;x=-666183648;
#10;x=-666083648;
#10;x=-665983648;
#10;x=-665883648;
#10;x=-665783648;
#10;x=-665683648;
#10;x=-665583648;
#10;x=-665483648;
#10;x=-665383648;
#10;x=-665283648;
#10;x=-665183648;
#10;x=-665083648;
#10;x=-664983648;
#10;x=-664883648;
#10;x=-664783648;
#10;x=-664683648;
#10;x=-664583648;
#10;x=-664483648;
#10;x=-664383648;
#10;x=-664283648;
#10;x=-664183648;
#10;x=-664083648;
#10;x=-663983648;
#10;x=-663883648;
#10;x=-663783648;
#10;x=-663683648;
#10;x=-663583648;
#10;x=-663483648;
#10;x=-663383648;
#10;x=-663283648;
#10;x=-663183648;
#10;x=-663083648;
#10;x=-662983648;
#10;x=-662883648;
#10;x=-662783648;
#10;x=-662683648;
#10;x=-662583648;
#10;x=-662483648;
#10;x=-662383648;
#10;x=-662283648;
#10;x=-662183648;
#10;x=-662083648;
#10;x=-661983648;
#10;x=-661883648;
#10;x=-661783648;
#10;x=-661683648;
#10;x=-661583648;
#10;x=-661483648;
#10;x=-661383648;
#10;x=-661283648;
#10;x=-661183648;
#10;x=-661083648;
#10;x=-660983648;
#10;x=-660883648;
#10;x=-660783648;
#10;x=-660683648;
#10;x=-660583648;
#10;x=-660483648;
#10;x=-660383648;
#10;x=-660283648;
#10;x=-660183648;
#10;x=-660083648;
#10;x=-659983648;
#10;x=-659883648;
#10;x=-659783648;
#10;x=-659683648;
#10;x=-659583648;
#10;x=-659483648;
#10;x=-659383648;
#10;x=-659283648;
#10;x=-659183648;
#10;x=-659083648;
#10;x=-658983648;
#10;x=-658883648;
#10;x=-658783648;
#10;x=-658683648;
#10;x=-658583648;
#10;x=-658483648;
#10;x=-658383648;
#10;x=-658283648;
#10;x=-658183648;
#10;x=-658083648;
#10;x=-657983648;
#10;x=-657883648;
#10;x=-657783648;
#10;x=-657683648;
#10;x=-657583648;
#10;x=-657483648;
#10;x=-657383648;
#10;x=-657283648;
#10;x=-657183648;
#10;x=-657083648;
#10;x=-656983648;
#10;x=-656883648;
#10;x=-656783648;
#10;x=-656683648;
#10;x=-656583648;
#10;x=-656483648;
#10;x=-656383648;
#10;x=-656283648;
#10;x=-656183648;
#10;x=-656083648;
#10;x=-655983648;
#10;x=-655883648;
#10;x=-655783648;
#10;x=-655683648;
#10;x=-655583648;
#10;x=-655483648;
#10;x=-655383648;
#10;x=-655283648;
#10;x=-655183648;
#10;x=-655083648;
#10;x=-654983648;
#10;x=-654883648;
#10;x=-654783648;
#10;x=-654683648;
#10;x=-654583648;
#10;x=-654483648;
#10;x=-654383648;
#10;x=-654283648;
#10;x=-654183648;
#10;x=-654083648;
#10;x=-653983648;
#10;x=-653883648;
#10;x=-653783648;
#10;x=-653683648;
#10;x=-653583648;
#10;x=-653483648;
#10;x=-653383648;
#10;x=-653283648;
#10;x=-653183648;
#10;x=-653083648;
#10;x=-652983648;
#10;x=-652883648;
#10;x=-652783648;
#10;x=-652683648;
#10;x=-652583648;
#10;x=-652483648;
#10;x=-652383648;
#10;x=-652283648;
#10;x=-652183648;
#10;x=-652083648;
#10;x=-651983648;
#10;x=-651883648;
#10;x=-651783648;
#10;x=-651683648;
#10;x=-651583648;
#10;x=-651483648;
#10;x=-651383648;
#10;x=-651283648;
#10;x=-651183648;
#10;x=-651083648;
#10;x=-650983648;
#10;x=-650883648;
#10;x=-650783648;
#10;x=-650683648;
#10;x=-650583648;
#10;x=-650483648;
#10;x=-650383648;
#10;x=-650283648;
#10;x=-650183648;
#10;x=-650083648;
#10;x=-649983648;
#10;x=-649883648;
#10;x=-649783648;
#10;x=-649683648;
#10;x=-649583648;
#10;x=-649483648;
#10;x=-649383648;
#10;x=-649283648;
#10;x=-649183648;
#10;x=-649083648;
#10;x=-648983648;
#10;x=-648883648;
#10;x=-648783648;
#10;x=-648683648;
#10;x=-648583648;
#10;x=-648483648;
#10;x=-648383648;
#10;x=-648283648;
#10;x=-648183648;
#10;x=-648083648;
#10;x=-647983648;
#10;x=-647883648;
#10;x=-647783648;
#10;x=-647683648;
#10;x=-647583648;
#10;x=-647483648;
#10;x=-647383648;
#10;x=-647283648;
#10;x=-647183648;
#10;x=-647083648;
#10;x=-646983648;
#10;x=-646883648;
#10;x=-646783648;
#10;x=-646683648;
#10;x=-646583648;
#10;x=-646483648;
#10;x=-646383648;
#10;x=-646283648;
#10;x=-646183648;
#10;x=-646083648;
#10;x=-645983648;
#10;x=-645883648;
#10;x=-645783648;
#10;x=-645683648;
#10;x=-645583648;
#10;x=-645483648;
#10;x=-645383648;
#10;x=-645283648;
#10;x=-645183648;
#10;x=-645083648;
#10;x=-644983648;
#10;x=-644883648;
#10;x=-644783648;
#10;x=-644683648;
#10;x=-644583648;
#10;x=-644483648;
#10;x=-644383648;
#10;x=-644283648;
#10;x=-644183648;
#10;x=-644083648;
#10;x=-643983648;
#10;x=-643883648;
#10;x=-643783648;
#10;x=-643683648;
#10;x=-643583648;
#10;x=-643483648;
#10;x=-643383648;
#10;x=-643283648;
#10;x=-643183648;
#10;x=-643083648;
#10;x=-642983648;
#10;x=-642883648;
#10;x=-642783648;
#10;x=-642683648;
#10;x=-642583648;
#10;x=-642483648;
#10;x=-642383648;
#10;x=-642283648;
#10;x=-642183648;
#10;x=-642083648;
#10;x=-641983648;
#10;x=-641883648;
#10;x=-641783648;
#10;x=-641683648;
#10;x=-641583648;
#10;x=-641483648;
#10;x=-641383648;
#10;x=-641283648;
#10;x=-641183648;
#10;x=-641083648;
#10;x=-640983648;
#10;x=-640883648;
#10;x=-640783648;
#10;x=-640683648;
#10;x=-640583648;
#10;x=-640483648;
#10;x=-640383648;
#10;x=-640283648;
#10;x=-640183648;
#10;x=-640083648;
#10;x=-639983648;
#10;x=-639883648;
#10;x=-639783648;
#10;x=-639683648;
#10;x=-639583648;
#10;x=-639483648;
#10;x=-639383648;
#10;x=-639283648;
#10;x=-639183648;
#10;x=-639083648;
#10;x=-638983648;
#10;x=-638883648;
#10;x=-638783648;
#10;x=-638683648;
#10;x=-638583648;
#10;x=-638483648;
#10;x=-638383648;
#10;x=-638283648;
#10;x=-638183648;
#10;x=-638083648;
#10;x=-637983648;
#10;x=-637883648;
#10;x=-637783648;
#10;x=-637683648;
#10;x=-637583648;
#10;x=-637483648;
#10;x=-637383648;
#10;x=-637283648;
#10;x=-637183648;
#10;x=-637083648;
#10;x=-636983648;
#10;x=-636883648;
#10;x=-636783648;
#10;x=-636683648;
#10;x=-636583648;
#10;x=-636483648;
#10;x=-636383648;
#10;x=-636283648;
#10;x=-636183648;
#10;x=-636083648;
#10;x=-635983648;
#10;x=-635883648;
#10;x=-635783648;
#10;x=-635683648;
#10;x=-635583648;
#10;x=-635483648;
#10;x=-635383648;
#10;x=-635283648;
#10;x=-635183648;
#10;x=-635083648;
#10;x=-634983648;
#10;x=-634883648;
#10;x=-634783648;
#10;x=-634683648;
#10;x=-634583648;
#10;x=-634483648;
#10;x=-634383648;
#10;x=-634283648;
#10;x=-634183648;
#10;x=-634083648;
#10;x=-633983648;
#10;x=-633883648;
#10;x=-633783648;
#10;x=-633683648;
#10;x=-633583648;
#10;x=-633483648;
#10;x=-633383648;
#10;x=-633283648;
#10;x=-633183648;
#10;x=-633083648;
#10;x=-632983648;
#10;x=-632883648;
#10;x=-632783648;
#10;x=-632683648;
#10;x=-632583648;
#10;x=-632483648;
#10;x=-632383648;
#10;x=-632283648;
#10;x=-632183648;
#10;x=-632083648;
#10;x=-631983648;
#10;x=-631883648;
#10;x=-631783648;
#10;x=-631683648;
#10;x=-631583648;
#10;x=-631483648;
#10;x=-631383648;
#10;x=-631283648;
#10;x=-631183648;
#10;x=-631083648;
#10;x=-630983648;
#10;x=-630883648;
#10;x=-630783648;
#10;x=-630683648;
#10;x=-630583648;
#10;x=-630483648;
#10;x=-630383648;
#10;x=-630283648;
#10;x=-630183648;
#10;x=-630083648;
#10;x=-629983648;
#10;x=-629883648;
#10;x=-629783648;
#10;x=-629683648;
#10;x=-629583648;
#10;x=-629483648;
#10;x=-629383648;
#10;x=-629283648;
#10;x=-629183648;
#10;x=-629083648;
#10;x=-628983648;
#10;x=-628883648;
#10;x=-628783648;
#10;x=-628683648;
#10;x=-628583648;
#10;x=-628483648;
#10;x=-628383648;
#10;x=-628283648;
#10;x=-628183648;
#10;x=-628083648;
#10;x=-627983648;
#10;x=-627883648;
#10;x=-627783648;
#10;x=-627683648;
#10;x=-627583648;
#10;x=-627483648;
#10;x=-627383648;
#10;x=-627283648;
#10;x=-627183648;
#10;x=-627083648;
#10;x=-626983648;
#10;x=-626883648;
#10;x=-626783648;
#10;x=-626683648;
#10;x=-626583648;
#10;x=-626483648;
#10;x=-626383648;
#10;x=-626283648;
#10;x=-626183648;
#10;x=-626083648;
#10;x=-625983648;
#10;x=-625883648;
#10;x=-625783648;
#10;x=-625683648;
#10;x=-625583648;
#10;x=-625483648;
#10;x=-625383648;
#10;x=-625283648;
#10;x=-625183648;
#10;x=-625083648;
#10;x=-624983648;
#10;x=-624883648;
#10;x=-624783648;
#10;x=-624683648;
#10;x=-624583648;
#10;x=-624483648;
#10;x=-624383648;
#10;x=-624283648;
#10;x=-624183648;
#10;x=-624083648;
#10;x=-623983648;
#10;x=-623883648;
#10;x=-623783648;
#10;x=-623683648;
#10;x=-623583648;
#10;x=-623483648;
#10;x=-623383648;
#10;x=-623283648;
#10;x=-623183648;
#10;x=-623083648;
#10;x=-622983648;
#10;x=-622883648;
#10;x=-622783648;
#10;x=-622683648;
#10;x=-622583648;
#10;x=-622483648;
#10;x=-622383648;
#10;x=-622283648;
#10;x=-622183648;
#10;x=-622083648;
#10;x=-621983648;
#10;x=-621883648;
#10;x=-621783648;
#10;x=-621683648;
#10;x=-621583648;
#10;x=-621483648;
#10;x=-621383648;
#10;x=-621283648;
#10;x=-621183648;
#10;x=-621083648;
#10;x=-620983648;
#10;x=-620883648;
#10;x=-620783648;
#10;x=-620683648;
#10;x=-620583648;
#10;x=-620483648;
#10;x=-620383648;
#10;x=-620283648;
#10;x=-620183648;
#10;x=-620083648;
#10;x=-619983648;
#10;x=-619883648;
#10;x=-619783648;
#10;x=-619683648;
#10;x=-619583648;
#10;x=-619483648;
#10;x=-619383648;
#10;x=-619283648;
#10;x=-619183648;
#10;x=-619083648;
#10;x=-618983648;
#10;x=-618883648;
#10;x=-618783648;
#10;x=-618683648;
#10;x=-618583648;
#10;x=-618483648;
#10;x=-618383648;
#10;x=-618283648;
#10;x=-618183648;
#10;x=-618083648;
#10;x=-617983648;
#10;x=-617883648;
#10;x=-617783648;
#10;x=-617683648;
#10;x=-617583648;
#10;x=-617483648;
#10;x=-617383648;
#10;x=-617283648;
#10;x=-617183648;
#10;x=-617083648;
#10;x=-616983648;
#10;x=-616883648;
#10;x=-616783648;
#10;x=-616683648;
#10;x=-616583648;
#10;x=-616483648;
#10;x=-616383648;
#10;x=-616283648;
#10;x=-616183648;
#10;x=-616083648;
#10;x=-615983648;
#10;x=-615883648;
#10;x=-615783648;
#10;x=-615683648;
#10;x=-615583648;
#10;x=-615483648;
#10;x=-615383648;
#10;x=-615283648;
#10;x=-615183648;
#10;x=-615083648;
#10;x=-614983648;
#10;x=-614883648;
#10;x=-614783648;
#10;x=-614683648;
#10;x=-614583648;
#10;x=-614483648;
#10;x=-614383648;
#10;x=-614283648;
#10;x=-614183648;
#10;x=-614083648;
#10;x=-613983648;
#10;x=-613883648;
#10;x=-613783648;
#10;x=-613683648;
#10;x=-613583648;
#10;x=-613483648;
#10;x=-613383648;
#10;x=-613283648;
#10;x=-613183648;
#10;x=-613083648;
#10;x=-612983648;
#10;x=-612883648;
#10;x=-612783648;
#10;x=-612683648;
#10;x=-612583648;
#10;x=-612483648;
#10;x=-612383648;
#10;x=-612283648;
#10;x=-612183648;
#10;x=-612083648;
#10;x=-611983648;
#10;x=-611883648;
#10;x=-611783648;
#10;x=-611683648;
#10;x=-611583648;
#10;x=-611483648;
#10;x=-611383648;
#10;x=-611283648;
#10;x=-611183648;
#10;x=-611083648;
#10;x=-610983648;
#10;x=-610883648;
#10;x=-610783648;
#10;x=-610683648;
#10;x=-610583648;
#10;x=-610483648;
#10;x=-610383648;
#10;x=-610283648;
#10;x=-610183648;
#10;x=-610083648;
#10;x=-609983648;
#10;x=-609883648;
#10;x=-609783648;
#10;x=-609683648;
#10;x=-609583648;
#10;x=-609483648;
#10;x=-609383648;
#10;x=-609283648;
#10;x=-609183648;
#10;x=-609083648;
#10;x=-608983648;
#10;x=-608883648;
#10;x=-608783648;
#10;x=-608683648;
#10;x=-608583648;
#10;x=-608483648;
#10;x=-608383648;
#10;x=-608283648;
#10;x=-608183648;
#10;x=-608083648;
#10;x=-607983648;
#10;x=-607883648;
#10;x=-607783648;
#10;x=-607683648;
#10;x=-607583648;
#10;x=-607483648;
#10;x=-607383648;
#10;x=-607283648;
#10;x=-607183648;
#10;x=-607083648;
#10;x=-606983648;
#10;x=-606883648;
#10;x=-606783648;
#10;x=-606683648;
#10;x=-606583648;
#10;x=-606483648;
#10;x=-606383648;
#10;x=-606283648;
#10;x=-606183648;
#10;x=-606083648;
#10;x=-605983648;
#10;x=-605883648;
#10;x=-605783648;
#10;x=-605683648;
#10;x=-605583648;
#10;x=-605483648;
#10;x=-605383648;
#10;x=-605283648;
#10;x=-605183648;
#10;x=-605083648;
#10;x=-604983648;
#10;x=-604883648;
#10;x=-604783648;
#10;x=-604683648;
#10;x=-604583648;
#10;x=-604483648;
#10;x=-604383648;
#10;x=-604283648;
#10;x=-604183648;
#10;x=-604083648;
#10;x=-603983648;
#10;x=-603883648;
#10;x=-603783648;
#10;x=-603683648;
#10;x=-603583648;
#10;x=-603483648;
#10;x=-603383648;
#10;x=-603283648;
#10;x=-603183648;
#10;x=-603083648;
#10;x=-602983648;
#10;x=-602883648;
#10;x=-602783648;
#10;x=-602683648;
#10;x=-602583648;
#10;x=-602483648;
#10;x=-602383648;
#10;x=-602283648;
#10;x=-602183648;
#10;x=-602083648;
#10;x=-601983648;
#10;x=-601883648;
#10;x=-601783648;
#10;x=-601683648;
#10;x=-601583648;
#10;x=-601483648;
#10;x=-601383648;
#10;x=-601283648;
#10;x=-601183648;
#10;x=-601083648;
#10;x=-600983648;
#10;x=-600883648;
#10;x=-600783648;
#10;x=-600683648;
#10;x=-600583648;
#10;x=-600483648;
#10;x=-600383648;
#10;x=-600283648;
#10;x=-600183648;
#10;x=-600083648;
#10;x=-599983648;
#10;x=-599883648;
#10;x=-599783648;
#10;x=-599683648;
#10;x=-599583648;
#10;x=-599483648;
#10;x=-599383648;
#10;x=-599283648;
#10;x=-599183648;
#10;x=-599083648;
#10;x=-598983648;
#10;x=-598883648;
#10;x=-598783648;
#10;x=-598683648;
#10;x=-598583648;
#10;x=-598483648;
#10;x=-598383648;
#10;x=-598283648;
#10;x=-598183648;
#10;x=-598083648;
#10;x=-597983648;
#10;x=-597883648;
#10;x=-597783648;
#10;x=-597683648;
#10;x=-597583648;
#10;x=-597483648;
#10;x=-597383648;
#10;x=-597283648;
#10;x=-597183648;
#10;x=-597083648;
#10;x=-596983648;
#10;x=-596883648;
#10;x=-596783648;
#10;x=-596683648;
#10;x=-596583648;
#10;x=-596483648;
#10;x=-596383648;
#10;x=-596283648;
#10;x=-596183648;
#10;x=-596083648;
#10;x=-595983648;
#10;x=-595883648;
#10;x=-595783648;
#10;x=-595683648;
#10;x=-595583648;
#10;x=-595483648;
#10;x=-595383648;
#10;x=-595283648;
#10;x=-595183648;
#10;x=-595083648;
#10;x=-594983648;
#10;x=-594883648;
#10;x=-594783648;
#10;x=-594683648;
#10;x=-594583648;
#10;x=-594483648;
#10;x=-594383648;
#10;x=-594283648;
#10;x=-594183648;
#10;x=-594083648;
#10;x=-593983648;
#10;x=-593883648;
#10;x=-593783648;
#10;x=-593683648;
#10;x=-593583648;
#10;x=-593483648;
#10;x=-593383648;
#10;x=-593283648;
#10;x=-593183648;
#10;x=-593083648;
#10;x=-592983648;
#10;x=-592883648;
#10;x=-592783648;
#10;x=-592683648;
#10;x=-592583648;
#10;x=-592483648;
#10;x=-592383648;
#10;x=-592283648;
#10;x=-592183648;
#10;x=-592083648;
#10;x=-591983648;
#10;x=-591883648;
#10;x=-591783648;
#10;x=-591683648;
#10;x=-591583648;
#10;x=-591483648;
#10;x=-591383648;
#10;x=-591283648;
#10;x=-591183648;
#10;x=-591083648;
#10;x=-590983648;
#10;x=-590883648;
#10;x=-590783648;
#10;x=-590683648;
#10;x=-590583648;
#10;x=-590483648;
#10;x=-590383648;
#10;x=-590283648;
#10;x=-590183648;
#10;x=-590083648;
#10;x=-589983648;
#10;x=-589883648;
#10;x=-589783648;
#10;x=-589683648;
#10;x=-589583648;
#10;x=-589483648;
#10;x=-589383648;
#10;x=-589283648;
#10;x=-589183648;
#10;x=-589083648;
#10;x=-588983648;
#10;x=-588883648;
#10;x=-588783648;
#10;x=-588683648;
#10;x=-588583648;
#10;x=-588483648;
#10;x=-588383648;
#10;x=-588283648;
#10;x=-588183648;
#10;x=-588083648;
#10;x=-587983648;
#10;x=-587883648;
#10;x=-587783648;
#10;x=-587683648;
#10;x=-587583648;
#10;x=-587483648;
#10;x=-587383648;
#10;x=-587283648;
#10;x=-587183648;
#10;x=-587083648;
#10;x=-586983648;
#10;x=-586883648;
#10;x=-586783648;
#10;x=-586683648;
#10;x=-586583648;
#10;x=-586483648;
#10;x=-586383648;
#10;x=-586283648;
#10;x=-586183648;
#10;x=-586083648;
#10;x=-585983648;
#10;x=-585883648;
#10;x=-585783648;
#10;x=-585683648;
#10;x=-585583648;
#10;x=-585483648;
#10;x=-585383648;
#10;x=-585283648;
#10;x=-585183648;
#10;x=-585083648;
#10;x=-584983648;
#10;x=-584883648;
#10;x=-584783648;
#10;x=-584683648;
#10;x=-584583648;
#10;x=-584483648;
#10;x=-584383648;
#10;x=-584283648;
#10;x=-584183648;
#10;x=-584083648;
#10;x=-583983648;
#10;x=-583883648;
#10;x=-583783648;
#10;x=-583683648;
#10;x=-583583648;
#10;x=-583483648;
#10;x=-583383648;
#10;x=-583283648;
#10;x=-583183648;
#10;x=-583083648;
#10;x=-582983648;
#10;x=-582883648;
#10;x=-582783648;
#10;x=-582683648;
#10;x=-582583648;
#10;x=-582483648;
#10;x=-582383648;
#10;x=-582283648;
#10;x=-582183648;
#10;x=-582083648;
#10;x=-581983648;
#10;x=-581883648;
#10;x=-581783648;
#10;x=-581683648;
#10;x=-581583648;
#10;x=-581483648;
#10;x=-581383648;
#10;x=-581283648;
#10;x=-581183648;
#10;x=-581083648;
#10;x=-580983648;
#10;x=-580883648;
#10;x=-580783648;
#10;x=-580683648;
#10;x=-580583648;
#10;x=-580483648;
#10;x=-580383648;
#10;x=-580283648;
#10;x=-580183648;
#10;x=-580083648;
#10;x=-579983648;
#10;x=-579883648;
#10;x=-579783648;
#10;x=-579683648;
#10;x=-579583648;
#10;x=-579483648;
#10;x=-579383648;
#10;x=-579283648;
#10;x=-579183648;
#10;x=-579083648;
#10;x=-578983648;
#10;x=-578883648;
#10;x=-578783648;
#10;x=-578683648;
#10;x=-578583648;
#10;x=-578483648;
#10;x=-578383648;
#10;x=-578283648;
#10;x=-578183648;
#10;x=-578083648;
#10;x=-577983648;
#10;x=-577883648;
#10;x=-577783648;
#10;x=-577683648;
#10;x=-577583648;
#10;x=-577483648;
#10;x=-577383648;
#10;x=-577283648;
#10;x=-577183648;
#10;x=-577083648;
#10;x=-576983648;
#10;x=-576883648;
#10;x=-576783648;
#10;x=-576683648;
#10;x=-576583648;
#10;x=-576483648;
#10;x=-576383648;
#10;x=-576283648;
#10;x=-576183648;
#10;x=-576083648;
#10;x=-575983648;
#10;x=-575883648;
#10;x=-575783648;
#10;x=-575683648;
#10;x=-575583648;
#10;x=-575483648;
#10;x=-575383648;
#10;x=-575283648;
#10;x=-575183648;
#10;x=-575083648;
#10;x=-574983648;
#10;x=-574883648;
#10;x=-574783648;
#10;x=-574683648;
#10;x=-574583648;
#10;x=-574483648;
#10;x=-574383648;
#10;x=-574283648;
#10;x=-574183648;
#10;x=-574083648;
#10;x=-573983648;
#10;x=-573883648;
#10;x=-573783648;
#10;x=-573683648;
#10;x=-573583648;
#10;x=-573483648;
#10;x=-573383648;
#10;x=-573283648;
#10;x=-573183648;
#10;x=-573083648;
#10;x=-572983648;
#10;x=-572883648;
#10;x=-572783648;
#10;x=-572683648;
#10;x=-572583648;
#10;x=-572483648;
#10;x=-572383648;
#10;x=-572283648;
#10;x=-572183648;
#10;x=-572083648;
#10;x=-571983648;
#10;x=-571883648;
#10;x=-571783648;
#10;x=-571683648;
#10;x=-571583648;
#10;x=-571483648;
#10;x=-571383648;
#10;x=-571283648;
#10;x=-571183648;
#10;x=-571083648;
#10;x=-570983648;
#10;x=-570883648;
#10;x=-570783648;
#10;x=-570683648;
#10;x=-570583648;
#10;x=-570483648;
#10;x=-570383648;
#10;x=-570283648;
#10;x=-570183648;
#10;x=-570083648;
#10;x=-569983648;
#10;x=-569883648;
#10;x=-569783648;
#10;x=-569683648;
#10;x=-569583648;
#10;x=-569483648;
#10;x=-569383648;
#10;x=-569283648;
#10;x=-569183648;
#10;x=-569083648;
#10;x=-568983648;
#10;x=-568883648;
#10;x=-568783648;
#10;x=-568683648;
#10;x=-568583648;
#10;x=-568483648;
#10;x=-568383648;
#10;x=-568283648;
#10;x=-568183648;
#10;x=-568083648;
#10;x=-567983648;
#10;x=-567883648;
#10;x=-567783648;
#10;x=-567683648;
#10;x=-567583648;
#10;x=-567483648;
#10;x=-567383648;
#10;x=-567283648;
#10;x=-567183648;
#10;x=-567083648;
#10;x=-566983648;
#10;x=-566883648;
#10;x=-566783648;
#10;x=-566683648;
#10;x=-566583648;
#10;x=-566483648;
#10;x=-566383648;
#10;x=-566283648;
#10;x=-566183648;
#10;x=-566083648;
#10;x=-565983648;
#10;x=-565883648;
#10;x=-565783648;
#10;x=-565683648;
#10;x=-565583648;
#10;x=-565483648;
#10;x=-565383648;
#10;x=-565283648;
#10;x=-565183648;
#10;x=-565083648;
#10;x=-564983648;
#10;x=-564883648;
#10;x=-564783648;
#10;x=-564683648;
#10;x=-564583648;
#10;x=-564483648;
#10;x=-564383648;
#10;x=-564283648;
#10;x=-564183648;
#10;x=-564083648;
#10;x=-563983648;
#10;x=-563883648;
#10;x=-563783648;
#10;x=-563683648;
#10;x=-563583648;
#10;x=-563483648;
#10;x=-563383648;
#10;x=-563283648;
#10;x=-563183648;
#10;x=-563083648;
#10;x=-562983648;
#10;x=-562883648;
#10;x=-562783648;
#10;x=-562683648;
#10;x=-562583648;
#10;x=-562483648;
#10;x=-562383648;
#10;x=-562283648;
#10;x=-562183648;
#10;x=-562083648;
#10;x=-561983648;
#10;x=-561883648;
#10;x=-561783648;
#10;x=-561683648;
#10;x=-561583648;
#10;x=-561483648;
#10;x=-561383648;
#10;x=-561283648;
#10;x=-561183648;
#10;x=-561083648;
#10;x=-560983648;
#10;x=-560883648;
#10;x=-560783648;
#10;x=-560683648;
#10;x=-560583648;
#10;x=-560483648;
#10;x=-560383648;
#10;x=-560283648;
#10;x=-560183648;
#10;x=-560083648;
#10;x=-559983648;
#10;x=-559883648;
#10;x=-559783648;
#10;x=-559683648;
#10;x=-559583648;
#10;x=-559483648;
#10;x=-559383648;
#10;x=-559283648;
#10;x=-559183648;
#10;x=-559083648;
#10;x=-558983648;
#10;x=-558883648;
#10;x=-558783648;
#10;x=-558683648;
#10;x=-558583648;
#10;x=-558483648;
#10;x=-558383648;
#10;x=-558283648;
#10;x=-558183648;
#10;x=-558083648;
#10;x=-557983648;
#10;x=-557883648;
#10;x=-557783648;
#10;x=-557683648;
#10;x=-557583648;
#10;x=-557483648;
#10;x=-557383648;
#10;x=-557283648;
#10;x=-557183648;
#10;x=-557083648;
#10;x=-556983648;
#10;x=-556883648;
#10;x=-556783648;
#10;x=-556683648;
#10;x=-556583648;
#10;x=-556483648;
#10;x=-556383648;
#10;x=-556283648;
#10;x=-556183648;
#10;x=-556083648;
#10;x=-555983648;
#10;x=-555883648;
#10;x=-555783648;
#10;x=-555683648;
#10;x=-555583648;
#10;x=-555483648;
#10;x=-555383648;
#10;x=-555283648;
#10;x=-555183648;
#10;x=-555083648;
#10;x=-554983648;
#10;x=-554883648;
#10;x=-554783648;
#10;x=-554683648;
#10;x=-554583648;
#10;x=-554483648;
#10;x=-554383648;
#10;x=-554283648;
#10;x=-554183648;
#10;x=-554083648;
#10;x=-553983648;
#10;x=-553883648;
#10;x=-553783648;
#10;x=-553683648;
#10;x=-553583648;
#10;x=-553483648;
#10;x=-553383648;
#10;x=-553283648;
#10;x=-553183648;
#10;x=-553083648;
#10;x=-552983648;
#10;x=-552883648;
#10;x=-552783648;
#10;x=-552683648;
#10;x=-552583648;
#10;x=-552483648;
#10;x=-552383648;
#10;x=-552283648;
#10;x=-552183648;
#10;x=-552083648;
#10;x=-551983648;
#10;x=-551883648;
#10;x=-551783648;
#10;x=-551683648;
#10;x=-551583648;
#10;x=-551483648;
#10;x=-551383648;
#10;x=-551283648;
#10;x=-551183648;
#10;x=-551083648;
#10;x=-550983648;
#10;x=-550883648;
#10;x=-550783648;
#10;x=-550683648;
#10;x=-550583648;
#10;x=-550483648;
#10;x=-550383648;
#10;x=-550283648;
#10;x=-550183648;
#10;x=-550083648;
#10;x=-549983648;
#10;x=-549883648;
#10;x=-549783648;
#10;x=-549683648;
#10;x=-549583648;
#10;x=-549483648;
#10;x=-549383648;
#10;x=-549283648;
#10;x=-549183648;
#10;x=-549083648;
#10;x=-548983648;
#10;x=-548883648;
#10;x=-548783648;
#10;x=-548683648;
#10;x=-548583648;
#10;x=-548483648;
#10;x=-548383648;
#10;x=-548283648;
#10;x=-548183648;
#10;x=-548083648;
#10;x=-547983648;
#10;x=-547883648;
#10;x=-547783648;
#10;x=-547683648;
#10;x=-547583648;
#10;x=-547483648;
#10;x=-547383648;
#10;x=-547283648;
#10;x=-547183648;
#10;x=-547083648;
#10;x=-546983648;
#10;x=-546883648;
#10;x=-546783648;
#10;x=-546683648;
#10;x=-546583648;
#10;x=-546483648;
#10;x=-546383648;
#10;x=-546283648;
#10;x=-546183648;
#10;x=-546083648;
#10;x=-545983648;
#10;x=-545883648;
#10;x=-545783648;
#10;x=-545683648;
#10;x=-545583648;
#10;x=-545483648;
#10;x=-545383648;
#10;x=-545283648;
#10;x=-545183648;
#10;x=-545083648;
#10;x=-544983648;
#10;x=-544883648;
#10;x=-544783648;
#10;x=-544683648;
#10;x=-544583648;
#10;x=-544483648;
#10;x=-544383648;
#10;x=-544283648;
#10;x=-544183648;
#10;x=-544083648;
#10;x=-543983648;
#10;x=-543883648;
#10;x=-543783648;
#10;x=-543683648;
#10;x=-543583648;
#10;x=-543483648;
#10;x=-543383648;
#10;x=-543283648;
#10;x=-543183648;
#10;x=-543083648;
#10;x=-542983648;
#10;x=-542883648;
#10;x=-542783648;
#10;x=-542683648;
#10;x=-542583648;
#10;x=-542483648;
#10;x=-542383648;
#10;x=-542283648;
#10;x=-542183648;
#10;x=-542083648;
#10;x=-541983648;
#10;x=-541883648;
#10;x=-541783648;
#10;x=-541683648;
#10;x=-541583648;
#10;x=-541483648;
#10;x=-541383648;
#10;x=-541283648;
#10;x=-541183648;
#10;x=-541083648;
#10;x=-540983648;
#10;x=-540883648;
#10;x=-540783648;
#10;x=-540683648;
#10;x=-540583648;
#10;x=-540483648;
#10;x=-540383648;
#10;x=-540283648;
#10;x=-540183648;
#10;x=-540083648;
#10;x=-539983648;
#10;x=-539883648;
#10;x=-539783648;
#10;x=-539683648;
#10;x=-539583648;
#10;x=-539483648;
#10;x=-539383648;
#10;x=-539283648;
#10;x=-539183648;
#10;x=-539083648;
#10;x=-538983648;
#10;x=-538883648;
#10;x=-538783648;
#10;x=-538683648;
#10;x=-538583648;
#10;x=-538483648;
#10;x=-538383648;
#10;x=-538283648;
#10;x=-538183648;
#10;x=-538083648;
#10;x=-537983648;
#10;x=-537883648;
#10;x=-537783648;
#10;x=-537683648;
#10;x=-537583648;
#10;x=-537483648;
#10;x=-537383648;
#10;x=-537283648;
#10;x=-537183648;
#10;x=-537083648;
#10;x=-536983648;
#10;x=-536883648;
#10;x=-536783648;
#10;x=-536683648;
#10;x=-536583648;
#10;x=-536483648;
#10;x=-536383648;
#10;x=-536283648;
#10;x=-536183648;
#10;x=-536083648;
#10;x=-535983648;
#10;x=-535883648;
#10;x=-535783648;
#10;x=-535683648;
#10;x=-535583648;
#10;x=-535483648;
#10;x=-535383648;
#10;x=-535283648;
#10;x=-535183648;
#10;x=-535083648;
#10;x=-534983648;
#10;x=-534883648;
#10;x=-534783648;
#10;x=-534683648;
#10;x=-534583648;
#10;x=-534483648;
#10;x=-534383648;
#10;x=-534283648;
#10;x=-534183648;
#10;x=-534083648;
#10;x=-533983648;
#10;x=-533883648;
#10;x=-533783648;
#10;x=-533683648;
#10;x=-533583648;
#10;x=-533483648;
#10;x=-533383648;
#10;x=-533283648;
#10;x=-533183648;
#10;x=-533083648;
#10;x=-532983648;
#10;x=-532883648;
#10;x=-532783648;
#10;x=-532683648;
#10;x=-532583648;
#10;x=-532483648;
#10;x=-532383648;
#10;x=-532283648;
#10;x=-532183648;
#10;x=-532083648;
#10;x=-531983648;
#10;x=-531883648;
#10;x=-531783648;
#10;x=-531683648;
#10;x=-531583648;
#10;x=-531483648;
#10;x=-531383648;
#10;x=-531283648;
#10;x=-531183648;
#10;x=-531083648;
#10;x=-530983648;
#10;x=-530883648;
#10;x=-530783648;
#10;x=-530683648;
#10;x=-530583648;
#10;x=-530483648;
#10;x=-530383648;
#10;x=-530283648;
#10;x=-530183648;
#10;x=-530083648;
#10;x=-529983648;
#10;x=-529883648;
#10;x=-529783648;
#10;x=-529683648;
#10;x=-529583648;
#10;x=-529483648;
#10;x=-529383648;
#10;x=-529283648;
#10;x=-529183648;
#10;x=-529083648;
#10;x=-528983648;
#10;x=-528883648;
#10;x=-528783648;
#10;x=-528683648;
#10;x=-528583648;
#10;x=-528483648;
#10;x=-528383648;
#10;x=-528283648;
#10;x=-528183648;
#10;x=-528083648;
#10;x=-527983648;
#10;x=-527883648;
#10;x=-527783648;
#10;x=-527683648;
#10;x=-527583648;
#10;x=-527483648;
#10;x=-527383648;
#10;x=-527283648;
#10;x=-527183648;
#10;x=-527083648;
#10;x=-526983648;
#10;x=-526883648;
#10;x=-526783648;
#10;x=-526683648;
#10;x=-526583648;
#10;x=-526483648;
#10;x=-526383648;
#10;x=-526283648;
#10;x=-526183648;
#10;x=-526083648;
#10;x=-525983648;
#10;x=-525883648;
#10;x=-525783648;
#10;x=-525683648;
#10;x=-525583648;
#10;x=-525483648;
#10;x=-525383648;
#10;x=-525283648;
#10;x=-525183648;
#10;x=-525083648;
#10;x=-524983648;
#10;x=-524883648;
#10;x=-524783648;
#10;x=-524683648;
#10;x=-524583648;
#10;x=-524483648;
#10;x=-524383648;
#10;x=-524283648;
#10;x=-524183648;
#10;x=-524083648;
#10;x=-523983648;
#10;x=-523883648;
#10;x=-523783648;
#10;x=-523683648;
#10;x=-523583648;
#10;x=-523483648;
#10;x=-523383648;
#10;x=-523283648;
#10;x=-523183648;
#10;x=-523083648;
#10;x=-522983648;
#10;x=-522883648;
#10;x=-522783648;
#10;x=-522683648;
#10;x=-522583648;
#10;x=-522483648;
#10;x=-522383648;
#10;x=-522283648;
#10;x=-522183648;
#10;x=-522083648;
#10;x=-521983648;
#10;x=-521883648;
#10;x=-521783648;
#10;x=-521683648;
#10;x=-521583648;
#10;x=-521483648;
#10;x=-521383648;
#10;x=-521283648;
#10;x=-521183648;
#10;x=-521083648;
#10;x=-520983648;
#10;x=-520883648;
#10;x=-520783648;
#10;x=-520683648;
#10;x=-520583648;
#10;x=-520483648;
#10;x=-520383648;
#10;x=-520283648;
#10;x=-520183648;
#10;x=-520083648;
#10;x=-519983648;
#10;x=-519883648;
#10;x=-519783648;
#10;x=-519683648;
#10;x=-519583648;
#10;x=-519483648;
#10;x=-519383648;
#10;x=-519283648;
#10;x=-519183648;
#10;x=-519083648;
#10;x=-518983648;
#10;x=-518883648;
#10;x=-518783648;
#10;x=-518683648;
#10;x=-518583648;
#10;x=-518483648;
#10;x=-518383648;
#10;x=-518283648;
#10;x=-518183648;
#10;x=-518083648;
#10;x=-517983648;
#10;x=-517883648;
#10;x=-517783648;
#10;x=-517683648;
#10;x=-517583648;
#10;x=-517483648;
#10;x=-517383648;
#10;x=-517283648;
#10;x=-517183648;
#10;x=-517083648;
#10;x=-516983648;
#10;x=-516883648;
#10;x=-516783648;
#10;x=-516683648;
#10;x=-516583648;
#10;x=-516483648;
#10;x=-516383648;
#10;x=-516283648;
#10;x=-516183648;
#10;x=-516083648;
#10;x=-515983648;
#10;x=-515883648;
#10;x=-515783648;
#10;x=-515683648;
#10;x=-515583648;
#10;x=-515483648;
#10;x=-515383648;
#10;x=-515283648;
#10;x=-515183648;
#10;x=-515083648;
#10;x=-514983648;
#10;x=-514883648;
#10;x=-514783648;
#10;x=-514683648;
#10;x=-514583648;
#10;x=-514483648;
#10;x=-514383648;
#10;x=-514283648;
#10;x=-514183648;
#10;x=-514083648;
#10;x=-513983648;
#10;x=-513883648;
#10;x=-513783648;
#10;x=-513683648;
#10;x=-513583648;
#10;x=-513483648;
#10;x=-513383648;
#10;x=-513283648;
#10;x=-513183648;
#10;x=-513083648;
#10;x=-512983648;
#10;x=-512883648;
#10;x=-512783648;
#10;x=-512683648;
#10;x=-512583648;
#10;x=-512483648;
#10;x=-512383648;
#10;x=-512283648;
#10;x=-512183648;
#10;x=-512083648;
#10;x=-511983648;
#10;x=-511883648;
#10;x=-511783648;
#10;x=-511683648;
#10;x=-511583648;
#10;x=-511483648;
#10;x=-511383648;
#10;x=-511283648;
#10;x=-511183648;
#10;x=-511083648;
#10;x=-510983648;
#10;x=-510883648;
#10;x=-510783648;
#10;x=-510683648;
#10;x=-510583648;
#10;x=-510483648;
#10;x=-510383648;
#10;x=-510283648;
#10;x=-510183648;
#10;x=-510083648;
#10;x=-509983648;
#10;x=-509883648;
#10;x=-509783648;
#10;x=-509683648;
#10;x=-509583648;
#10;x=-509483648;
#10;x=-509383648;
#10;x=-509283648;
#10;x=-509183648;
#10;x=-509083648;
#10;x=-508983648;
#10;x=-508883648;
#10;x=-508783648;
#10;x=-508683648;
#10;x=-508583648;
#10;x=-508483648;
#10;x=-508383648;
#10;x=-508283648;
#10;x=-508183648;
#10;x=-508083648;
#10;x=-507983648;
#10;x=-507883648;
#10;x=-507783648;
#10;x=-507683648;
#10;x=-507583648;
#10;x=-507483648;
#10;x=-507383648;
#10;x=-507283648;
#10;x=-507183648;
#10;x=-507083648;
#10;x=-506983648;
#10;x=-506883648;
#10;x=-506783648;
#10;x=-506683648;
#10;x=-506583648;
#10;x=-506483648;
#10;x=-506383648;
#10;x=-506283648;
#10;x=-506183648;
#10;x=-506083648;
#10;x=-505983648;
#10;x=-505883648;
#10;x=-505783648;
#10;x=-505683648;
#10;x=-505583648;
#10;x=-505483648;
#10;x=-505383648;
#10;x=-505283648;
#10;x=-505183648;
#10;x=-505083648;
#10;x=-504983648;
#10;x=-504883648;
#10;x=-504783648;
#10;x=-504683648;
#10;x=-504583648;
#10;x=-504483648;
#10;x=-504383648;
#10;x=-504283648;
#10;x=-504183648;
#10;x=-504083648;
#10;x=-503983648;
#10;x=-503883648;
#10;x=-503783648;
#10;x=-503683648;
#10;x=-503583648;
#10;x=-503483648;
#10;x=-503383648;
#10;x=-503283648;
#10;x=-503183648;
#10;x=-503083648;
#10;x=-502983648;
#10;x=-502883648;
#10;x=-502783648;
#10;x=-502683648;
#10;x=-502583648;
#10;x=-502483648;
#10;x=-502383648;
#10;x=-502283648;
#10;x=-502183648;
#10;x=-502083648;
#10;x=-501983648;
#10;x=-501883648;
#10;x=-501783648;
#10;x=-501683648;
#10;x=-501583648;
#10;x=-501483648;
#10;x=-501383648;
#10;x=-501283648;
#10;x=-501183648;
#10;x=-501083648;
#10;x=-500983648;
#10;x=-500883648;
#10;x=-500783648;
#10;x=-500683648;
#10;x=-500583648;
#10;x=-500483648;
#10;x=-500383648;
#10;x=-500283648;
#10;x=-500183648;
#10;x=-500083648;
#10;x=-499983648;
#10;x=-499883648;
#10;x=-499783648;
#10;x=-499683648;
#10;x=-499583648;
#10;x=-499483648;
#10;x=-499383648;
#10;x=-499283648;
#10;x=-499183648;
#10;x=-499083648;
#10;x=-498983648;
#10;x=-498883648;
#10;x=-498783648;
#10;x=-498683648;
#10;x=-498583648;
#10;x=-498483648;
#10;x=-498383648;
#10;x=-498283648;
#10;x=-498183648;
#10;x=-498083648;
#10;x=-497983648;
#10;x=-497883648;
#10;x=-497783648;
#10;x=-497683648;
#10;x=-497583648;
#10;x=-497483648;
#10;x=-497383648;
#10;x=-497283648;
#10;x=-497183648;
#10;x=-497083648;
#10;x=-496983648;
#10;x=-496883648;
#10;x=-496783648;
#10;x=-496683648;
#10;x=-496583648;
#10;x=-496483648;
#10;x=-496383648;
#10;x=-496283648;
#10;x=-496183648;
#10;x=-496083648;
#10;x=-495983648;
#10;x=-495883648;
#10;x=-495783648;
#10;x=-495683648;
#10;x=-495583648;
#10;x=-495483648;
#10;x=-495383648;
#10;x=-495283648;
#10;x=-495183648;
#10;x=-495083648;
#10;x=-494983648;
#10;x=-494883648;
#10;x=-494783648;
#10;x=-494683648;
#10;x=-494583648;
#10;x=-494483648;
#10;x=-494383648;
#10;x=-494283648;
#10;x=-494183648;
#10;x=-494083648;
#10;x=-493983648;
#10;x=-493883648;
#10;x=-493783648;
#10;x=-493683648;
#10;x=-493583648;
#10;x=-493483648;
#10;x=-493383648;
#10;x=-493283648;
#10;x=-493183648;
#10;x=-493083648;
#10;x=-492983648;
#10;x=-492883648;
#10;x=-492783648;
#10;x=-492683648;
#10;x=-492583648;
#10;x=-492483648;
#10;x=-492383648;
#10;x=-492283648;
#10;x=-492183648;
#10;x=-492083648;
#10;x=-491983648;
#10;x=-491883648;
#10;x=-491783648;
#10;x=-491683648;
#10;x=-491583648;
#10;x=-491483648;
#10;x=-491383648;
#10;x=-491283648;
#10;x=-491183648;
#10;x=-491083648;
#10;x=-490983648;
#10;x=-490883648;
#10;x=-490783648;
#10;x=-490683648;
#10;x=-490583648;
#10;x=-490483648;
#10;x=-490383648;
#10;x=-490283648;
#10;x=-490183648;
#10;x=-490083648;
#10;x=-489983648;
#10;x=-489883648;
#10;x=-489783648;
#10;x=-489683648;
#10;x=-489583648;
#10;x=-489483648;
#10;x=-489383648;
#10;x=-489283648;
#10;x=-489183648;
#10;x=-489083648;
#10;x=-488983648;
#10;x=-488883648;
#10;x=-488783648;
#10;x=-488683648;
#10;x=-488583648;
#10;x=-488483648;
#10;x=-488383648;
#10;x=-488283648;
#10;x=-488183648;
#10;x=-488083648;
#10;x=-487983648;
#10;x=-487883648;
#10;x=-487783648;
#10;x=-487683648;
#10;x=-487583648;
#10;x=-487483648;
#10;x=-487383648;
#10;x=-487283648;
#10;x=-487183648;
#10;x=-487083648;
#10;x=-486983648;
#10;x=-486883648;
#10;x=-486783648;
#10;x=-486683648;
#10;x=-486583648;
#10;x=-486483648;
#10;x=-486383648;
#10;x=-486283648;
#10;x=-486183648;
#10;x=-486083648;
#10;x=-485983648;
#10;x=-485883648;
#10;x=-485783648;
#10;x=-485683648;
#10;x=-485583648;
#10;x=-485483648;
#10;x=-485383648;
#10;x=-485283648;
#10;x=-485183648;
#10;x=-485083648;
#10;x=-484983648;
#10;x=-484883648;
#10;x=-484783648;
#10;x=-484683648;
#10;x=-484583648;
#10;x=-484483648;
#10;x=-484383648;
#10;x=-484283648;
#10;x=-484183648;
#10;x=-484083648;
#10;x=-483983648;
#10;x=-483883648;
#10;x=-483783648;
#10;x=-483683648;
#10;x=-483583648;
#10;x=-483483648;
#10;x=-483383648;
#10;x=-483283648;
#10;x=-483183648;
#10;x=-483083648;
#10;x=-482983648;
#10;x=-482883648;
#10;x=-482783648;
#10;x=-482683648;
#10;x=-482583648;
#10;x=-482483648;
#10;x=-482383648;
#10;x=-482283648;
#10;x=-482183648;
#10;x=-482083648;
#10;x=-481983648;
#10;x=-481883648;
#10;x=-481783648;
#10;x=-481683648;
#10;x=-481583648;
#10;x=-481483648;
#10;x=-481383648;
#10;x=-481283648;
#10;x=-481183648;
#10;x=-481083648;
#10;x=-480983648;
#10;x=-480883648;
#10;x=-480783648;
#10;x=-480683648;
#10;x=-480583648;
#10;x=-480483648;
#10;x=-480383648;
#10;x=-480283648;
#10;x=-480183648;
#10;x=-480083648;
#10;x=-479983648;
#10;x=-479883648;
#10;x=-479783648;
#10;x=-479683648;
#10;x=-479583648;
#10;x=-479483648;
#10;x=-479383648;
#10;x=-479283648;
#10;x=-479183648;
#10;x=-479083648;
#10;x=-478983648;
#10;x=-478883648;
#10;x=-478783648;
#10;x=-478683648;
#10;x=-478583648;
#10;x=-478483648;
#10;x=-478383648;
#10;x=-478283648;
#10;x=-478183648;
#10;x=-478083648;
#10;x=-477983648;
#10;x=-477883648;
#10;x=-477783648;
#10;x=-477683648;
#10;x=-477583648;
#10;x=-477483648;
#10;x=-477383648;
#10;x=-477283648;
#10;x=-477183648;
#10;x=-477083648;
#10;x=-476983648;
#10;x=-476883648;
#10;x=-476783648;
#10;x=-476683648;
#10;x=-476583648;
#10;x=-476483648;
#10;x=-476383648;
#10;x=-476283648;
#10;x=-476183648;
#10;x=-476083648;
#10;x=-475983648;
#10;x=-475883648;
#10;x=-475783648;
#10;x=-475683648;
#10;x=-475583648;
#10;x=-475483648;
#10;x=-475383648;
#10;x=-475283648;
#10;x=-475183648;
#10;x=-475083648;
#10;x=-474983648;
#10;x=-474883648;
#10;x=-474783648;
#10;x=-474683648;
#10;x=-474583648;
#10;x=-474483648;
#10;x=-474383648;
#10;x=-474283648;
#10;x=-474183648;
#10;x=-474083648;
#10;x=-473983648;
#10;x=-473883648;
#10;x=-473783648;
#10;x=-473683648;
#10;x=-473583648;
#10;x=-473483648;
#10;x=-473383648;
#10;x=-473283648;
#10;x=-473183648;
#10;x=-473083648;
#10;x=-472983648;
#10;x=-472883648;
#10;x=-472783648;
#10;x=-472683648;
#10;x=-472583648;
#10;x=-472483648;
#10;x=-472383648;
#10;x=-472283648;
#10;x=-472183648;
#10;x=-472083648;
#10;x=-471983648;
#10;x=-471883648;
#10;x=-471783648;
#10;x=-471683648;
#10;x=-471583648;
#10;x=-471483648;
#10;x=-471383648;
#10;x=-471283648;
#10;x=-471183648;
#10;x=-471083648;
#10;x=-470983648;
#10;x=-470883648;
#10;x=-470783648;
#10;x=-470683648;
#10;x=-470583648;
#10;x=-470483648;
#10;x=-470383648;
#10;x=-470283648;
#10;x=-470183648;
#10;x=-470083648;
#10;x=-469983648;
#10;x=-469883648;
#10;x=-469783648;
#10;x=-469683648;
#10;x=-469583648;
#10;x=-469483648;
#10;x=-469383648;
#10;x=-469283648;
#10;x=-469183648;
#10;x=-469083648;
#10;x=-468983648;
#10;x=-468883648;
#10;x=-468783648;
#10;x=-468683648;
#10;x=-468583648;
#10;x=-468483648;
#10;x=-468383648;
#10;x=-468283648;
#10;x=-468183648;
#10;x=-468083648;
#10;x=-467983648;
#10;x=-467883648;
#10;x=-467783648;
#10;x=-467683648;
#10;x=-467583648;
#10;x=-467483648;
#10;x=-467383648;
#10;x=-467283648;
#10;x=-467183648;
#10;x=-467083648;
#10;x=-466983648;
#10;x=-466883648;
#10;x=-466783648;
#10;x=-466683648;
#10;x=-466583648;
#10;x=-466483648;
#10;x=-466383648;
#10;x=-466283648;
#10;x=-466183648;
#10;x=-466083648;
#10;x=-465983648;
#10;x=-465883648;
#10;x=-465783648;
#10;x=-465683648;
#10;x=-465583648;
#10;x=-465483648;
#10;x=-465383648;
#10;x=-465283648;
#10;x=-465183648;
#10;x=-465083648;
#10;x=-464983648;
#10;x=-464883648;
#10;x=-464783648;
#10;x=-464683648;
#10;x=-464583648;
#10;x=-464483648;
#10;x=-464383648;
#10;x=-464283648;
#10;x=-464183648;
#10;x=-464083648;
#10;x=-463983648;
#10;x=-463883648;
#10;x=-463783648;
#10;x=-463683648;
#10;x=-463583648;
#10;x=-463483648;
#10;x=-463383648;
#10;x=-463283648;
#10;x=-463183648;
#10;x=-463083648;
#10;x=-462983648;
#10;x=-462883648;
#10;x=-462783648;
#10;x=-462683648;
#10;x=-462583648;
#10;x=-462483648;
#10;x=-462383648;
#10;x=-462283648;
#10;x=-462183648;
#10;x=-462083648;
#10;x=-461983648;
#10;x=-461883648;
#10;x=-461783648;
#10;x=-461683648;
#10;x=-461583648;
#10;x=-461483648;
#10;x=-461383648;
#10;x=-461283648;
#10;x=-461183648;
#10;x=-461083648;
#10;x=-460983648;
#10;x=-460883648;
#10;x=-460783648;
#10;x=-460683648;
#10;x=-460583648;
#10;x=-460483648;
#10;x=-460383648;
#10;x=-460283648;
#10;x=-460183648;
#10;x=-460083648;
#10;x=-459983648;
#10;x=-459883648;
#10;x=-459783648;
#10;x=-459683648;
#10;x=-459583648;
#10;x=-459483648;
#10;x=-459383648;
#10;x=-459283648;
#10;x=-459183648;
#10;x=-459083648;
#10;x=-458983648;
#10;x=-458883648;
#10;x=-458783648;
#10;x=-458683648;
#10;x=-458583648;
#10;x=-458483648;
#10;x=-458383648;
#10;x=-458283648;
#10;x=-458183648;
#10;x=-458083648;
#10;x=-457983648;
#10;x=-457883648;
#10;x=-457783648;
#10;x=-457683648;
#10;x=-457583648;
#10;x=-457483648;
#10;x=-457383648;
#10;x=-457283648;
#10;x=-457183648;
#10;x=-457083648;
#10;x=-456983648;
#10;x=-456883648;
#10;x=-456783648;
#10;x=-456683648;
#10;x=-456583648;
#10;x=-456483648;
#10;x=-456383648;
#10;x=-456283648;
#10;x=-456183648;
#10;x=-456083648;
#10;x=-455983648;
#10;x=-455883648;
#10;x=-455783648;
#10;x=-455683648;
#10;x=-455583648;
#10;x=-455483648;
#10;x=-455383648;
#10;x=-455283648;
#10;x=-455183648;
#10;x=-455083648;
#10;x=-454983648;
#10;x=-454883648;
#10;x=-454783648;
#10;x=-454683648;
#10;x=-454583648;
#10;x=-454483648;
#10;x=-454383648;
#10;x=-454283648;
#10;x=-454183648;
#10;x=-454083648;
#10;x=-453983648;
#10;x=-453883648;
#10;x=-453783648;
#10;x=-453683648;
#10;x=-453583648;
#10;x=-453483648;
#10;x=-453383648;
#10;x=-453283648;
#10;x=-453183648;
#10;x=-453083648;
#10;x=-452983648;
#10;x=-452883648;
#10;x=-452783648;
#10;x=-452683648;
#10;x=-452583648;
#10;x=-452483648;
#10;x=-452383648;
#10;x=-452283648;
#10;x=-452183648;
#10;x=-452083648;
#10;x=-451983648;
#10;x=-451883648;
#10;x=-451783648;
#10;x=-451683648;
#10;x=-451583648;
#10;x=-451483648;
#10;x=-451383648;
#10;x=-451283648;
#10;x=-451183648;
#10;x=-451083648;
#10;x=-450983648;
#10;x=-450883648;
#10;x=-450783648;
#10;x=-450683648;
#10;x=-450583648;
#10;x=-450483648;
#10;x=-450383648;
#10;x=-450283648;
#10;x=-450183648;
#10;x=-450083648;
#10;x=-449983648;
#10;x=-449883648;
#10;x=-449783648;
#10;x=-449683648;
#10;x=-449583648;
#10;x=-449483648;
#10;x=-449383648;
#10;x=-449283648;
#10;x=-449183648;
#10;x=-449083648;
#10;x=-448983648;
#10;x=-448883648;
#10;x=-448783648;
#10;x=-448683648;
#10;x=-448583648;
#10;x=-448483648;
#10;x=-448383648;
#10;x=-448283648;
#10;x=-448183648;
#10;x=-448083648;
#10;x=-447983648;
#10;x=-447883648;
#10;x=-447783648;
#10;x=-447683648;
#10;x=-447583648;
#10;x=-447483648;
#10;x=-447383648;
#10;x=-447283648;
#10;x=-447183648;
#10;x=-447083648;
#10;x=-446983648;
#10;x=-446883648;
#10;x=-446783648;
#10;x=-446683648;
#10;x=-446583648;
#10;x=-446483648;
#10;x=-446383648;
#10;x=-446283648;
#10;x=-446183648;
#10;x=-446083648;
#10;x=-445983648;
#10;x=-445883648;
#10;x=-445783648;
#10;x=-445683648;
#10;x=-445583648;
#10;x=-445483648;
#10;x=-445383648;
#10;x=-445283648;
#10;x=-445183648;
#10;x=-445083648;
#10;x=-444983648;
#10;x=-444883648;
#10;x=-444783648;
#10;x=-444683648;
#10;x=-444583648;
#10;x=-444483648;
#10;x=-444383648;
#10;x=-444283648;
#10;x=-444183648;
#10;x=-444083648;
#10;x=-443983648;
#10;x=-443883648;
#10;x=-443783648;
#10;x=-443683648;
#10;x=-443583648;
#10;x=-443483648;
#10;x=-443383648;
#10;x=-443283648;
#10;x=-443183648;
#10;x=-443083648;
#10;x=-442983648;
#10;x=-442883648;
#10;x=-442783648;
#10;x=-442683648;
#10;x=-442583648;
#10;x=-442483648;
#10;x=-442383648;
#10;x=-442283648;
#10;x=-442183648;
#10;x=-442083648;
#10;x=-441983648;
#10;x=-441883648;
#10;x=-441783648;
#10;x=-441683648;
#10;x=-441583648;
#10;x=-441483648;
#10;x=-441383648;
#10;x=-441283648;
#10;x=-441183648;
#10;x=-441083648;
#10;x=-440983648;
#10;x=-440883648;
#10;x=-440783648;
#10;x=-440683648;
#10;x=-440583648;
#10;x=-440483648;
#10;x=-440383648;
#10;x=-440283648;
#10;x=-440183648;
#10;x=-440083648;
#10;x=-439983648;
#10;x=-439883648;
#10;x=-439783648;
#10;x=-439683648;
#10;x=-439583648;
#10;x=-439483648;
#10;x=-439383648;
#10;x=-439283648;
#10;x=-439183648;
#10;x=-439083648;
#10;x=-438983648;
#10;x=-438883648;
#10;x=-438783648;
#10;x=-438683648;
#10;x=-438583648;
#10;x=-438483648;
#10;x=-438383648;
#10;x=-438283648;
#10;x=-438183648;
#10;x=-438083648;
#10;x=-437983648;
#10;x=-437883648;
#10;x=-437783648;
#10;x=-437683648;
#10;x=-437583648;
#10;x=-437483648;
#10;x=-437383648;
#10;x=-437283648;
#10;x=-437183648;
#10;x=-437083648;
#10;x=-436983648;
#10;x=-436883648;
#10;x=-436783648;
#10;x=-436683648;
#10;x=-436583648;
#10;x=-436483648;
#10;x=-436383648;
#10;x=-436283648;
#10;x=-436183648;
#10;x=-436083648;
#10;x=-435983648;
#10;x=-435883648;
#10;x=-435783648;
#10;x=-435683648;
#10;x=-435583648;
#10;x=-435483648;
#10;x=-435383648;
#10;x=-435283648;
#10;x=-435183648;
#10;x=-435083648;
#10;x=-434983648;
#10;x=-434883648;
#10;x=-434783648;
#10;x=-434683648;
#10;x=-434583648;
#10;x=-434483648;
#10;x=-434383648;
#10;x=-434283648;
#10;x=-434183648;
#10;x=-434083648;
#10;x=-433983648;
#10;x=-433883648;
#10;x=-433783648;
#10;x=-433683648;
#10;x=-433583648;
#10;x=-433483648;
#10;x=-433383648;
#10;x=-433283648;
#10;x=-433183648;
#10;x=-433083648;
#10;x=-432983648;
#10;x=-432883648;
#10;x=-432783648;
#10;x=-432683648;
#10;x=-432583648;
#10;x=-432483648;
#10;x=-432383648;
#10;x=-432283648;
#10;x=-432183648;
#10;x=-432083648;
#10;x=-431983648;
#10;x=-431883648;
#10;x=-431783648;
#10;x=-431683648;
#10;x=-431583648;
#10;x=-431483648;
#10;x=-431383648;
#10;x=-431283648;
#10;x=-431183648;
#10;x=-431083648;
#10;x=-430983648;
#10;x=-430883648;
#10;x=-430783648;
#10;x=-430683648;
#10;x=-430583648;
#10;x=-430483648;
#10;x=-430383648;
#10;x=-430283648;
#10;x=-430183648;
#10;x=-430083648;
#10;x=-429983648;
#10;x=-429883648;
#10;x=-429783648;
#10;x=-429683648;
#10;x=-429583648;
#10;x=-429483648;
#10;x=-429383648;
#10;x=-429283648;
#10;x=-429183648;
#10;x=-429083648;
#10;x=-428983648;
#10;x=-428883648;
#10;x=-428783648;
#10;x=-428683648;
#10;x=-428583648;
#10;x=-428483648;
#10;x=-428383648;
#10;x=-428283648;
#10;x=-428183648;
#10;x=-428083648;
#10;x=-427983648;
#10;x=-427883648;
#10;x=-427783648;
#10;x=-427683648;
#10;x=-427583648;
#10;x=-427483648;
#10;x=-427383648;
#10;x=-427283648;
#10;x=-427183648;
#10;x=-427083648;
#10;x=-426983648;
#10;x=-426883648;
#10;x=-426783648;
#10;x=-426683648;
#10;x=-426583648;
#10;x=-426483648;
#10;x=-426383648;
#10;x=-426283648;
#10;x=-426183648;
#10;x=-426083648;
#10;x=-425983648;
#10;x=-425883648;
#10;x=-425783648;
#10;x=-425683648;
#10;x=-425583648;
#10;x=-425483648;
#10;x=-425383648;
#10;x=-425283648;
#10;x=-425183648;
#10;x=-425083648;
#10;x=-424983648;
#10;x=-424883648;
#10;x=-424783648;
#10;x=-424683648;
#10;x=-424583648;
#10;x=-424483648;
#10;x=-424383648;
#10;x=-424283648;
#10;x=-424183648;
#10;x=-424083648;
#10;x=-423983648;
#10;x=-423883648;
#10;x=-423783648;
#10;x=-423683648;
#10;x=-423583648;
#10;x=-423483648;
#10;x=-423383648;
#10;x=-423283648;
#10;x=-423183648;
#10;x=-423083648;
#10;x=-422983648;
#10;x=-422883648;
#10;x=-422783648;
#10;x=-422683648;
#10;x=-422583648;
#10;x=-422483648;
#10;x=-422383648;
#10;x=-422283648;
#10;x=-422183648;
#10;x=-422083648;
#10;x=-421983648;
#10;x=-421883648;
#10;x=-421783648;
#10;x=-421683648;
#10;x=-421583648;
#10;x=-421483648;
#10;x=-421383648;
#10;x=-421283648;
#10;x=-421183648;
#10;x=-421083648;
#10;x=-420983648;
#10;x=-420883648;
#10;x=-420783648;
#10;x=-420683648;
#10;x=-420583648;
#10;x=-420483648;
#10;x=-420383648;
#10;x=-420283648;
#10;x=-420183648;
#10;x=-420083648;
#10;x=-419983648;
#10;x=-419883648;
#10;x=-419783648;
#10;x=-419683648;
#10;x=-419583648;
#10;x=-419483648;
#10;x=-419383648;
#10;x=-419283648;
#10;x=-419183648;
#10;x=-419083648;
#10;x=-418983648;
#10;x=-418883648;
#10;x=-418783648;
#10;x=-418683648;
#10;x=-418583648;
#10;x=-418483648;
#10;x=-418383648;
#10;x=-418283648;
#10;x=-418183648;
#10;x=-418083648;
#10;x=-417983648;
#10;x=-417883648;
#10;x=-417783648;
#10;x=-417683648;
#10;x=-417583648;
#10;x=-417483648;
#10;x=-417383648;
#10;x=-417283648;
#10;x=-417183648;
#10;x=-417083648;
#10;x=-416983648;
#10;x=-416883648;
#10;x=-416783648;
#10;x=-416683648;
#10;x=-416583648;
#10;x=-416483648;
#10;x=-416383648;
#10;x=-416283648;
#10;x=-416183648;
#10;x=-416083648;
#10;x=-415983648;
#10;x=-415883648;
#10;x=-415783648;
#10;x=-415683648;
#10;x=-415583648;
#10;x=-415483648;
#10;x=-415383648;
#10;x=-415283648;
#10;x=-415183648;
#10;x=-415083648;
#10;x=-414983648;
#10;x=-414883648;
#10;x=-414783648;
#10;x=-414683648;
#10;x=-414583648;
#10;x=-414483648;
#10;x=-414383648;
#10;x=-414283648;
#10;x=-414183648;
#10;x=-414083648;
#10;x=-413983648;
#10;x=-413883648;
#10;x=-413783648;
#10;x=-413683648;
#10;x=-413583648;
#10;x=-413483648;
#10;x=-413383648;
#10;x=-413283648;
#10;x=-413183648;
#10;x=-413083648;
#10;x=-412983648;
#10;x=-412883648;
#10;x=-412783648;
#10;x=-412683648;
#10;x=-412583648;
#10;x=-412483648;
#10;x=-412383648;
#10;x=-412283648;
#10;x=-412183648;
#10;x=-412083648;
#10;x=-411983648;
#10;x=-411883648;
#10;x=-411783648;
#10;x=-411683648;
#10;x=-411583648;
#10;x=-411483648;
#10;x=-411383648;
#10;x=-411283648;
#10;x=-411183648;
#10;x=-411083648;
#10;x=-410983648;
#10;x=-410883648;
#10;x=-410783648;
#10;x=-410683648;
#10;x=-410583648;
#10;x=-410483648;
#10;x=-410383648;
#10;x=-410283648;
#10;x=-410183648;
#10;x=-410083648;
#10;x=-409983648;
#10;x=-409883648;
#10;x=-409783648;
#10;x=-409683648;
#10;x=-409583648;
#10;x=-409483648;
#10;x=-409383648;
#10;x=-409283648;
#10;x=-409183648;
#10;x=-409083648;
#10;x=-408983648;
#10;x=-408883648;
#10;x=-408783648;
#10;x=-408683648;
#10;x=-408583648;
#10;x=-408483648;
#10;x=-408383648;
#10;x=-408283648;
#10;x=-408183648;
#10;x=-408083648;
#10;x=-407983648;
#10;x=-407883648;
#10;x=-407783648;
#10;x=-407683648;
#10;x=-407583648;
#10;x=-407483648;
#10;x=-407383648;
#10;x=-407283648;
#10;x=-407183648;
#10;x=-407083648;
#10;x=-406983648;
#10;x=-406883648;
#10;x=-406783648;
#10;x=-406683648;
#10;x=-406583648;
#10;x=-406483648;
#10;x=-406383648;
#10;x=-406283648;
#10;x=-406183648;
#10;x=-406083648;
#10;x=-405983648;
#10;x=-405883648;
#10;x=-405783648;
#10;x=-405683648;
#10;x=-405583648;
#10;x=-405483648;
#10;x=-405383648;
#10;x=-405283648;
#10;x=-405183648;
#10;x=-405083648;
#10;x=-404983648;
#10;x=-404883648;
#10;x=-404783648;
#10;x=-404683648;
#10;x=-404583648;
#10;x=-404483648;
#10;x=-404383648;
#10;x=-404283648;
#10;x=-404183648;
#10;x=-404083648;
#10;x=-403983648;
#10;x=-403883648;
#10;x=-403783648;
#10;x=-403683648;
#10;x=-403583648;
#10;x=-403483648;
#10;x=-403383648;
#10;x=-403283648;
#10;x=-403183648;
#10;x=-403083648;
#10;x=-402983648;
#10;x=-402883648;
#10;x=-402783648;
#10;x=-402683648;
#10;x=-402583648;
#10;x=-402483648;
#10;x=-402383648;
#10;x=-402283648;
#10;x=-402183648;
#10;x=-402083648;
#10;x=-401983648;
#10;x=-401883648;
#10;x=-401783648;
#10;x=-401683648;
#10;x=-401583648;
#10;x=-401483648;
#10;x=-401383648;
#10;x=-401283648;
#10;x=-401183648;
#10;x=-401083648;
#10;x=-400983648;
#10;x=-400883648;
#10;x=-400783648;
#10;x=-400683648;
#10;x=-400583648;
#10;x=-400483648;
#10;x=-400383648;
#10;x=-400283648;
#10;x=-400183648;
#10;x=-400083648;
#10;x=-399983648;
#10;x=-399883648;
#10;x=-399783648;
#10;x=-399683648;
#10;x=-399583648;
#10;x=-399483648;
#10;x=-399383648;
#10;x=-399283648;
#10;x=-399183648;
#10;x=-399083648;
#10;x=-398983648;
#10;x=-398883648;
#10;x=-398783648;
#10;x=-398683648;
#10;x=-398583648;
#10;x=-398483648;
#10;x=-398383648;
#10;x=-398283648;
#10;x=-398183648;
#10;x=-398083648;
#10;x=-397983648;
#10;x=-397883648;
#10;x=-397783648;
#10;x=-397683648;
#10;x=-397583648;
#10;x=-397483648;
#10;x=-397383648;
#10;x=-397283648;
#10;x=-397183648;
#10;x=-397083648;
#10;x=-396983648;
#10;x=-396883648;
#10;x=-396783648;
#10;x=-396683648;
#10;x=-396583648;
#10;x=-396483648;
#10;x=-396383648;
#10;x=-396283648;
#10;x=-396183648;
#10;x=-396083648;
#10;x=-395983648;
#10;x=-395883648;
#10;x=-395783648;
#10;x=-395683648;
#10;x=-395583648;
#10;x=-395483648;
#10;x=-395383648;
#10;x=-395283648;
#10;x=-395183648;
#10;x=-395083648;
#10;x=-394983648;
#10;x=-394883648;
#10;x=-394783648;
#10;x=-394683648;
#10;x=-394583648;
#10;x=-394483648;
#10;x=-394383648;
#10;x=-394283648;
#10;x=-394183648;
#10;x=-394083648;
#10;x=-393983648;
#10;x=-393883648;
#10;x=-393783648;
#10;x=-393683648;
#10;x=-393583648;
#10;x=-393483648;
#10;x=-393383648;
#10;x=-393283648;
#10;x=-393183648;
#10;x=-393083648;
#10;x=-392983648;
#10;x=-392883648;
#10;x=-392783648;
#10;x=-392683648;
#10;x=-392583648;
#10;x=-392483648;
#10;x=-392383648;
#10;x=-392283648;
#10;x=-392183648;
#10;x=-392083648;
#10;x=-391983648;
#10;x=-391883648;
#10;x=-391783648;
#10;x=-391683648;
#10;x=-391583648;
#10;x=-391483648;
#10;x=-391383648;
#10;x=-391283648;
#10;x=-391183648;
#10;x=-391083648;
#10;x=-390983648;
#10;x=-390883648;
#10;x=-390783648;
#10;x=-390683648;
#10;x=-390583648;
#10;x=-390483648;
#10;x=-390383648;
#10;x=-390283648;
#10;x=-390183648;
#10;x=-390083648;
#10;x=-389983648;
#10;x=-389883648;
#10;x=-389783648;
#10;x=-389683648;
#10;x=-389583648;
#10;x=-389483648;
#10;x=-389383648;
#10;x=-389283648;
#10;x=-389183648;
#10;x=-389083648;
#10;x=-388983648;
#10;x=-388883648;
#10;x=-388783648;
#10;x=-388683648;
#10;x=-388583648;
#10;x=-388483648;
#10;x=-388383648;
#10;x=-388283648;
#10;x=-388183648;
#10;x=-388083648;
#10;x=-387983648;
#10;x=-387883648;
#10;x=-387783648;
#10;x=-387683648;
#10;x=-387583648;
#10;x=-387483648;
#10;x=-387383648;
#10;x=-387283648;
#10;x=-387183648;
#10;x=-387083648;
#10;x=-386983648;
#10;x=-386883648;
#10;x=-386783648;
#10;x=-386683648;
#10;x=-386583648;
#10;x=-386483648;
#10;x=-386383648;
#10;x=-386283648;
#10;x=-386183648;
#10;x=-386083648;
#10;x=-385983648;
#10;x=-385883648;
#10;x=-385783648;
#10;x=-385683648;
#10;x=-385583648;
#10;x=-385483648;
#10;x=-385383648;
#10;x=-385283648;
#10;x=-385183648;
#10;x=-385083648;
#10;x=-384983648;
#10;x=-384883648;
#10;x=-384783648;
#10;x=-384683648;
#10;x=-384583648;
#10;x=-384483648;
#10;x=-384383648;
#10;x=-384283648;
#10;x=-384183648;
#10;x=-384083648;
#10;x=-383983648;
#10;x=-383883648;
#10;x=-383783648;
#10;x=-383683648;
#10;x=-383583648;
#10;x=-383483648;
#10;x=-383383648;
#10;x=-383283648;
#10;x=-383183648;
#10;x=-383083648;
#10;x=-382983648;
#10;x=-382883648;
#10;x=-382783648;
#10;x=-382683648;
#10;x=-382583648;
#10;x=-382483648;
#10;x=-382383648;
#10;x=-382283648;
#10;x=-382183648;
#10;x=-382083648;
#10;x=-381983648;
#10;x=-381883648;
#10;x=-381783648;
#10;x=-381683648;
#10;x=-381583648;
#10;x=-381483648;
#10;x=-381383648;
#10;x=-381283648;
#10;x=-381183648;
#10;x=-381083648;
#10;x=-380983648;
#10;x=-380883648;
#10;x=-380783648;
#10;x=-380683648;
#10;x=-380583648;
#10;x=-380483648;
#10;x=-380383648;
#10;x=-380283648;
#10;x=-380183648;
#10;x=-380083648;
#10;x=-379983648;
#10;x=-379883648;
#10;x=-379783648;
#10;x=-379683648;
#10;x=-379583648;
#10;x=-379483648;
#10;x=-379383648;
#10;x=-379283648;
#10;x=-379183648;
#10;x=-379083648;
#10;x=-378983648;
#10;x=-378883648;
#10;x=-378783648;
#10;x=-378683648;
#10;x=-378583648;
#10;x=-378483648;
#10;x=-378383648;
#10;x=-378283648;
#10;x=-378183648;
#10;x=-378083648;
#10;x=-377983648;
#10;x=-377883648;
#10;x=-377783648;
#10;x=-377683648;
#10;x=-377583648;
#10;x=-377483648;
#10;x=-377383648;
#10;x=-377283648;
#10;x=-377183648;
#10;x=-377083648;
#10;x=-376983648;
#10;x=-376883648;
#10;x=-376783648;
#10;x=-376683648;
#10;x=-376583648;
#10;x=-376483648;
#10;x=-376383648;
#10;x=-376283648;
#10;x=-376183648;
#10;x=-376083648;
#10;x=-375983648;
#10;x=-375883648;
#10;x=-375783648;
#10;x=-375683648;
#10;x=-375583648;
#10;x=-375483648;
#10;x=-375383648;
#10;x=-375283648;
#10;x=-375183648;
#10;x=-375083648;
#10;x=-374983648;
#10;x=-374883648;
#10;x=-374783648;
#10;x=-374683648;
#10;x=-374583648;
#10;x=-374483648;
#10;x=-374383648;
#10;x=-374283648;
#10;x=-374183648;
#10;x=-374083648;
#10;x=-373983648;
#10;x=-373883648;
#10;x=-373783648;
#10;x=-373683648;
#10;x=-373583648;
#10;x=-373483648;
#10;x=-373383648;
#10;x=-373283648;
#10;x=-373183648;
#10;x=-373083648;
#10;x=-372983648;
#10;x=-372883648;
#10;x=-372783648;
#10;x=-372683648;
#10;x=-372583648;
#10;x=-372483648;
#10;x=-372383648;
#10;x=-372283648;
#10;x=-372183648;
#10;x=-372083648;
#10;x=-371983648;
#10;x=-371883648;
#10;x=-371783648;
#10;x=-371683648;
#10;x=-371583648;
#10;x=-371483648;
#10;x=-371383648;
#10;x=-371283648;
#10;x=-371183648;
#10;x=-371083648;
#10;x=-370983648;
#10;x=-370883648;
#10;x=-370783648;
#10;x=-370683648;
#10;x=-370583648;
#10;x=-370483648;
#10;x=-370383648;
#10;x=-370283648;
#10;x=-370183648;
#10;x=-370083648;
#10;x=-369983648;
#10;x=-369883648;
#10;x=-369783648;
#10;x=-369683648;
#10;x=-369583648;
#10;x=-369483648;
#10;x=-369383648;
#10;x=-369283648;
#10;x=-369183648;
#10;x=-369083648;
#10;x=-368983648;
#10;x=-368883648;
#10;x=-368783648;
#10;x=-368683648;
#10;x=-368583648;
#10;x=-368483648;
#10;x=-368383648;
#10;x=-368283648;
#10;x=-368183648;
#10;x=-368083648;
#10;x=-367983648;
#10;x=-367883648;
#10;x=-367783648;
#10;x=-367683648;
#10;x=-367583648;
#10;x=-367483648;
#10;x=-367383648;
#10;x=-367283648;
#10;x=-367183648;
#10;x=-367083648;
#10;x=-366983648;
#10;x=-366883648;
#10;x=-366783648;
#10;x=-366683648;
#10;x=-366583648;
#10;x=-366483648;
#10;x=-366383648;
#10;x=-366283648;
#10;x=-366183648;
#10;x=-366083648;
#10;x=-365983648;
#10;x=-365883648;
#10;x=-365783648;
#10;x=-365683648;
#10;x=-365583648;
#10;x=-365483648;
#10;x=-365383648;
#10;x=-365283648;
#10;x=-365183648;
#10;x=-365083648;
#10;x=-364983648;
#10;x=-364883648;
#10;x=-364783648;
#10;x=-364683648;
#10;x=-364583648;
#10;x=-364483648;
#10;x=-364383648;
#10;x=-364283648;
#10;x=-364183648;
#10;x=-364083648;
#10;x=-363983648;
#10;x=-363883648;
#10;x=-363783648;
#10;x=-363683648;
#10;x=-363583648;
#10;x=-363483648;
#10;x=-363383648;
#10;x=-363283648;
#10;x=-363183648;
#10;x=-363083648;
#10;x=-362983648;
#10;x=-362883648;
#10;x=-362783648;
#10;x=-362683648;
#10;x=-362583648;
#10;x=-362483648;
#10;x=-362383648;
#10;x=-362283648;
#10;x=-362183648;
#10;x=-362083648;
#10;x=-361983648;
#10;x=-361883648;
#10;x=-361783648;
#10;x=-361683648;
#10;x=-361583648;
#10;x=-361483648;
#10;x=-361383648;
#10;x=-361283648;
#10;x=-361183648;
#10;x=-361083648;
#10;x=-360983648;
#10;x=-360883648;
#10;x=-360783648;
#10;x=-360683648;
#10;x=-360583648;
#10;x=-360483648;
#10;x=-360383648;
#10;x=-360283648;
#10;x=-360183648;
#10;x=-360083648;
#10;x=-359983648;
#10;x=-359883648;
#10;x=-359783648;
#10;x=-359683648;
#10;x=-359583648;
#10;x=-359483648;
#10;x=-359383648;
#10;x=-359283648;
#10;x=-359183648;
#10;x=-359083648;
#10;x=-358983648;
#10;x=-358883648;
#10;x=-358783648;
#10;x=-358683648;
#10;x=-358583648;
#10;x=-358483648;
#10;x=-358383648;
#10;x=-358283648;
#10;x=-358183648;
#10;x=-358083648;
#10;x=-357983648;
#10;x=-357883648;
#10;x=-357783648;
#10;x=-357683648;
#10;x=-357583648;
#10;x=-357483648;
#10;x=-357383648;
#10;x=-357283648;
#10;x=-357183648;
#10;x=-357083648;
#10;x=-356983648;
#10;x=-356883648;
#10;x=-356783648;
#10;x=-356683648;
#10;x=-356583648;
#10;x=-356483648;
#10;x=-356383648;
#10;x=-356283648;
#10;x=-356183648;
#10;x=-356083648;
#10;x=-355983648;
#10;x=-355883648;
#10;x=-355783648;
#10;x=-355683648;
#10;x=-355583648;
#10;x=-355483648;
#10;x=-355383648;
#10;x=-355283648;
#10;x=-355183648;
#10;x=-355083648;
#10;x=-354983648;
#10;x=-354883648;
#10;x=-354783648;
#10;x=-354683648;
#10;x=-354583648;
#10;x=-354483648;
#10;x=-354383648;
#10;x=-354283648;
#10;x=-354183648;
#10;x=-354083648;
#10;x=-353983648;
#10;x=-353883648;
#10;x=-353783648;
#10;x=-353683648;
#10;x=-353583648;
#10;x=-353483648;
#10;x=-353383648;
#10;x=-353283648;
#10;x=-353183648;
#10;x=-353083648;
#10;x=-352983648;
#10;x=-352883648;
#10;x=-352783648;
#10;x=-352683648;
#10;x=-352583648;
#10;x=-352483648;
#10;x=-352383648;
#10;x=-352283648;
#10;x=-352183648;
#10;x=-352083648;
#10;x=-351983648;
#10;x=-351883648;
#10;x=-351783648;
#10;x=-351683648;
#10;x=-351583648;
#10;x=-351483648;
#10;x=-351383648;
#10;x=-351283648;
#10;x=-351183648;
#10;x=-351083648;
#10;x=-350983648;
#10;x=-350883648;
#10;x=-350783648;
#10;x=-350683648;
#10;x=-350583648;
#10;x=-350483648;
#10;x=-350383648;
#10;x=-350283648;
#10;x=-350183648;
#10;x=-350083648;
#10;x=-349983648;
#10;x=-349883648;
#10;x=-349783648;
#10;x=-349683648;
#10;x=-349583648;
#10;x=-349483648;
#10;x=-349383648;
#10;x=-349283648;
#10;x=-349183648;
#10;x=-349083648;
#10;x=-348983648;
#10;x=-348883648;
#10;x=-348783648;
#10;x=-348683648;
#10;x=-348583648;
#10;x=-348483648;
#10;x=-348383648;
#10;x=-348283648;
#10;x=-348183648;
#10;x=-348083648;
#10;x=-347983648;
#10;x=-347883648;
#10;x=-347783648;
#10;x=-347683648;
#10;x=-347583648;
#10;x=-347483648;
#10;x=-347383648;
#10;x=-347283648;
#10;x=-347183648;
#10;x=-347083648;
#10;x=-346983648;
#10;x=-346883648;
#10;x=-346783648;
#10;x=-346683648;
#10;x=-346583648;
#10;x=-346483648;
#10;x=-346383648;
#10;x=-346283648;
#10;x=-346183648;
#10;x=-346083648;
#10;x=-345983648;
#10;x=-345883648;
#10;x=-345783648;
#10;x=-345683648;
#10;x=-345583648;
#10;x=-345483648;
#10;x=-345383648;
#10;x=-345283648;
#10;x=-345183648;
#10;x=-345083648;
#10;x=-344983648;
#10;x=-344883648;
#10;x=-344783648;
#10;x=-344683648;
#10;x=-344583648;
#10;x=-344483648;
#10;x=-344383648;
#10;x=-344283648;
#10;x=-344183648;
#10;x=-344083648;
#10;x=-343983648;
#10;x=-343883648;
#10;x=-343783648;
#10;x=-343683648;
#10;x=-343583648;
#10;x=-343483648;
#10;x=-343383648;
#10;x=-343283648;
#10;x=-343183648;
#10;x=-343083648;
#10;x=-342983648;
#10;x=-342883648;
#10;x=-342783648;
#10;x=-342683648;
#10;x=-342583648;
#10;x=-342483648;
#10;x=-342383648;
#10;x=-342283648;
#10;x=-342183648;
#10;x=-342083648;
#10;x=-341983648;
#10;x=-341883648;
#10;x=-341783648;
#10;x=-341683648;
#10;x=-341583648;
#10;x=-341483648;
#10;x=-341383648;
#10;x=-341283648;
#10;x=-341183648;
#10;x=-341083648;
#10;x=-340983648;
#10;x=-340883648;
#10;x=-340783648;
#10;x=-340683648;
#10;x=-340583648;
#10;x=-340483648;
#10;x=-340383648;
#10;x=-340283648;
#10;x=-340183648;
#10;x=-340083648;
#10;x=-339983648;
#10;x=-339883648;
#10;x=-339783648;
#10;x=-339683648;
#10;x=-339583648;
#10;x=-339483648;
#10;x=-339383648;
#10;x=-339283648;
#10;x=-339183648;
#10;x=-339083648;
#10;x=-338983648;
#10;x=-338883648;
#10;x=-338783648;
#10;x=-338683648;
#10;x=-338583648;
#10;x=-338483648;
#10;x=-338383648;
#10;x=-338283648;
#10;x=-338183648;
#10;x=-338083648;
#10;x=-337983648;
#10;x=-337883648;
#10;x=-337783648;
#10;x=-337683648;
#10;x=-337583648;
#10;x=-337483648;
#10;x=-337383648;
#10;x=-337283648;
#10;x=-337183648;
#10;x=-337083648;
#10;x=-336983648;
#10;x=-336883648;
#10;x=-336783648;
#10;x=-336683648;
#10;x=-336583648;
#10;x=-336483648;
#10;x=-336383648;
#10;x=-336283648;
#10;x=-336183648;
#10;x=-336083648;
#10;x=-335983648;
#10;x=-335883648;
#10;x=-335783648;
#10;x=-335683648;
#10;x=-335583648;
#10;x=-335483648;
#10;x=-335383648;
#10;x=-335283648;
#10;x=-335183648;
#10;x=-335083648;
#10;x=-334983648;
#10;x=-334883648;
#10;x=-334783648;
#10;x=-334683648;
#10;x=-334583648;
#10;x=-334483648;
#10;x=-334383648;
#10;x=-334283648;
#10;x=-334183648;
#10;x=-334083648;
#10;x=-333983648;
#10;x=-333883648;
#10;x=-333783648;
#10;x=-333683648;
#10;x=-333583648;
#10;x=-333483648;
#10;x=-333383648;
#10;x=-333283648;
#10;x=-333183648;
#10;x=-333083648;
#10;x=-332983648;
#10;x=-332883648;
#10;x=-332783648;
#10;x=-332683648;
#10;x=-332583648;
#10;x=-332483648;
#10;x=-332383648;
#10;x=-332283648;
#10;x=-332183648;
#10;x=-332083648;
#10;x=-331983648;
#10;x=-331883648;
#10;x=-331783648;
#10;x=-331683648;
#10;x=-331583648;
#10;x=-331483648;
#10;x=-331383648;
#10;x=-331283648;
#10;x=-331183648;
#10;x=-331083648;
#10;x=-330983648;
#10;x=-330883648;
#10;x=-330783648;
#10;x=-330683648;
#10;x=-330583648;
#10;x=-330483648;
#10;x=-330383648;
#10;x=-330283648;
#10;x=-330183648;
#10;x=-330083648;
#10;x=-329983648;
#10;x=-329883648;
#10;x=-329783648;
#10;x=-329683648;
#10;x=-329583648;
#10;x=-329483648;
#10;x=-329383648;
#10;x=-329283648;
#10;x=-329183648;
#10;x=-329083648;
#10;x=-328983648;
#10;x=-328883648;
#10;x=-328783648;
#10;x=-328683648;
#10;x=-328583648;
#10;x=-328483648;
#10;x=-328383648;
#10;x=-328283648;
#10;x=-328183648;
#10;x=-328083648;
#10;x=-327983648;
#10;x=-327883648;
#10;x=-327783648;
#10;x=-327683648;
#10;x=-327583648;
#10;x=-327483648;
#10;x=-327383648;
#10;x=-327283648;
#10;x=-327183648;
#10;x=-327083648;
#10;x=-326983648;
#10;x=-326883648;
#10;x=-326783648;
#10;x=-326683648;
#10;x=-326583648;
#10;x=-326483648;
#10;x=-326383648;
#10;x=-326283648;
#10;x=-326183648;
#10;x=-326083648;
#10;x=-325983648;
#10;x=-325883648;
#10;x=-325783648;
#10;x=-325683648;
#10;x=-325583648;
#10;x=-325483648;
#10;x=-325383648;
#10;x=-325283648;
#10;x=-325183648;
#10;x=-325083648;
#10;x=-324983648;
#10;x=-324883648;
#10;x=-324783648;
#10;x=-324683648;
#10;x=-324583648;
#10;x=-324483648;
#10;x=-324383648;
#10;x=-324283648;
#10;x=-324183648;
#10;x=-324083648;
#10;x=-323983648;
#10;x=-323883648;
#10;x=-323783648;
#10;x=-323683648;
#10;x=-323583648;
#10;x=-323483648;
#10;x=-323383648;
#10;x=-323283648;
#10;x=-323183648;
#10;x=-323083648;
#10;x=-322983648;
#10;x=-322883648;
#10;x=-322783648;
#10;x=-322683648;
#10;x=-322583648;
#10;x=-322483648;
#10;x=-322383648;
#10;x=-322283648;
#10;x=-322183648;
#10;x=-322083648;
#10;x=-321983648;
#10;x=-321883648;
#10;x=-321783648;
#10;x=-321683648;
#10;x=-321583648;
#10;x=-321483648;
#10;x=-321383648;
#10;x=-321283648;
#10;x=-321183648;
#10;x=-321083648;
#10;x=-320983648;
#10;x=-320883648;
#10;x=-320783648;
#10;x=-320683648;
#10;x=-320583648;
#10;x=-320483648;
#10;x=-320383648;
#10;x=-320283648;
#10;x=-320183648;
#10;x=-320083648;
#10;x=-319983648;
#10;x=-319883648;
#10;x=-319783648;
#10;x=-319683648;
#10;x=-319583648;
#10;x=-319483648;
#10;x=-319383648;
#10;x=-319283648;
#10;x=-319183648;
#10;x=-319083648;
#10;x=-318983648;
#10;x=-318883648;
#10;x=-318783648;
#10;x=-318683648;
#10;x=-318583648;
#10;x=-318483648;
#10;x=-318383648;
#10;x=-318283648;
#10;x=-318183648;
#10;x=-318083648;
#10;x=-317983648;
#10;x=-317883648;
#10;x=-317783648;
#10;x=-317683648;
#10;x=-317583648;
#10;x=-317483648;
#10;x=-317383648;
#10;x=-317283648;
#10;x=-317183648;
#10;x=-317083648;
#10;x=-316983648;
#10;x=-316883648;
#10;x=-316783648;
#10;x=-316683648;
#10;x=-316583648;
#10;x=-316483648;
#10;x=-316383648;
#10;x=-316283648;
#10;x=-316183648;
#10;x=-316083648;
#10;x=-315983648;
#10;x=-315883648;
#10;x=-315783648;
#10;x=-315683648;
#10;x=-315583648;
#10;x=-315483648;
#10;x=-315383648;
#10;x=-315283648;
#10;x=-315183648;
#10;x=-315083648;
#10;x=-314983648;
#10;x=-314883648;
#10;x=-314783648;
#10;x=-314683648;
#10;x=-314583648;
#10;x=-314483648;
#10;x=-314383648;
#10;x=-314283648;
#10;x=-314183648;
#10;x=-314083648;
#10;x=-313983648;
#10;x=-313883648;
#10;x=-313783648;
#10;x=-313683648;
#10;x=-313583648;
#10;x=-313483648;
#10;x=-313383648;
#10;x=-313283648;
#10;x=-313183648;
#10;x=-313083648;
#10;x=-312983648;
#10;x=-312883648;
#10;x=-312783648;
#10;x=-312683648;
#10;x=-312583648;
#10;x=-312483648;
#10;x=-312383648;
#10;x=-312283648;
#10;x=-312183648;
#10;x=-312083648;
#10;x=-311983648;
#10;x=-311883648;
#10;x=-311783648;
#10;x=-311683648;
#10;x=-311583648;
#10;x=-311483648;
#10;x=-311383648;
#10;x=-311283648;
#10;x=-311183648;
#10;x=-311083648;
#10;x=-310983648;
#10;x=-310883648;
#10;x=-310783648;
#10;x=-310683648;
#10;x=-310583648;
#10;x=-310483648;
#10;x=-310383648;
#10;x=-310283648;
#10;x=-310183648;
#10;x=-310083648;
#10;x=-309983648;
#10;x=-309883648;
#10;x=-309783648;
#10;x=-309683648;
#10;x=-309583648;
#10;x=-309483648;
#10;x=-309383648;
#10;x=-309283648;
#10;x=-309183648;
#10;x=-309083648;
#10;x=-308983648;
#10;x=-308883648;
#10;x=-308783648;
#10;x=-308683648;
#10;x=-308583648;
#10;x=-308483648;
#10;x=-308383648;
#10;x=-308283648;
#10;x=-308183648;
#10;x=-308083648;
#10;x=-307983648;
#10;x=-307883648;
#10;x=-307783648;
#10;x=-307683648;
#10;x=-307583648;
#10;x=-307483648;
#10;x=-307383648;
#10;x=-307283648;
#10;x=-307183648;
#10;x=-307083648;
#10;x=-306983648;
#10;x=-306883648;
#10;x=-306783648;
#10;x=-306683648;
#10;x=-306583648;
#10;x=-306483648;
#10;x=-306383648;
#10;x=-306283648;
#10;x=-306183648;
#10;x=-306083648;
#10;x=-305983648;
#10;x=-305883648;
#10;x=-305783648;
#10;x=-305683648;
#10;x=-305583648;
#10;x=-305483648;
#10;x=-305383648;
#10;x=-305283648;
#10;x=-305183648;
#10;x=-305083648;
#10;x=-304983648;
#10;x=-304883648;
#10;x=-304783648;
#10;x=-304683648;
#10;x=-304583648;
#10;x=-304483648;
#10;x=-304383648;
#10;x=-304283648;
#10;x=-304183648;
#10;x=-304083648;
#10;x=-303983648;
#10;x=-303883648;
#10;x=-303783648;
#10;x=-303683648;
#10;x=-303583648;
#10;x=-303483648;
#10;x=-303383648;
#10;x=-303283648;
#10;x=-303183648;
#10;x=-303083648;
#10;x=-302983648;
#10;x=-302883648;
#10;x=-302783648;
#10;x=-302683648;
#10;x=-302583648;
#10;x=-302483648;
#10;x=-302383648;
#10;x=-302283648;
#10;x=-302183648;
#10;x=-302083648;
#10;x=-301983648;
#10;x=-301883648;
#10;x=-301783648;
#10;x=-301683648;
#10;x=-301583648;
#10;x=-301483648;
#10;x=-301383648;
#10;x=-301283648;
#10;x=-301183648;
#10;x=-301083648;
#10;x=-300983648;
#10;x=-300883648;
#10;x=-300783648;
#10;x=-300683648;
#10;x=-300583648;
#10;x=-300483648;
#10;x=-300383648;
#10;x=-300283648;
#10;x=-300183648;
#10;x=-300083648;
#10;x=-299983648;
#10;x=-299883648;
#10;x=-299783648;
#10;x=-299683648;
#10;x=-299583648;
#10;x=-299483648;
#10;x=-299383648;
#10;x=-299283648;
#10;x=-299183648;
#10;x=-299083648;
#10;x=-298983648;
#10;x=-298883648;
#10;x=-298783648;
#10;x=-298683648;
#10;x=-298583648;
#10;x=-298483648;
#10;x=-298383648;
#10;x=-298283648;
#10;x=-298183648;
#10;x=-298083648;
#10;x=-297983648;
#10;x=-297883648;
#10;x=-297783648;
#10;x=-297683648;
#10;x=-297583648;
#10;x=-297483648;
#10;x=-297383648;
#10;x=-297283648;
#10;x=-297183648;
#10;x=-297083648;
#10;x=-296983648;
#10;x=-296883648;
#10;x=-296783648;
#10;x=-296683648;
#10;x=-296583648;
#10;x=-296483648;
#10;x=-296383648;
#10;x=-296283648;
#10;x=-296183648;
#10;x=-296083648;
#10;x=-295983648;
#10;x=-295883648;
#10;x=-295783648;
#10;x=-295683648;
#10;x=-295583648;
#10;x=-295483648;
#10;x=-295383648;
#10;x=-295283648;
#10;x=-295183648;
#10;x=-295083648;
#10;x=-294983648;
#10;x=-294883648;
#10;x=-294783648;
#10;x=-294683648;
#10;x=-294583648;
#10;x=-294483648;
#10;x=-294383648;
#10;x=-294283648;
#10;x=-294183648;
#10;x=-294083648;
#10;x=-293983648;
#10;x=-293883648;
#10;x=-293783648;
#10;x=-293683648;
#10;x=-293583648;
#10;x=-293483648;
#10;x=-293383648;
#10;x=-293283648;
#10;x=-293183648;
#10;x=-293083648;
#10;x=-292983648;
#10;x=-292883648;
#10;x=-292783648;
#10;x=-292683648;
#10;x=-292583648;
#10;x=-292483648;
#10;x=-292383648;
#10;x=-292283648;
#10;x=-292183648;
#10;x=-292083648;
#10;x=-291983648;
#10;x=-291883648;
#10;x=-291783648;
#10;x=-291683648;
#10;x=-291583648;
#10;x=-291483648;
#10;x=-291383648;
#10;x=-291283648;
#10;x=-291183648;
#10;x=-291083648;
#10;x=-290983648;
#10;x=-290883648;
#10;x=-290783648;
#10;x=-290683648;
#10;x=-290583648;
#10;x=-290483648;
#10;x=-290383648;
#10;x=-290283648;
#10;x=-290183648;
#10;x=-290083648;
#10;x=-289983648;
#10;x=-289883648;
#10;x=-289783648;
#10;x=-289683648;
#10;x=-289583648;
#10;x=-289483648;
#10;x=-289383648;
#10;x=-289283648;
#10;x=-289183648;
#10;x=-289083648;
#10;x=-288983648;
#10;x=-288883648;
#10;x=-288783648;
#10;x=-288683648;
#10;x=-288583648;
#10;x=-288483648;
#10;x=-288383648;
#10;x=-288283648;
#10;x=-288183648;
#10;x=-288083648;
#10;x=-287983648;
#10;x=-287883648;
#10;x=-287783648;
#10;x=-287683648;
#10;x=-287583648;
#10;x=-287483648;
#10;x=-287383648;
#10;x=-287283648;
#10;x=-287183648;
#10;x=-287083648;
#10;x=-286983648;
#10;x=-286883648;
#10;x=-286783648;
#10;x=-286683648;
#10;x=-286583648;
#10;x=-286483648;
#10;x=-286383648;
#10;x=-286283648;
#10;x=-286183648;
#10;x=-286083648;
#10;x=-285983648;
#10;x=-285883648;
#10;x=-285783648;
#10;x=-285683648;
#10;x=-285583648;
#10;x=-285483648;
#10;x=-285383648;
#10;x=-285283648;
#10;x=-285183648;
#10;x=-285083648;
#10;x=-284983648;
#10;x=-284883648;
#10;x=-284783648;
#10;x=-284683648;
#10;x=-284583648;
#10;x=-284483648;
#10;x=-284383648;
#10;x=-284283648;
#10;x=-284183648;
#10;x=-284083648;
#10;x=-283983648;
#10;x=-283883648;
#10;x=-283783648;
#10;x=-283683648;
#10;x=-283583648;
#10;x=-283483648;
#10;x=-283383648;
#10;x=-283283648;
#10;x=-283183648;
#10;x=-283083648;
#10;x=-282983648;
#10;x=-282883648;
#10;x=-282783648;
#10;x=-282683648;
#10;x=-282583648;
#10;x=-282483648;
#10;x=-282383648;
#10;x=-282283648;
#10;x=-282183648;
#10;x=-282083648;
#10;x=-281983648;
#10;x=-281883648;
#10;x=-281783648;
#10;x=-281683648;
#10;x=-281583648;
#10;x=-281483648;
#10;x=-281383648;
#10;x=-281283648;
#10;x=-281183648;
#10;x=-281083648;
#10;x=-280983648;
#10;x=-280883648;
#10;x=-280783648;
#10;x=-280683648;
#10;x=-280583648;
#10;x=-280483648;
#10;x=-280383648;
#10;x=-280283648;
#10;x=-280183648;
#10;x=-280083648;
#10;x=-279983648;
#10;x=-279883648;
#10;x=-279783648;
#10;x=-279683648;
#10;x=-279583648;
#10;x=-279483648;
#10;x=-279383648;
#10;x=-279283648;
#10;x=-279183648;
#10;x=-279083648;
#10;x=-278983648;
#10;x=-278883648;
#10;x=-278783648;
#10;x=-278683648;
#10;x=-278583648;
#10;x=-278483648;
#10;x=-278383648;
#10;x=-278283648;
#10;x=-278183648;
#10;x=-278083648;
#10;x=-277983648;
#10;x=-277883648;
#10;x=-277783648;
#10;x=-277683648;
#10;x=-277583648;
#10;x=-277483648;
#10;x=-277383648;
#10;x=-277283648;
#10;x=-277183648;
#10;x=-277083648;
#10;x=-276983648;
#10;x=-276883648;
#10;x=-276783648;
#10;x=-276683648;
#10;x=-276583648;
#10;x=-276483648;
#10;x=-276383648;
#10;x=-276283648;
#10;x=-276183648;
#10;x=-276083648;
#10;x=-275983648;
#10;x=-275883648;
#10;x=-275783648;
#10;x=-275683648;
#10;x=-275583648;
#10;x=-275483648;
#10;x=-275383648;
#10;x=-275283648;
#10;x=-275183648;
#10;x=-275083648;
#10;x=-274983648;
#10;x=-274883648;
#10;x=-274783648;
#10;x=-274683648;
#10;x=-274583648;
#10;x=-274483648;
#10;x=-274383648;
#10;x=-274283648;
#10;x=-274183648;
#10;x=-274083648;
#10;x=-273983648;
#10;x=-273883648;
#10;x=-273783648;
#10;x=-273683648;
#10;x=-273583648;
#10;x=-273483648;
#10;x=-273383648;
#10;x=-273283648;
#10;x=-273183648;
#10;x=-273083648;
#10;x=-272983648;
#10;x=-272883648;
#10;x=-272783648;
#10;x=-272683648;
#10;x=-272583648;
#10;x=-272483648;
#10;x=-272383648;
#10;x=-272283648;
#10;x=-272183648;
#10;x=-272083648;
#10;x=-271983648;
#10;x=-271883648;
#10;x=-271783648;
#10;x=-271683648;
#10;x=-271583648;
#10;x=-271483648;
#10;x=-271383648;
#10;x=-271283648;
#10;x=-271183648;
#10;x=-271083648;
#10;x=-270983648;
#10;x=-270883648;
#10;x=-270783648;
#10;x=-270683648;
#10;x=-270583648;
#10;x=-270483648;
#10;x=-270383648;
#10;x=-270283648;
#10;x=-270183648;
#10;x=-270083648;
#10;x=-269983648;
#10;x=-269883648;
#10;x=-269783648;
#10;x=-269683648;
#10;x=-269583648;
#10;x=-269483648;
#10;x=-269383648;
#10;x=-269283648;
#10;x=-269183648;
#10;x=-269083648;
#10;x=-268983648;
#10;x=-268883648;
#10;x=-268783648;
#10;x=-268683648;
#10;x=-268583648;
#10;x=-268483648;
#10;x=-268383648;
#10;x=-268283648;
#10;x=-268183648;
#10;x=-268083648;
#10;x=-267983648;
#10;x=-267883648;
#10;x=-267783648;
#10;x=-267683648;
#10;x=-267583648;
#10;x=-267483648;
#10;x=-267383648;
#10;x=-267283648;
#10;x=-267183648;
#10;x=-267083648;
#10;x=-266983648;
#10;x=-266883648;
#10;x=-266783648;
#10;x=-266683648;
#10;x=-266583648;
#10;x=-266483648;
#10;x=-266383648;
#10;x=-266283648;
#10;x=-266183648;
#10;x=-266083648;
#10;x=-265983648;
#10;x=-265883648;
#10;x=-265783648;
#10;x=-265683648;
#10;x=-265583648;
#10;x=-265483648;
#10;x=-265383648;
#10;x=-265283648;
#10;x=-265183648;
#10;x=-265083648;
#10;x=-264983648;
#10;x=-264883648;
#10;x=-264783648;
#10;x=-264683648;
#10;x=-264583648;
#10;x=-264483648;
#10;x=-264383648;
#10;x=-264283648;
#10;x=-264183648;
#10;x=-264083648;
#10;x=-263983648;
#10;x=-263883648;
#10;x=-263783648;
#10;x=-263683648;
#10;x=-263583648;
#10;x=-263483648;
#10;x=-263383648;
#10;x=-263283648;
#10;x=-263183648;
#10;x=-263083648;
#10;x=-262983648;
#10;x=-262883648;
#10;x=-262783648;
#10;x=-262683648;
#10;x=-262583648;
#10;x=-262483648;
#10;x=-262383648;
#10;x=-262283648;
#10;x=-262183648;
#10;x=-262083648;
#10;x=-261983648;
#10;x=-261883648;
#10;x=-261783648;
#10;x=-261683648;
#10;x=-261583648;
#10;x=-261483648;
#10;x=-261383648;
#10;x=-261283648;
#10;x=-261183648;
#10;x=-261083648;
#10;x=-260983648;
#10;x=-260883648;
#10;x=-260783648;
#10;x=-260683648;
#10;x=-260583648;
#10;x=-260483648;
#10;x=-260383648;
#10;x=-260283648;
#10;x=-260183648;
#10;x=-260083648;
#10;x=-259983648;
#10;x=-259883648;
#10;x=-259783648;
#10;x=-259683648;
#10;x=-259583648;
#10;x=-259483648;
#10;x=-259383648;
#10;x=-259283648;
#10;x=-259183648;
#10;x=-259083648;
#10;x=-258983648;
#10;x=-258883648;
#10;x=-258783648;
#10;x=-258683648;
#10;x=-258583648;
#10;x=-258483648;
#10;x=-258383648;
#10;x=-258283648;
#10;x=-258183648;
#10;x=-258083648;
#10;x=-257983648;
#10;x=-257883648;
#10;x=-257783648;
#10;x=-257683648;
#10;x=-257583648;
#10;x=-257483648;
#10;x=-257383648;
#10;x=-257283648;
#10;x=-257183648;
#10;x=-257083648;
#10;x=-256983648;
#10;x=-256883648;
#10;x=-256783648;
#10;x=-256683648;
#10;x=-256583648;
#10;x=-256483648;
#10;x=-256383648;
#10;x=-256283648;
#10;x=-256183648;
#10;x=-256083648;
#10;x=-255983648;
#10;x=-255883648;
#10;x=-255783648;
#10;x=-255683648;
#10;x=-255583648;
#10;x=-255483648;
#10;x=-255383648;
#10;x=-255283648;
#10;x=-255183648;
#10;x=-255083648;
#10;x=-254983648;
#10;x=-254883648;
#10;x=-254783648;
#10;x=-254683648;
#10;x=-254583648;
#10;x=-254483648;
#10;x=-254383648;
#10;x=-254283648;
#10;x=-254183648;
#10;x=-254083648;
#10;x=-253983648;
#10;x=-253883648;
#10;x=-253783648;
#10;x=-253683648;
#10;x=-253583648;
#10;x=-253483648;
#10;x=-253383648;
#10;x=-253283648;
#10;x=-253183648;
#10;x=-253083648;
#10;x=-252983648;
#10;x=-252883648;
#10;x=-252783648;
#10;x=-252683648;
#10;x=-252583648;
#10;x=-252483648;
#10;x=-252383648;
#10;x=-252283648;
#10;x=-252183648;
#10;x=-252083648;
#10;x=-251983648;
#10;x=-251883648;
#10;x=-251783648;
#10;x=-251683648;
#10;x=-251583648;
#10;x=-251483648;
#10;x=-251383648;
#10;x=-251283648;
#10;x=-251183648;
#10;x=-251083648;
#10;x=-250983648;
#10;x=-250883648;
#10;x=-250783648;
#10;x=-250683648;
#10;x=-250583648;
#10;x=-250483648;
#10;x=-250383648;
#10;x=-250283648;
#10;x=-250183648;
#10;x=-250083648;
#10;x=-249983648;
#10;x=-249883648;
#10;x=-249783648;
#10;x=-249683648;
#10;x=-249583648;
#10;x=-249483648;
#10;x=-249383648;
#10;x=-249283648;
#10;x=-249183648;
#10;x=-249083648;
#10;x=-248983648;
#10;x=-248883648;
#10;x=-248783648;
#10;x=-248683648;
#10;x=-248583648;
#10;x=-248483648;
#10;x=-248383648;
#10;x=-248283648;
#10;x=-248183648;
#10;x=-248083648;
#10;x=-247983648;
#10;x=-247883648;
#10;x=-247783648;
#10;x=-247683648;
#10;x=-247583648;
#10;x=-247483648;
#10;x=-247383648;
#10;x=-247283648;
#10;x=-247183648;
#10;x=-247083648;
#10;x=-246983648;
#10;x=-246883648;
#10;x=-246783648;
#10;x=-246683648;
#10;x=-246583648;
#10;x=-246483648;
#10;x=-246383648;
#10;x=-246283648;
#10;x=-246183648;
#10;x=-246083648;
#10;x=-245983648;
#10;x=-245883648;
#10;x=-245783648;
#10;x=-245683648;
#10;x=-245583648;
#10;x=-245483648;
#10;x=-245383648;
#10;x=-245283648;
#10;x=-245183648;
#10;x=-245083648;
#10;x=-244983648;
#10;x=-244883648;
#10;x=-244783648;
#10;x=-244683648;
#10;x=-244583648;
#10;x=-244483648;
#10;x=-244383648;
#10;x=-244283648;
#10;x=-244183648;
#10;x=-244083648;
#10;x=-243983648;
#10;x=-243883648;
#10;x=-243783648;
#10;x=-243683648;
#10;x=-243583648;
#10;x=-243483648;
#10;x=-243383648;
#10;x=-243283648;
#10;x=-243183648;
#10;x=-243083648;
#10;x=-242983648;
#10;x=-242883648;
#10;x=-242783648;
#10;x=-242683648;
#10;x=-242583648;
#10;x=-242483648;
#10;x=-242383648;
#10;x=-242283648;
#10;x=-242183648;
#10;x=-242083648;
#10;x=-241983648;
#10;x=-241883648;
#10;x=-241783648;
#10;x=-241683648;
#10;x=-241583648;
#10;x=-241483648;
#10;x=-241383648;
#10;x=-241283648;
#10;x=-241183648;
#10;x=-241083648;
#10;x=-240983648;
#10;x=-240883648;
#10;x=-240783648;
#10;x=-240683648;
#10;x=-240583648;
#10;x=-240483648;
#10;x=-240383648;
#10;x=-240283648;
#10;x=-240183648;
#10;x=-240083648;
#10;x=-239983648;
#10;x=-239883648;
#10;x=-239783648;
#10;x=-239683648;
#10;x=-239583648;
#10;x=-239483648;
#10;x=-239383648;
#10;x=-239283648;
#10;x=-239183648;
#10;x=-239083648;
#10;x=-238983648;
#10;x=-238883648;
#10;x=-238783648;
#10;x=-238683648;
#10;x=-238583648;
#10;x=-238483648;
#10;x=-238383648;
#10;x=-238283648;
#10;x=-238183648;
#10;x=-238083648;
#10;x=-237983648;
#10;x=-237883648;
#10;x=-237783648;
#10;x=-237683648;
#10;x=-237583648;
#10;x=-237483648;
#10;x=-237383648;
#10;x=-237283648;
#10;x=-237183648;
#10;x=-237083648;
#10;x=-236983648;
#10;x=-236883648;
#10;x=-236783648;
#10;x=-236683648;
#10;x=-236583648;
#10;x=-236483648;
#10;x=-236383648;
#10;x=-236283648;
#10;x=-236183648;
#10;x=-236083648;
#10;x=-235983648;
#10;x=-235883648;
#10;x=-235783648;
#10;x=-235683648;
#10;x=-235583648;
#10;x=-235483648;
#10;x=-235383648;
#10;x=-235283648;
#10;x=-235183648;
#10;x=-235083648;
#10;x=-234983648;
#10;x=-234883648;
#10;x=-234783648;
#10;x=-234683648;
#10;x=-234583648;
#10;x=-234483648;
#10;x=-234383648;
#10;x=-234283648;
#10;x=-234183648;
#10;x=-234083648;
#10;x=-233983648;
#10;x=-233883648;
#10;x=-233783648;
#10;x=-233683648;
#10;x=-233583648;
#10;x=-233483648;
#10;x=-233383648;
#10;x=-233283648;
#10;x=-233183648;
#10;x=-233083648;
#10;x=-232983648;
#10;x=-232883648;
#10;x=-232783648;
#10;x=-232683648;
#10;x=-232583648;
#10;x=-232483648;
#10;x=-232383648;
#10;x=-232283648;
#10;x=-232183648;
#10;x=-232083648;
#10;x=-231983648;
#10;x=-231883648;
#10;x=-231783648;
#10;x=-231683648;
#10;x=-231583648;
#10;x=-231483648;
#10;x=-231383648;
#10;x=-231283648;
#10;x=-231183648;
#10;x=-231083648;
#10;x=-230983648;
#10;x=-230883648;
#10;x=-230783648;
#10;x=-230683648;
#10;x=-230583648;
#10;x=-230483648;
#10;x=-230383648;
#10;x=-230283648;
#10;x=-230183648;
#10;x=-230083648;
#10;x=-229983648;
#10;x=-229883648;
#10;x=-229783648;
#10;x=-229683648;
#10;x=-229583648;
#10;x=-229483648;
#10;x=-229383648;
#10;x=-229283648;
#10;x=-229183648;
#10;x=-229083648;
#10;x=-228983648;
#10;x=-228883648;
#10;x=-228783648;
#10;x=-228683648;
#10;x=-228583648;
#10;x=-228483648;
#10;x=-228383648;
#10;x=-228283648;
#10;x=-228183648;
#10;x=-228083648;
#10;x=-227983648;
#10;x=-227883648;
#10;x=-227783648;
#10;x=-227683648;
#10;x=-227583648;
#10;x=-227483648;
#10;x=-227383648;
#10;x=-227283648;
#10;x=-227183648;
#10;x=-227083648;
#10;x=-226983648;
#10;x=-226883648;
#10;x=-226783648;
#10;x=-226683648;
#10;x=-226583648;
#10;x=-226483648;
#10;x=-226383648;
#10;x=-226283648;
#10;x=-226183648;
#10;x=-226083648;
#10;x=-225983648;
#10;x=-225883648;
#10;x=-225783648;
#10;x=-225683648;
#10;x=-225583648;
#10;x=-225483648;
#10;x=-225383648;
#10;x=-225283648;
#10;x=-225183648;
#10;x=-225083648;
#10;x=-224983648;
#10;x=-224883648;
#10;x=-224783648;
#10;x=-224683648;
#10;x=-224583648;
#10;x=-224483648;
#10;x=-224383648;
#10;x=-224283648;
#10;x=-224183648;
#10;x=-224083648;
#10;x=-223983648;
#10;x=-223883648;
#10;x=-223783648;
#10;x=-223683648;
#10;x=-223583648;
#10;x=-223483648;
#10;x=-223383648;
#10;x=-223283648;
#10;x=-223183648;
#10;x=-223083648;
#10;x=-222983648;
#10;x=-222883648;
#10;x=-222783648;
#10;x=-222683648;
#10;x=-222583648;
#10;x=-222483648;
#10;x=-222383648;
#10;x=-222283648;
#10;x=-222183648;
#10;x=-222083648;
#10;x=-221983648;
#10;x=-221883648;
#10;x=-221783648;
#10;x=-221683648;
#10;x=-221583648;
#10;x=-221483648;
#10;x=-221383648;
#10;x=-221283648;
#10;x=-221183648;
#10;x=-221083648;
#10;x=-220983648;
#10;x=-220883648;
#10;x=-220783648;
#10;x=-220683648;
#10;x=-220583648;
#10;x=-220483648;
#10;x=-220383648;
#10;x=-220283648;
#10;x=-220183648;
#10;x=-220083648;
#10;x=-219983648;
#10;x=-219883648;
#10;x=-219783648;
#10;x=-219683648;
#10;x=-219583648;
#10;x=-219483648;
#10;x=-219383648;
#10;x=-219283648;
#10;x=-219183648;
#10;x=-219083648;
#10;x=-218983648;
#10;x=-218883648;
#10;x=-218783648;
#10;x=-218683648;
#10;x=-218583648;
#10;x=-218483648;
#10;x=-218383648;
#10;x=-218283648;
#10;x=-218183648;
#10;x=-218083648;
#10;x=-217983648;
#10;x=-217883648;
#10;x=-217783648;
#10;x=-217683648;
#10;x=-217583648;
#10;x=-217483648;
#10;x=-217383648;
#10;x=-217283648;
#10;x=-217183648;
#10;x=-217083648;
#10;x=-216983648;
#10;x=-216883648;
#10;x=-216783648;
#10;x=-216683648;
#10;x=-216583648;
#10;x=-216483648;
#10;x=-216383648;
#10;x=-216283648;
#10;x=-216183648;
#10;x=-216083648;
#10;x=-215983648;
#10;x=-215883648;
#10;x=-215783648;
#10;x=-215683648;
#10;x=-215583648;
#10;x=-215483648;
#10;x=-215383648;
#10;x=-215283648;
#10;x=-215183648;
#10;x=-215083648;
#10;x=-214983648;
#10;x=-214883648;
#10;x=-214783648;
#10;x=-214683648;
#10;x=-214583648;
#10;x=-214483648;
#10;x=-214383648;
#10;x=-214283648;
#10;x=-214183648;
#10;x=-214083648;
#10;x=-213983648;
#10;x=-213883648;
#10;x=-213783648;
#10;x=-213683648;
#10;x=-213583648;
#10;x=-213483648;
#10;x=-213383648;
#10;x=-213283648;
#10;x=-213183648;
#10;x=-213083648;
#10;x=-212983648;
#10;x=-212883648;
#10;x=-212783648;
#10;x=-212683648;
#10;x=-212583648;
#10;x=-212483648;
#10;x=-212383648;
#10;x=-212283648;
#10;x=-212183648;
#10;x=-212083648;
#10;x=-211983648;
#10;x=-211883648;
#10;x=-211783648;
#10;x=-211683648;
#10;x=-211583648;
#10;x=-211483648;
#10;x=-211383648;
#10;x=-211283648;
#10;x=-211183648;
#10;x=-211083648;
#10;x=-210983648;
#10;x=-210883648;
#10;x=-210783648;
#10;x=-210683648;
#10;x=-210583648;
#10;x=-210483648;
#10;x=-210383648;
#10;x=-210283648;
#10;x=-210183648;
#10;x=-210083648;
#10;x=-209983648;
#10;x=-209883648;
#10;x=-209783648;
#10;x=-209683648;
#10;x=-209583648;
#10;x=-209483648;
#10;x=-209383648;
#10;x=-209283648;
#10;x=-209183648;
#10;x=-209083648;
#10;x=-208983648;
#10;x=-208883648;
#10;x=-208783648;
#10;x=-208683648;
#10;x=-208583648;
#10;x=-208483648;
#10;x=-208383648;
#10;x=-208283648;
#10;x=-208183648;
#10;x=-208083648;
#10;x=-207983648;
#10;x=-207883648;
#10;x=-207783648;
#10;x=-207683648;
#10;x=-207583648;
#10;x=-207483648;
#10;x=-207383648;
#10;x=-207283648;
#10;x=-207183648;
#10;x=-207083648;
#10;x=-206983648;
#10;x=-206883648;
#10;x=-206783648;
#10;x=-206683648;
#10;x=-206583648;
#10;x=-206483648;
#10;x=-206383648;
#10;x=-206283648;
#10;x=-206183648;
#10;x=-206083648;
#10;x=-205983648;
#10;x=-205883648;
#10;x=-205783648;
#10;x=-205683648;
#10;x=-205583648;
#10;x=-205483648;
#10;x=-205383648;
#10;x=-205283648;
#10;x=-205183648;
#10;x=-205083648;
#10;x=-204983648;
#10;x=-204883648;
#10;x=-204783648;
#10;x=-204683648;
#10;x=-204583648;
#10;x=-204483648;
#10;x=-204383648;
#10;x=-204283648;
#10;x=-204183648;
#10;x=-204083648;
#10;x=-203983648;
#10;x=-203883648;
#10;x=-203783648;
#10;x=-203683648;
#10;x=-203583648;
#10;x=-203483648;
#10;x=-203383648;
#10;x=-203283648;
#10;x=-203183648;
#10;x=-203083648;
#10;x=-202983648;
#10;x=-202883648;
#10;x=-202783648;
#10;x=-202683648;
#10;x=-202583648;
#10;x=-202483648;
#10;x=-202383648;
#10;x=-202283648;
#10;x=-202183648;
#10;x=-202083648;
#10;x=-201983648;
#10;x=-201883648;
#10;x=-201783648;
#10;x=-201683648;
#10;x=-201583648;
#10;x=-201483648;
#10;x=-201383648;
#10;x=-201283648;
#10;x=-201183648;
#10;x=-201083648;
#10;x=-200983648;
#10;x=-200883648;
#10;x=-200783648;
#10;x=-200683648;
#10;x=-200583648;
#10;x=-200483648;
#10;x=-200383648;
#10;x=-200283648;
#10;x=-200183648;
#10;x=-200083648;
#10;x=-199983648;
#10;x=-199883648;
#10;x=-199783648;
#10;x=-199683648;
#10;x=-199583648;
#10;x=-199483648;
#10;x=-199383648;
#10;x=-199283648;
#10;x=-199183648;
#10;x=-199083648;
#10;x=-198983648;
#10;x=-198883648;
#10;x=-198783648;
#10;x=-198683648;
#10;x=-198583648;
#10;x=-198483648;
#10;x=-198383648;
#10;x=-198283648;
#10;x=-198183648;
#10;x=-198083648;
#10;x=-197983648;
#10;x=-197883648;
#10;x=-197783648;
#10;x=-197683648;
#10;x=-197583648;
#10;x=-197483648;
#10;x=-197383648;
#10;x=-197283648;
#10;x=-197183648;
#10;x=-197083648;
#10;x=-196983648;
#10;x=-196883648;
#10;x=-196783648;
#10;x=-196683648;
#10;x=-196583648;
#10;x=-196483648;
#10;x=-196383648;
#10;x=-196283648;
#10;x=-196183648;
#10;x=-196083648;
#10;x=-195983648;
#10;x=-195883648;
#10;x=-195783648;
#10;x=-195683648;
#10;x=-195583648;
#10;x=-195483648;
#10;x=-195383648;
#10;x=-195283648;
#10;x=-195183648;
#10;x=-195083648;
#10;x=-194983648;
#10;x=-194883648;
#10;x=-194783648;
#10;x=-194683648;
#10;x=-194583648;
#10;x=-194483648;
#10;x=-194383648;
#10;x=-194283648;
#10;x=-194183648;
#10;x=-194083648;
#10;x=-193983648;
#10;x=-193883648;
#10;x=-193783648;
#10;x=-193683648;
#10;x=-193583648;
#10;x=-193483648;
#10;x=-193383648;
#10;x=-193283648;
#10;x=-193183648;
#10;x=-193083648;
#10;x=-192983648;
#10;x=-192883648;
#10;x=-192783648;
#10;x=-192683648;
#10;x=-192583648;
#10;x=-192483648;
#10;x=-192383648;
#10;x=-192283648;
#10;x=-192183648;
#10;x=-192083648;
#10;x=-191983648;
#10;x=-191883648;
#10;x=-191783648;
#10;x=-191683648;
#10;x=-191583648;
#10;x=-191483648;
#10;x=-191383648;
#10;x=-191283648;
#10;x=-191183648;
#10;x=-191083648;
#10;x=-190983648;
#10;x=-190883648;
#10;x=-190783648;
#10;x=-190683648;
#10;x=-190583648;
#10;x=-190483648;
#10;x=-190383648;
#10;x=-190283648;
#10;x=-190183648;
#10;x=-190083648;
#10;x=-189983648;
#10;x=-189883648;
#10;x=-189783648;
#10;x=-189683648;
#10;x=-189583648;
#10;x=-189483648;
#10;x=-189383648;
#10;x=-189283648;
#10;x=-189183648;
#10;x=-189083648;
#10;x=-188983648;
#10;x=-188883648;
#10;x=-188783648;
#10;x=-188683648;
#10;x=-188583648;
#10;x=-188483648;
#10;x=-188383648;
#10;x=-188283648;
#10;x=-188183648;
#10;x=-188083648;
#10;x=-187983648;
#10;x=-187883648;
#10;x=-187783648;
#10;x=-187683648;
#10;x=-187583648;
#10;x=-187483648;
#10;x=-187383648;
#10;x=-187283648;
#10;x=-187183648;
#10;x=-187083648;
#10;x=-186983648;
#10;x=-186883648;
#10;x=-186783648;
#10;x=-186683648;
#10;x=-186583648;
#10;x=-186483648;
#10;x=-186383648;
#10;x=-186283648;
#10;x=-186183648;
#10;x=-186083648;
#10;x=-185983648;
#10;x=-185883648;
#10;x=-185783648;
#10;x=-185683648;
#10;x=-185583648;
#10;x=-185483648;
#10;x=-185383648;
#10;x=-185283648;
#10;x=-185183648;
#10;x=-185083648;
#10;x=-184983648;
#10;x=-184883648;
#10;x=-184783648;
#10;x=-184683648;
#10;x=-184583648;
#10;x=-184483648;
#10;x=-184383648;
#10;x=-184283648;
#10;x=-184183648;
#10;x=-184083648;
#10;x=-183983648;
#10;x=-183883648;
#10;x=-183783648;
#10;x=-183683648;
#10;x=-183583648;
#10;x=-183483648;
#10;x=-183383648;
#10;x=-183283648;
#10;x=-183183648;
#10;x=-183083648;
#10;x=-182983648;
#10;x=-182883648;
#10;x=-182783648;
#10;x=-182683648;
#10;x=-182583648;
#10;x=-182483648;
#10;x=-182383648;
#10;x=-182283648;
#10;x=-182183648;
#10;x=-182083648;
#10;x=-181983648;
#10;x=-181883648;
#10;x=-181783648;
#10;x=-181683648;
#10;x=-181583648;
#10;x=-181483648;
#10;x=-181383648;
#10;x=-181283648;
#10;x=-181183648;
#10;x=-181083648;
#10;x=-180983648;
#10;x=-180883648;
#10;x=-180783648;
#10;x=-180683648;
#10;x=-180583648;
#10;x=-180483648;
#10;x=-180383648;
#10;x=-180283648;
#10;x=-180183648;
#10;x=-180083648;
#10;x=-179983648;
#10;x=-179883648;
#10;x=-179783648;
#10;x=-179683648;
#10;x=-179583648;
#10;x=-179483648;
#10;x=-179383648;
#10;x=-179283648;
#10;x=-179183648;
#10;x=-179083648;
#10;x=-178983648;
#10;x=-178883648;
#10;x=-178783648;
#10;x=-178683648;
#10;x=-178583648;
#10;x=-178483648;
#10;x=-178383648;
#10;x=-178283648;
#10;x=-178183648;
#10;x=-178083648;
#10;x=-177983648;
#10;x=-177883648;
#10;x=-177783648;
#10;x=-177683648;
#10;x=-177583648;
#10;x=-177483648;
#10;x=-177383648;
#10;x=-177283648;
#10;x=-177183648;
#10;x=-177083648;
#10;x=-176983648;
#10;x=-176883648;
#10;x=-176783648;
#10;x=-176683648;
#10;x=-176583648;
#10;x=-176483648;
#10;x=-176383648;
#10;x=-176283648;
#10;x=-176183648;
#10;x=-176083648;
#10;x=-175983648;
#10;x=-175883648;
#10;x=-175783648;
#10;x=-175683648;
#10;x=-175583648;
#10;x=-175483648;
#10;x=-175383648;
#10;x=-175283648;
#10;x=-175183648;
#10;x=-175083648;
#10;x=-174983648;
#10;x=-174883648;
#10;x=-174783648;
#10;x=-174683648;
#10;x=-174583648;
#10;x=-174483648;
#10;x=-174383648;
#10;x=-174283648;
#10;x=-174183648;
#10;x=-174083648;
#10;x=-173983648;
#10;x=-173883648;
#10;x=-173783648;
#10;x=-173683648;
#10;x=-173583648;
#10;x=-173483648;
#10;x=-173383648;
#10;x=-173283648;
#10;x=-173183648;
#10;x=-173083648;
#10;x=-172983648;
#10;x=-172883648;
#10;x=-172783648;
#10;x=-172683648;
#10;x=-172583648;
#10;x=-172483648;
#10;x=-172383648;
#10;x=-172283648;
#10;x=-172183648;
#10;x=-172083648;
#10;x=-171983648;
#10;x=-171883648;
#10;x=-171783648;
#10;x=-171683648;
#10;x=-171583648;
#10;x=-171483648;
#10;x=-171383648;
#10;x=-171283648;
#10;x=-171183648;
#10;x=-171083648;
#10;x=-170983648;
#10;x=-170883648;
#10;x=-170783648;
#10;x=-170683648;
#10;x=-170583648;
#10;x=-170483648;
#10;x=-170383648;
#10;x=-170283648;
#10;x=-170183648;
#10;x=-170083648;
#10;x=-169983648;
#10;x=-169883648;
#10;x=-169783648;
#10;x=-169683648;
#10;x=-169583648;
#10;x=-169483648;
#10;x=-169383648;
#10;x=-169283648;
#10;x=-169183648;
#10;x=-169083648;
#10;x=-168983648;
#10;x=-168883648;
#10;x=-168783648;
#10;x=-168683648;
#10;x=-168583648;
#10;x=-168483648;
#10;x=-168383648;
#10;x=-168283648;
#10;x=-168183648;
#10;x=-168083648;
#10;x=-167983648;
#10;x=-167883648;
#10;x=-167783648;
#10;x=-167683648;
#10;x=-167583648;
#10;x=-167483648;
#10;x=-167383648;
#10;x=-167283648;
#10;x=-167183648;
#10;x=-167083648;
#10;x=-166983648;
#10;x=-166883648;
#10;x=-166783648;
#10;x=-166683648;
#10;x=-166583648;
#10;x=-166483648;
#10;x=-166383648;
#10;x=-166283648;
#10;x=-166183648;
#10;x=-166083648;
#10;x=-165983648;
#10;x=-165883648;
#10;x=-165783648;
#10;x=-165683648;
#10;x=-165583648;
#10;x=-165483648;
#10;x=-165383648;
#10;x=-165283648;
#10;x=-165183648;
#10;x=-165083648;
#10;x=-164983648;
#10;x=-164883648;
#10;x=-164783648;
#10;x=-164683648;
#10;x=-164583648;
#10;x=-164483648;
#10;x=-164383648;
#10;x=-164283648;
#10;x=-164183648;
#10;x=-164083648;
#10;x=-163983648;
#10;x=-163883648;
#10;x=-163783648;
#10;x=-163683648;
#10;x=-163583648;
#10;x=-163483648;
#10;x=-163383648;
#10;x=-163283648;
#10;x=-163183648;
#10;x=-163083648;
#10;x=-162983648;
#10;x=-162883648;
#10;x=-162783648;
#10;x=-162683648;
#10;x=-162583648;
#10;x=-162483648;
#10;x=-162383648;
#10;x=-162283648;
#10;x=-162183648;
#10;x=-162083648;
#10;x=-161983648;
#10;x=-161883648;
#10;x=-161783648;
#10;x=-161683648;
#10;x=-161583648;
#10;x=-161483648;
#10;x=-161383648;
#10;x=-161283648;
#10;x=-161183648;
#10;x=-161083648;
#10;x=-160983648;
#10;x=-160883648;
#10;x=-160783648;
#10;x=-160683648;
#10;x=-160583648;
#10;x=-160483648;
#10;x=-160383648;
#10;x=-160283648;
#10;x=-160183648;
#10;x=-160083648;
#10;x=-159983648;
#10;x=-159883648;
#10;x=-159783648;
#10;x=-159683648;
#10;x=-159583648;
#10;x=-159483648;
#10;x=-159383648;
#10;x=-159283648;
#10;x=-159183648;
#10;x=-159083648;
#10;x=-158983648;
#10;x=-158883648;
#10;x=-158783648;
#10;x=-158683648;
#10;x=-158583648;
#10;x=-158483648;
#10;x=-158383648;
#10;x=-158283648;
#10;x=-158183648;
#10;x=-158083648;
#10;x=-157983648;
#10;x=-157883648;
#10;x=-157783648;
#10;x=-157683648;
#10;x=-157583648;
#10;x=-157483648;
#10;x=-157383648;
#10;x=-157283648;
#10;x=-157183648;
#10;x=-157083648;
#10;x=-156983648;
#10;x=-156883648;
#10;x=-156783648;
#10;x=-156683648;
#10;x=-156583648;
#10;x=-156483648;
#10;x=-156383648;
#10;x=-156283648;
#10;x=-156183648;
#10;x=-156083648;
#10;x=-155983648;
#10;x=-155883648;
#10;x=-155783648;
#10;x=-155683648;
#10;x=-155583648;
#10;x=-155483648;
#10;x=-155383648;
#10;x=-155283648;
#10;x=-155183648;
#10;x=-155083648;
#10;x=-154983648;
#10;x=-154883648;
#10;x=-154783648;
#10;x=-154683648;
#10;x=-154583648;
#10;x=-154483648;
#10;x=-154383648;
#10;x=-154283648;
#10;x=-154183648;
#10;x=-154083648;
#10;x=-153983648;
#10;x=-153883648;
#10;x=-153783648;
#10;x=-153683648;
#10;x=-153583648;
#10;x=-153483648;
#10;x=-153383648;
#10;x=-153283648;
#10;x=-153183648;
#10;x=-153083648;
#10;x=-152983648;
#10;x=-152883648;
#10;x=-152783648;
#10;x=-152683648;
#10;x=-152583648;
#10;x=-152483648;
#10;x=-152383648;
#10;x=-152283648;
#10;x=-152183648;
#10;x=-152083648;
#10;x=-151983648;
#10;x=-151883648;
#10;x=-151783648;
#10;x=-151683648;
#10;x=-151583648;
#10;x=-151483648;
#10;x=-151383648;
#10;x=-151283648;
#10;x=-151183648;
#10;x=-151083648;
#10;x=-150983648;
#10;x=-150883648;
#10;x=-150783648;
#10;x=-150683648;
#10;x=-150583648;
#10;x=-150483648;
#10;x=-150383648;
#10;x=-150283648;
#10;x=-150183648;
#10;x=-150083648;
#10;x=-149983648;
#10;x=-149883648;
#10;x=-149783648;
#10;x=-149683648;
#10;x=-149583648;
#10;x=-149483648;
#10;x=-149383648;
#10;x=-149283648;
#10;x=-149183648;
#10;x=-149083648;
#10;x=-148983648;
#10;x=-148883648;
#10;x=-148783648;
#10;x=-148683648;
#10;x=-148583648;
#10;x=-148483648;
#10;x=-148383648;
#10;x=-148283648;
#10;x=-148183648;
#10;x=-148083648;
#10;x=-147983648;
#10;x=-147883648;
#10;x=-147783648;
#10;x=-147683648;
#10;x=-147583648;
#10;x=-147483648;
#10;x=-147383648;
#10;x=-147283648;
#10;x=-147183648;
#10;x=-147083648;
#10;x=-146983648;
#10;x=-146883648;
#10;x=-146783648;
#10;x=-146683648;
#10;x=-146583648;
#10;x=-146483648;
#10;x=-146383648;
#10;x=-146283648;
#10;x=-146183648;
#10;x=-146083648;
#10;x=-145983648;
#10;x=-145883648;
#10;x=-145783648;
#10;x=-145683648;
#10;x=-145583648;
#10;x=-145483648;
#10;x=-145383648;
#10;x=-145283648;
#10;x=-145183648;
#10;x=-145083648;
#10;x=-144983648;
#10;x=-144883648;
#10;x=-144783648;
#10;x=-144683648;
#10;x=-144583648;
#10;x=-144483648;
#10;x=-144383648;
#10;x=-144283648;
#10;x=-144183648;
#10;x=-144083648;
#10;x=-143983648;
#10;x=-143883648;
#10;x=-143783648;
#10;x=-143683648;
#10;x=-143583648;
#10;x=-143483648;
#10;x=-143383648;
#10;x=-143283648;
#10;x=-143183648;
#10;x=-143083648;
#10;x=-142983648;
#10;x=-142883648;
#10;x=-142783648;
#10;x=-142683648;
#10;x=-142583648;
#10;x=-142483648;
#10;x=-142383648;
#10;x=-142283648;
#10;x=-142183648;
#10;x=-142083648;
#10;x=-141983648;
#10;x=-141883648;
#10;x=-141783648;
#10;x=-141683648;
#10;x=-141583648;
#10;x=-141483648;
#10;x=-141383648;
#10;x=-141283648;
#10;x=-141183648;
#10;x=-141083648;
#10;x=-140983648;
#10;x=-140883648;
#10;x=-140783648;
#10;x=-140683648;
#10;x=-140583648;
#10;x=-140483648;
#10;x=-140383648;
#10;x=-140283648;
#10;x=-140183648;
#10;x=-140083648;
#10;x=-139983648;
#10;x=-139883648;
#10;x=-139783648;
#10;x=-139683648;
#10;x=-139583648;
#10;x=-139483648;
#10;x=-139383648;
#10;x=-139283648;
#10;x=-139183648;
#10;x=-139083648;
#10;x=-138983648;
#10;x=-138883648;
#10;x=-138783648;
#10;x=-138683648;
#10;x=-138583648;
#10;x=-138483648;
#10;x=-138383648;
#10;x=-138283648;
#10;x=-138183648;
#10;x=-138083648;
#10;x=-137983648;
#10;x=-137883648;
#10;x=-137783648;
#10;x=-137683648;
#10;x=-137583648;
#10;x=-137483648;
#10;x=-137383648;
#10;x=-137283648;
#10;x=-137183648;
#10;x=-137083648;
#10;x=-136983648;
#10;x=-136883648;
#10;x=-136783648;
#10;x=-136683648;
#10;x=-136583648;
#10;x=-136483648;
#10;x=-136383648;
#10;x=-136283648;
#10;x=-136183648;
#10;x=-136083648;
#10;x=-135983648;
#10;x=-135883648;
#10;x=-135783648;
#10;x=-135683648;
#10;x=-135583648;
#10;x=-135483648;
#10;x=-135383648;
#10;x=-135283648;
#10;x=-135183648;
#10;x=-135083648;
#10;x=-134983648;
#10;x=-134883648;
#10;x=-134783648;
#10;x=-134683648;
#10;x=-134583648;
#10;x=-134483648;
#10;x=-134383648;
#10;x=-134283648;
#10;x=-134183648;
#10;x=-134083648;
#10;x=-133983648;
#10;x=-133883648;
#10;x=-133783648;
#10;x=-133683648;
#10;x=-133583648;
#10;x=-133483648;
#10;x=-133383648;
#10;x=-133283648;
#10;x=-133183648;
#10;x=-133083648;
#10;x=-132983648;
#10;x=-132883648;
#10;x=-132783648;
#10;x=-132683648;
#10;x=-132583648;
#10;x=-132483648;
#10;x=-132383648;
#10;x=-132283648;
#10;x=-132183648;
#10;x=-132083648;
#10;x=-131983648;
#10;x=-131883648;
#10;x=-131783648;
#10;x=-131683648;
#10;x=-131583648;
#10;x=-131483648;
#10;x=-131383648;
#10;x=-131283648;
#10;x=-131183648;
#10;x=-131083648;
#10;x=-130983648;
#10;x=-130883648;
#10;x=-130783648;
#10;x=-130683648;
#10;x=-130583648;
#10;x=-130483648;
#10;x=-130383648;
#10;x=-130283648;
#10;x=-130183648;
#10;x=-130083648;
#10;x=-129983648;
#10;x=-129883648;
#10;x=-129783648;
#10;x=-129683648;
#10;x=-129583648;
#10;x=-129483648;
#10;x=-129383648;
#10;x=-129283648;
#10;x=-129183648;
#10;x=-129083648;
#10;x=-128983648;
#10;x=-128883648;
#10;x=-128783648;
#10;x=-128683648;
#10;x=-128583648;
#10;x=-128483648;
#10;x=-128383648;
#10;x=-128283648;
#10;x=-128183648;
#10;x=-128083648;
#10;x=-127983648;
#10;x=-127883648;
#10;x=-127783648;
#10;x=-127683648;
#10;x=-127583648;
#10;x=-127483648;
#10;x=-127383648;
#10;x=-127283648;
#10;x=-127183648;
#10;x=-127083648;
#10;x=-126983648;
#10;x=-126883648;
#10;x=-126783648;
#10;x=-126683648;
#10;x=-126583648;
#10;x=-126483648;
#10;x=-126383648;
#10;x=-126283648;
#10;x=-126183648;
#10;x=-126083648;
#10;x=-125983648;
#10;x=-125883648;
#10;x=-125783648;
#10;x=-125683648;
#10;x=-125583648;
#10;x=-125483648;
#10;x=-125383648;
#10;x=-125283648;
#10;x=-125183648;
#10;x=-125083648;
#10;x=-124983648;
#10;x=-124883648;
#10;x=-124783648;
#10;x=-124683648;
#10;x=-124583648;
#10;x=-124483648;
#10;x=-124383648;
#10;x=-124283648;
#10;x=-124183648;
#10;x=-124083648;
#10;x=-123983648;
#10;x=-123883648;
#10;x=-123783648;
#10;x=-123683648;
#10;x=-123583648;
#10;x=-123483648;
#10;x=-123383648;
#10;x=-123283648;
#10;x=-123183648;
#10;x=-123083648;
#10;x=-122983648;
#10;x=-122883648;
#10;x=-122783648;
#10;x=-122683648;
#10;x=-122583648;
#10;x=-122483648;
#10;x=-122383648;
#10;x=-122283648;
#10;x=-122183648;
#10;x=-122083648;
#10;x=-121983648;
#10;x=-121883648;
#10;x=-121783648;
#10;x=-121683648;
#10;x=-121583648;
#10;x=-121483648;
#10;x=-121383648;
#10;x=-121283648;
#10;x=-121183648;
#10;x=-121083648;
#10;x=-120983648;
#10;x=-120883648;
#10;x=-120783648;
#10;x=-120683648;
#10;x=-120583648;
#10;x=-120483648;
#10;x=-120383648;
#10;x=-120283648;
#10;x=-120183648;
#10;x=-120083648;
#10;x=-119983648;
#10;x=-119883648;
#10;x=-119783648;
#10;x=-119683648;
#10;x=-119583648;
#10;x=-119483648;
#10;x=-119383648;
#10;x=-119283648;
#10;x=-119183648;
#10;x=-119083648;
#10;x=-118983648;
#10;x=-118883648;
#10;x=-118783648;
#10;x=-118683648;
#10;x=-118583648;
#10;x=-118483648;
#10;x=-118383648;
#10;x=-118283648;
#10;x=-118183648;
#10;x=-118083648;
#10;x=-117983648;
#10;x=-117883648;
#10;x=-117783648;
#10;x=-117683648;
#10;x=-117583648;
#10;x=-117483648;
#10;x=-117383648;
#10;x=-117283648;
#10;x=-117183648;
#10;x=-117083648;
#10;x=-116983648;
#10;x=-116883648;
#10;x=-116783648;
#10;x=-116683648;
#10;x=-116583648;
#10;x=-116483648;
#10;x=-116383648;
#10;x=-116283648;
#10;x=-116183648;
#10;x=-116083648;
#10;x=-115983648;
#10;x=-115883648;
#10;x=-115783648;
#10;x=-115683648;
#10;x=-115583648;
#10;x=-115483648;
#10;x=-115383648;
#10;x=-115283648;
#10;x=-115183648;
#10;x=-115083648;
#10;x=-114983648;
#10;x=-114883648;
#10;x=-114783648;
#10;x=-114683648;
#10;x=-114583648;
#10;x=-114483648;
#10;x=-114383648;
#10;x=-114283648;
#10;x=-114183648;
#10;x=-114083648;
#10;x=-113983648;
#10;x=-113883648;
#10;x=-113783648;
#10;x=-113683648;
#10;x=-113583648;
#10;x=-113483648;
#10;x=-113383648;
#10;x=-113283648;
#10;x=-113183648;
#10;x=-113083648;
#10;x=-112983648;
#10;x=-112883648;
#10;x=-112783648;
#10;x=-112683648;
#10;x=-112583648;
#10;x=-112483648;
#10;x=-112383648;
#10;x=-112283648;
#10;x=-112183648;
#10;x=-112083648;
#10;x=-111983648;
#10;x=-111883648;
#10;x=-111783648;
#10;x=-111683648;
#10;x=-111583648;
#10;x=-111483648;
#10;x=-111383648;
#10;x=-111283648;
#10;x=-111183648;
#10;x=-111083648;
#10;x=-110983648;
#10;x=-110883648;
#10;x=-110783648;
#10;x=-110683648;
#10;x=-110583648;
#10;x=-110483648;
#10;x=-110383648;
#10;x=-110283648;
#10;x=-110183648;
#10;x=-110083648;
#10;x=-109983648;
#10;x=-109883648;
#10;x=-109783648;
#10;x=-109683648;
#10;x=-109583648;
#10;x=-109483648;
#10;x=-109383648;
#10;x=-109283648;
#10;x=-109183648;
#10;x=-109083648;
#10;x=-108983648;
#10;x=-108883648;
#10;x=-108783648;
#10;x=-108683648;
#10;x=-108583648;
#10;x=-108483648;
#10;x=-108383648;
#10;x=-108283648;
#10;x=-108183648;
#10;x=-108083648;
#10;x=-107983648;
#10;x=-107883648;
#10;x=-107783648;
#10;x=-107683648;
#10;x=-107583648;
#10;x=-107483648;
#10;x=-107383648;
#10;x=-107283648;
#10;x=-107183648;
#10;x=-107083648;
#10;x=-106983648;
#10;x=-106883648;
#10;x=-106783648;
#10;x=-106683648;
#10;x=-106583648;
#10;x=-106483648;
#10;x=-106383648;
#10;x=-106283648;
#10;x=-106183648;
#10;x=-106083648;
#10;x=-105983648;
#10;x=-105883648;
#10;x=-105783648;
#10;x=-105683648;
#10;x=-105583648;
#10;x=-105483648;
#10;x=-105383648;
#10;x=-105283648;
#10;x=-105183648;
#10;x=-105083648;
#10;x=-104983648;
#10;x=-104883648;
#10;x=-104783648;
#10;x=-104683648;
#10;x=-104583648;
#10;x=-104483648;
#10;x=-104383648;
#10;x=-104283648;
#10;x=-104183648;
#10;x=-104083648;
#10;x=-103983648;
#10;x=-103883648;
#10;x=-103783648;
#10;x=-103683648;
#10;x=-103583648;
#10;x=-103483648;
#10;x=-103383648;
#10;x=-103283648;
#10;x=-103183648;
#10;x=-103083648;
#10;x=-102983648;
#10;x=-102883648;
#10;x=-102783648;
#10;x=-102683648;
#10;x=-102583648;
#10;x=-102483648;
#10;x=-102383648;
#10;x=-102283648;
#10;x=-102183648;
#10;x=-102083648;
#10;x=-101983648;
#10;x=-101883648;
#10;x=-101783648;
#10;x=-101683648;
#10;x=-101583648;
#10;x=-101483648;
#10;x=-101383648;
#10;x=-101283648;
#10;x=-101183648;
#10;x=-101083648;
#10;x=-100983648;
#10;x=-100883648;
#10;x=-100783648;
#10;x=-100683648;
#10;x=-100583648;
#10;x=-100483648;
#10;x=-100383648;
#10;x=-100283648;
#10;x=-100183648;
#10;x=-100083648;
#10;x=-99983648;
#10;x=-99883648;
#10;x=-99783648;
#10;x=-99683648;
#10;x=-99583648;
#10;x=-99483648;
#10;x=-99383648;
#10;x=-99283648;
#10;x=-99183648;
#10;x=-99083648;
#10;x=-98983648;
#10;x=-98883648;
#10;x=-98783648;
#10;x=-98683648;
#10;x=-98583648;
#10;x=-98483648;
#10;x=-98383648;
#10;x=-98283648;
#10;x=-98183648;
#10;x=-98083648;
#10;x=-97983648;
#10;x=-97883648;
#10;x=-97783648;
#10;x=-97683648;
#10;x=-97583648;
#10;x=-97483648;
#10;x=-97383648;
#10;x=-97283648;
#10;x=-97183648;
#10;x=-97083648;
#10;x=-96983648;
#10;x=-96883648;
#10;x=-96783648;
#10;x=-96683648;
#10;x=-96583648;
#10;x=-96483648;
#10;x=-96383648;
#10;x=-96283648;
#10;x=-96183648;
#10;x=-96083648;
#10;x=-95983648;
#10;x=-95883648;
#10;x=-95783648;
#10;x=-95683648;
#10;x=-95583648;
#10;x=-95483648;
#10;x=-95383648;
#10;x=-95283648;
#10;x=-95183648;
#10;x=-95083648;
#10;x=-94983648;
#10;x=-94883648;
#10;x=-94783648;
#10;x=-94683648;
#10;x=-94583648;
#10;x=-94483648;
#10;x=-94383648;
#10;x=-94283648;
#10;x=-94183648;
#10;x=-94083648;
#10;x=-93983648;
#10;x=-93883648;
#10;x=-93783648;
#10;x=-93683648;
#10;x=-93583648;
#10;x=-93483648;
#10;x=-93383648;
#10;x=-93283648;
#10;x=-93183648;
#10;x=-93083648;
#10;x=-92983648;
#10;x=-92883648;
#10;x=-92783648;
#10;x=-92683648;
#10;x=-92583648;
#10;x=-92483648;
#10;x=-92383648;
#10;x=-92283648;
#10;x=-92183648;
#10;x=-92083648;
#10;x=-91983648;
#10;x=-91883648;
#10;x=-91783648;
#10;x=-91683648;
#10;x=-91583648;
#10;x=-91483648;
#10;x=-91383648;
#10;x=-91283648;
#10;x=-91183648;
#10;x=-91083648;
#10;x=-90983648;
#10;x=-90883648;
#10;x=-90783648;
#10;x=-90683648;
#10;x=-90583648;
#10;x=-90483648;
#10;x=-90383648;
#10;x=-90283648;
#10;x=-90183648;
#10;x=-90083648;
#10;x=-89983648;
#10;x=-89883648;
#10;x=-89783648;
#10;x=-89683648;
#10;x=-89583648;
#10;x=-89483648;
#10;x=-89383648;
#10;x=-89283648;
#10;x=-89183648;
#10;x=-89083648;
#10;x=-88983648;
#10;x=-88883648;
#10;x=-88783648;
#10;x=-88683648;
#10;x=-88583648;
#10;x=-88483648;
#10;x=-88383648;
#10;x=-88283648;
#10;x=-88183648;
#10;x=-88083648;
#10;x=-87983648;
#10;x=-87883648;
#10;x=-87783648;
#10;x=-87683648;
#10;x=-87583648;
#10;x=-87483648;
#10;x=-87383648;
#10;x=-87283648;
#10;x=-87183648;
#10;x=-87083648;
#10;x=-86983648;
#10;x=-86883648;
#10;x=-86783648;
#10;x=-86683648;
#10;x=-86583648;
#10;x=-86483648;
#10;x=-86383648;
#10;x=-86283648;
#10;x=-86183648;
#10;x=-86083648;
#10;x=-85983648;
#10;x=-85883648;
#10;x=-85783648;
#10;x=-85683648;
#10;x=-85583648;
#10;x=-85483648;
#10;x=-85383648;
#10;x=-85283648;
#10;x=-85183648;
#10;x=-85083648;
#10;x=-84983648;
#10;x=-84883648;
#10;x=-84783648;
#10;x=-84683648;
#10;x=-84583648;
#10;x=-84483648;
#10;x=-84383648;
#10;x=-84283648;
#10;x=-84183648;
#10;x=-84083648;
#10;x=-83983648;
#10;x=-83883648;
#10;x=-83783648;
#10;x=-83683648;
#10;x=-83583648;
#10;x=-83483648;
#10;x=-83383648;
#10;x=-83283648;
#10;x=-83183648;
#10;x=-83083648;
#10;x=-82983648;
#10;x=-82883648;
#10;x=-82783648;
#10;x=-82683648;
#10;x=-82583648;
#10;x=-82483648;
#10;x=-82383648;
#10;x=-82283648;
#10;x=-82183648;
#10;x=-82083648;
#10;x=-81983648;
#10;x=-81883648;
#10;x=-81783648;
#10;x=-81683648;
#10;x=-81583648;
#10;x=-81483648;
#10;x=-81383648;
#10;x=-81283648;
#10;x=-81183648;
#10;x=-81083648;
#10;x=-80983648;
#10;x=-80883648;
#10;x=-80783648;
#10;x=-80683648;
#10;x=-80583648;
#10;x=-80483648;
#10;x=-80383648;
#10;x=-80283648;
#10;x=-80183648;
#10;x=-80083648;
#10;x=-79983648;
#10;x=-79883648;
#10;x=-79783648;
#10;x=-79683648;
#10;x=-79583648;
#10;x=-79483648;
#10;x=-79383648;
#10;x=-79283648;
#10;x=-79183648;
#10;x=-79083648;
#10;x=-78983648;
#10;x=-78883648;
#10;x=-78783648;
#10;x=-78683648;
#10;x=-78583648;
#10;x=-78483648;
#10;x=-78383648;
#10;x=-78283648;
#10;x=-78183648;
#10;x=-78083648;
#10;x=-77983648;
#10;x=-77883648;
#10;x=-77783648;
#10;x=-77683648;
#10;x=-77583648;
#10;x=-77483648;
#10;x=-77383648;
#10;x=-77283648;
#10;x=-77183648;
#10;x=-77083648;
#10;x=-76983648;
#10;x=-76883648;
#10;x=-76783648;
#10;x=-76683648;
#10;x=-76583648;
#10;x=-76483648;
#10;x=-76383648;
#10;x=-76283648;
#10;x=-76183648;
#10;x=-76083648;
#10;x=-75983648;
#10;x=-75883648;
#10;x=-75783648;
#10;x=-75683648;
#10;x=-75583648;
#10;x=-75483648;
#10;x=-75383648;
#10;x=-75283648;
#10;x=-75183648;
#10;x=-75083648;
#10;x=-74983648;
#10;x=-74883648;
#10;x=-74783648;
#10;x=-74683648;
#10;x=-74583648;
#10;x=-74483648;
#10;x=-74383648;
#10;x=-74283648;
#10;x=-74183648;
#10;x=-74083648;
#10;x=-73983648;
#10;x=-73883648;
#10;x=-73783648;
#10;x=-73683648;
#10;x=-73583648;
#10;x=-73483648;
#10;x=-73383648;
#10;x=-73283648;
#10;x=-73183648;
#10;x=-73083648;
#10;x=-72983648;
#10;x=-72883648;
#10;x=-72783648;
#10;x=-72683648;
#10;x=-72583648;
#10;x=-72483648;
#10;x=-72383648;
#10;x=-72283648;
#10;x=-72183648;
#10;x=-72083648;
#10;x=-71983648;
#10;x=-71883648;
#10;x=-71783648;
#10;x=-71683648;
#10;x=-71583648;
#10;x=-71483648;
#10;x=-71383648;
#10;x=-71283648;
#10;x=-71183648;
#10;x=-71083648;
#10;x=-70983648;
#10;x=-70883648;
#10;x=-70783648;
#10;x=-70683648;
#10;x=-70583648;
#10;x=-70483648;
#10;x=-70383648;
#10;x=-70283648;
#10;x=-70183648;
#10;x=-70083648;
#10;x=-69983648;
#10;x=-69883648;
#10;x=-69783648;
#10;x=-69683648;
#10;x=-69583648;
#10;x=-69483648;
#10;x=-69383648;
#10;x=-69283648;
#10;x=-69183648;
#10;x=-69083648;
#10;x=-68983648;
#10;x=-68883648;
#10;x=-68783648;
#10;x=-68683648;
#10;x=-68583648;
#10;x=-68483648;
#10;x=-68383648;
#10;x=-68283648;
#10;x=-68183648;
#10;x=-68083648;
#10;x=-67983648;
#10;x=-67883648;
#10;x=-67783648;
#10;x=-67683648;
#10;x=-67583648;
#10;x=-67483648;
#10;x=-67383648;
#10;x=-67283648;
#10;x=-67183648;
#10;x=-67083648;
#10;x=-66983648;
#10;x=-66883648;
#10;x=-66783648;
#10;x=-66683648;
#10;x=-66583648;
#10;x=-66483648;
#10;x=-66383648;
#10;x=-66283648;
#10;x=-66183648;
#10;x=-66083648;
#10;x=-65983648;
#10;x=-65883648;
#10;x=-65783648;
#10;x=-65683648;
#10;x=-65583648;
#10;x=-65483648;
#10;x=-65383648;
#10;x=-65283648;
#10;x=-65183648;
#10;x=-65083648;
#10;x=-64983648;
#10;x=-64883648;
#10;x=-64783648;
#10;x=-64683648;
#10;x=-64583648;
#10;x=-64483648;
#10;x=-64383648;
#10;x=-64283648;
#10;x=-64183648;
#10;x=-64083648;
#10;x=-63983648;
#10;x=-63883648;
#10;x=-63783648;
#10;x=-63683648;
#10;x=-63583648;
#10;x=-63483648;
#10;x=-63383648;
#10;x=-63283648;
#10;x=-63183648;
#10;x=-63083648;
#10;x=-62983648;
#10;x=-62883648;
#10;x=-62783648;
#10;x=-62683648;
#10;x=-62583648;
#10;x=-62483648;
#10;x=-62383648;
#10;x=-62283648;
#10;x=-62183648;
#10;x=-62083648;
#10;x=-61983648;
#10;x=-61883648;
#10;x=-61783648;
#10;x=-61683648;
#10;x=-61583648;
#10;x=-61483648;
#10;x=-61383648;
#10;x=-61283648;
#10;x=-61183648;
#10;x=-61083648;
#10;x=-60983648;
#10;x=-60883648;
#10;x=-60783648;
#10;x=-60683648;
#10;x=-60583648;
#10;x=-60483648;
#10;x=-60383648;
#10;x=-60283648;
#10;x=-60183648;
#10;x=-60083648;
#10;x=-59983648;
#10;x=-59883648;
#10;x=-59783648;
#10;x=-59683648;
#10;x=-59583648;
#10;x=-59483648;
#10;x=-59383648;
#10;x=-59283648;
#10;x=-59183648;
#10;x=-59083648;
#10;x=-58983648;
#10;x=-58883648;
#10;x=-58783648;
#10;x=-58683648;
#10;x=-58583648;
#10;x=-58483648;
#10;x=-58383648;
#10;x=-58283648;
#10;x=-58183648;
#10;x=-58083648;
#10;x=-57983648;
#10;x=-57883648;
#10;x=-57783648;
#10;x=-57683648;
#10;x=-57583648;
#10;x=-57483648;
#10;x=-57383648;
#10;x=-57283648;
#10;x=-57183648;
#10;x=-57083648;
#10;x=-56983648;
#10;x=-56883648;
#10;x=-56783648;
#10;x=-56683648;
#10;x=-56583648;
#10;x=-56483648;
#10;x=-56383648;
#10;x=-56283648;
#10;x=-56183648;
#10;x=-56083648;
#10;x=-55983648;
#10;x=-55883648;
#10;x=-55783648;
#10;x=-55683648;
#10;x=-55583648;
#10;x=-55483648;
#10;x=-55383648;
#10;x=-55283648;
#10;x=-55183648;
#10;x=-55083648;
#10;x=-54983648;
#10;x=-54883648;
#10;x=-54783648;
#10;x=-54683648;
#10;x=-54583648;
#10;x=-54483648;
#10;x=-54383648;
#10;x=-54283648;
#10;x=-54183648;
#10;x=-54083648;
#10;x=-53983648;
#10;x=-53883648;
#10;x=-53783648;
#10;x=-53683648;
#10;x=-53583648;
#10;x=-53483648;
#10;x=-53383648;
#10;x=-53283648;
#10;x=-53183648;
#10;x=-53083648;
#10;x=-52983648;
#10;x=-52883648;
#10;x=-52783648;
#10;x=-52683648;
#10;x=-52583648;
#10;x=-52483648;
#10;x=-52383648;
#10;x=-52283648;
#10;x=-52183648;
#10;x=-52083648;
#10;x=-51983648;
#10;x=-51883648;
#10;x=-51783648;
#10;x=-51683648;
#10;x=-51583648;
#10;x=-51483648;
#10;x=-51383648;
#10;x=-51283648;
#10;x=-51183648;
#10;x=-51083648;
#10;x=-50983648;
#10;x=-50883648;
#10;x=-50783648;
#10;x=-50683648;
#10;x=-50583648;
#10;x=-50483648;
#10;x=-50383648;
#10;x=-50283648;
#10;x=-50183648;
#10;x=-50083648;
#10;x=-49983648;
#10;x=-49883648;
#10;x=-49783648;
#10;x=-49683648;
#10;x=-49583648;
#10;x=-49483648;
#10;x=-49383648;
#10;x=-49283648;
#10;x=-49183648;
#10;x=-49083648;
#10;x=-48983648;
#10;x=-48883648;
#10;x=-48783648;
#10;x=-48683648;
#10;x=-48583648;
#10;x=-48483648;
#10;x=-48383648;
#10;x=-48283648;
#10;x=-48183648;
#10;x=-48083648;
#10;x=-47983648;
#10;x=-47883648;
#10;x=-47783648;
#10;x=-47683648;
#10;x=-47583648;
#10;x=-47483648;
#10;x=-47383648;
#10;x=-47283648;
#10;x=-47183648;
#10;x=-47083648;
#10;x=-46983648;
#10;x=-46883648;
#10;x=-46783648;
#10;x=-46683648;
#10;x=-46583648;
#10;x=-46483648;
#10;x=-46383648;
#10;x=-46283648;
#10;x=-46183648;
#10;x=-46083648;
#10;x=-45983648;
#10;x=-45883648;
#10;x=-45783648;
#10;x=-45683648;
#10;x=-45583648;
#10;x=-45483648;
#10;x=-45383648;
#10;x=-45283648;
#10;x=-45183648;
#10;x=-45083648;
#10;x=-44983648;
#10;x=-44883648;
#10;x=-44783648;
#10;x=-44683648;
#10;x=-44583648;
#10;x=-44483648;
#10;x=-44383648;
#10;x=-44283648;
#10;x=-44183648;
#10;x=-44083648;
#10;x=-43983648;
#10;x=-43883648;
#10;x=-43783648;
#10;x=-43683648;
#10;x=-43583648;
#10;x=-43483648;
#10;x=-43383648;
#10;x=-43283648;
#10;x=-43183648;
#10;x=-43083648;
#10;x=-42983648;
#10;x=-42883648;
#10;x=-42783648;
#10;x=-42683648;
#10;x=-42583648;
#10;x=-42483648;
#10;x=-42383648;
#10;x=-42283648;
#10;x=-42183648;
#10;x=-42083648;
#10;x=-41983648;
#10;x=-41883648;
#10;x=-41783648;
#10;x=-41683648;
#10;x=-41583648;
#10;x=-41483648;
#10;x=-41383648;
#10;x=-41283648;
#10;x=-41183648;
#10;x=-41083648;
#10;x=-40983648;
#10;x=-40883648;
#10;x=-40783648;
#10;x=-40683648;
#10;x=-40583648;
#10;x=-40483648;
#10;x=-40383648;
#10;x=-40283648;
#10;x=-40183648;
#10;x=-40083648;
#10;x=-39983648;
#10;x=-39883648;
#10;x=-39783648;
#10;x=-39683648;
#10;x=-39583648;
#10;x=-39483648;
#10;x=-39383648;
#10;x=-39283648;
#10;x=-39183648;
#10;x=-39083648;
#10;x=-38983648;
#10;x=-38883648;
#10;x=-38783648;
#10;x=-38683648;
#10;x=-38583648;
#10;x=-38483648;
#10;x=-38383648;
#10;x=-38283648;
#10;x=-38183648;
#10;x=-38083648;
#10;x=-37983648;
#10;x=-37883648;
#10;x=-37783648;
#10;x=-37683648;
#10;x=-37583648;
#10;x=-37483648;
#10;x=-37383648;
#10;x=-37283648;
#10;x=-37183648;
#10;x=-37083648;
#10;x=-36983648;
#10;x=-36883648;
#10;x=-36783648;
#10;x=-36683648;
#10;x=-36583648;
#10;x=-36483648;
#10;x=-36383648;
#10;x=-36283648;
#10;x=-36183648;
#10;x=-36083648;
#10;x=-35983648;
#10;x=-35883648;
#10;x=-35783648;
#10;x=-35683648;
#10;x=-35583648;
#10;x=-35483648;
#10;x=-35383648;
#10;x=-35283648;
#10;x=-35183648;
#10;x=-35083648;
#10;x=-34983648;
#10;x=-34883648;
#10;x=-34783648;
#10;x=-34683648;
#10;x=-34583648;
#10;x=-34483648;
#10;x=-34383648;
#10;x=-34283648;
#10;x=-34183648;
#10;x=-34083648;
#10;x=-33983648;
#10;x=-33883648;
#10;x=-33783648;
#10;x=-33683648;
#10;x=-33583648;
#10;x=-33483648;
#10;x=-33383648;
#10;x=-33283648;
#10;x=-33183648;
#10;x=-33083648;
#10;x=-32983648;
#10;x=-32883648;
#10;x=-32783648;
#10;x=-32683648;
#10;x=-32583648;
#10;x=-32483648;
#10;x=-32383648;
#10;x=-32283648;
#10;x=-32183648;
#10;x=-32083648;
#10;x=-31983648;
#10;x=-31883648;
#10;x=-31783648;
#10;x=-31683648;
#10;x=-31583648;
#10;x=-31483648;
#10;x=-31383648;
#10;x=-31283648;
#10;x=-31183648;
#10;x=-31083648;
#10;x=-30983648;
#10;x=-30883648;
#10;x=-30783648;
#10;x=-30683648;
#10;x=-30583648;
#10;x=-30483648;
#10;x=-30383648;
#10;x=-30283648;
#10;x=-30183648;
#10;x=-30083648;
#10;x=-29983648;
#10;x=-29883648;
#10;x=-29783648;
#10;x=-29683648;
#10;x=-29583648;
#10;x=-29483648;
#10;x=-29383648;
#10;x=-29283648;
#10;x=-29183648;
#10;x=-29083648;
#10;x=-28983648;
#10;x=-28883648;
#10;x=-28783648;
#10;x=-28683648;
#10;x=-28583648;
#10;x=-28483648;
#10;x=-28383648;
#10;x=-28283648;
#10;x=-28183648;
#10;x=-28083648;
#10;x=-27983648;
#10;x=-27883648;
#10;x=-27783648;
#10;x=-27683648;
#10;x=-27583648;
#10;x=-27483648;
#10;x=-27383648;
#10;x=-27283648;
#10;x=-27183648;
#10;x=-27083648;
#10;x=-26983648;
#10;x=-26883648;
#10;x=-26783648;
#10;x=-26683648;
#10;x=-26583648;
#10;x=-26483648;
#10;x=-26383648;
#10;x=-26283648;
#10;x=-26183648;
#10;x=-26083648;
#10;x=-25983648;
#10;x=-25883648;
#10;x=-25783648;
#10;x=-25683648;
#10;x=-25583648;
#10;x=-25483648;
#10;x=-25383648;
#10;x=-25283648;
#10;x=-25183648;
#10;x=-25083648;
#10;x=-24983648;
#10;x=-24883648;
#10;x=-24783648;
#10;x=-24683648;
#10;x=-24583648;
#10;x=-24483648;
#10;x=-24383648;
#10;x=-24283648;
#10;x=-24183648;
#10;x=-24083648;
#10;x=-23983648;
#10;x=-23883648;
#10;x=-23783648;
#10;x=-23683648;
#10;x=-23583648;
#10;x=-23483648;
#10;x=-23383648;
#10;x=-23283648;
#10;x=-23183648;
#10;x=-23083648;
#10;x=-22983648;
#10;x=-22883648;
#10;x=-22783648;
#10;x=-22683648;
#10;x=-22583648;
#10;x=-22483648;
#10;x=-22383648;
#10;x=-22283648;
#10;x=-22183648;
#10;x=-22083648;
#10;x=-21983648;
#10;x=-21883648;
#10;x=-21783648;
#10;x=-21683648;
#10;x=-21583648;
#10;x=-21483648;
#10;x=-21383648;
#10;x=-21283648;
#10;x=-21183648;
#10;x=-21083648;
#10;x=-20983648;
#10;x=-20883648;
#10;x=-20783648;
#10;x=-20683648;
#10;x=-20583648;
#10;x=-20483648;
#10;x=-20383648;
#10;x=-20283648;
#10;x=-20183648;
#10;x=-20083648;
#10;x=-19983648;
#10;x=-19883648;
#10;x=-19783648;
#10;x=-19683648;
#10;x=-19583648;
#10;x=-19483648;
#10;x=-19383648;
#10;x=-19283648;
#10;x=-19183648;
#10;x=-19083648;
#10;x=-18983648;
#10;x=-18883648;
#10;x=-18783648;
#10;x=-18683648;
#10;x=-18583648;
#10;x=-18483648;
#10;x=-18383648;
#10;x=-18283648;
#10;x=-18183648;
#10;x=-18083648;
#10;x=-17983648;
#10;x=-17883648;
#10;x=-17783648;
#10;x=-17683648;
#10;x=-17583648;
#10;x=-17483648;
#10;x=-17383648;
#10;x=-17283648;
#10;x=-17183648;
#10;x=-17083648;
#10;x=-16983648;
#10;x=-16883648;
#10;x=-16783648;
#10;x=-16683648;
#10;x=-16583648;
#10;x=-16483648;
#10;x=-16383648;
#10;x=-16283648;
#10;x=-16183648;
#10;x=-16083648;
#10;x=-15983648;
#10;x=-15883648;
#10;x=-15783648;
#10;x=-15683648;
#10;x=-15583648;
#10;x=-15483648;
#10;x=-15383648;
#10;x=-15283648;
#10;x=-15183648;
#10;x=-15083648;
#10;x=-14983648;
#10;x=-14883648;
#10;x=-14783648;
#10;x=-14683648;
#10;x=-14583648;
#10;x=-14483648;
#10;x=-14383648;
#10;x=-14283648;
#10;x=-14183648;
#10;x=-14083648;
#10;x=-13983648;
#10;x=-13883648;
#10;x=-13783648;
#10;x=-13683648;
#10;x=-13583648;
#10;x=-13483648;
#10;x=-13383648;
#10;x=-13283648;
#10;x=-13183648;
#10;x=-13083648;
#10;x=-12983648;
#10;x=-12883648;
#10;x=-12783648;
#10;x=-12683648;
#10;x=-12583648;
#10;x=-12483648;
#10;x=-12383648;
#10;x=-12283648;
#10;x=-12183648;
#10;x=-12083648;
#10;x=-11983648;
#10;x=-11883648;
#10;x=-11783648;
#10;x=-11683648;
#10;x=-11583648;
#10;x=-11483648;
#10;x=-11383648;
#10;x=-11283648;
#10;x=-11183648;
#10;x=-11083648;
#10;x=-10983648;
#10;x=-10883648;
#10;x=-10783648;
#10;x=-10683648;
#10;x=-10583648;
#10;x=-10483648;
#10;x=-10383648;
#10;x=-10283648;
#10;x=-10183648;
#10;x=-10083648;
#10;x=-9983648;
#10;x=-9883648;
#10;x=-9783648;
#10;x=-9683648;
#10;x=-9583648;
#10;x=-9483648;
#10;x=-9383648;
#10;x=-9283648;
#10;x=-9183648;
#10;x=-9083648;
#10;x=-8983648;
#10;x=-8883648;
#10;x=-8783648;
#10;x=-8683648;
#10;x=-8583648;
#10;x=-8483648;
#10;x=-8383648;
#10;x=-8283648;
#10;x=-8183648;
#10;x=-8083648;
#10;x=-7983648;
#10;x=-7883648;
#10;x=-7783648;
#10;x=-7683648;
#10;x=-7583648;
#10;x=-7483648;
#10;x=-7383648;
#10;x=-7283648;
#10;x=-7183648;
#10;x=-7083648;
#10;x=-6983648;
#10;x=-6883648;
#10;x=-6783648;
#10;x=-6683648;
#10;x=-6583648;
#10;x=-6483648;
#10;x=-6383648;
#10;x=-6283648;
#10;x=-6183648;
#10;x=-6083648;
#10;x=-5983648;
#10;x=-5883648;
#10;x=-5783648;
#10;x=-5683648;
#10;x=-5583648;
#10;x=-5483648;
#10;x=-5383648;
#10;x=-5283648;
#10;x=-5183648;
#10;x=-5083648;
#10;x=-4983648;
#10;x=-4883648;
#10;x=-4783648;
#10;x=-4683648;
#10;x=-4583648;
#10;x=-4483648;
#10;x=-4383648;
#10;x=-4283648;
#10;x=-4183648;
#10;x=-4083648;
#10;x=-3983648;
#10;x=-3883648;
#10;x=-3783648;
#10;x=-3683648;
#10;x=-3583648;
#10;x=-3483648;
#10;x=-3383648;
#10;x=-3283648;
#10;x=-3183648;
#10;x=-3083648;
#10;x=-2983648;
#10;x=-2883648;
#10;x=-2783648;
#10;x=-2683648;
#10;x=-2583648;
#10;x=-2483648;
#10;x=-2383648;
#10;x=-2283648;
#10;x=-2183648;
#10;x=-2083648;
#10;x=-1983648;
#10;x=-1883648;
#10;x=-1783648;
#10;x=-1683648;
#10;x=-1583648;
#10;x=-1483648;
#10;x=-1383648;
#10;x=-1283648;
#10;x=-1183648;
#10;x=-1083648;
#10;x=-983648;
#10;x=-883648;
#10;x=-783648;
#10;x=-683648;
#10;x=-583648;
#10;x=-483648;
#10;x=-383648;
#10;x=-283648;
#10;x=-183648;
#10;x=-83648;
#10;x=16352;
#10;x=116352;
#10;x=216352;
#10;x=316352;
#10;x=416352;
#10;x=516352;
#10;x=616352;
#10;x=716352;
#10;x=816352;
#10;x=916352;
#10;x=1016352;
#10;x=1116352;
#10;x=1216352;
#10;x=1316352;
#10;x=1416352;
#10;x=1516352;
#10;x=1616352;
#10;x=1716352;
#10;x=1816352;
#10;x=1916352;
#10;x=2016352;
#10;x=2116352;
#10;x=2216352;
#10;x=2316352;
#10;x=2416352;
#10;x=2516352;
#10;x=2616352;
#10;x=2716352;
#10;x=2816352;
#10;x=2916352;
#10;x=3016352;
#10;x=3116352;
#10;x=3216352;
#10;x=3316352;
#10;x=3416352;
#10;x=3516352;
#10;x=3616352;
#10;x=3716352;
#10;x=3816352;
#10;x=3916352;
#10;x=4016352;
#10;x=4116352;
#10;x=4216352;
#10;x=4316352;
#10;x=4416352;
#10;x=4516352;
#10;x=4616352;
#10;x=4716352;
#10;x=4816352;
#10;x=4916352;
#10;x=5016352;
#10;x=5116352;
#10;x=5216352;
#10;x=5316352;
#10;x=5416352;
#10;x=5516352;
#10;x=5616352;
#10;x=5716352;
#10;x=5816352;
#10;x=5916352;
#10;x=6016352;
#10;x=6116352;
#10;x=6216352;
#10;x=6316352;
#10;x=6416352;
#10;x=6516352;
#10;x=6616352;
#10;x=6716352;
#10;x=6816352;
#10;x=6916352;
#10;x=7016352;
#10;x=7116352;
#10;x=7216352;
#10;x=7316352;
#10;x=7416352;
#10;x=7516352;
#10;x=7616352;
#10;x=7716352;
#10;x=7816352;
#10;x=7916352;
#10;x=8016352;
#10;x=8116352;
#10;x=8216352;
#10;x=8316352;
#10;x=8416352;
#10;x=8516352;
#10;x=8616352;
#10;x=8716352;
#10;x=8816352;
#10;x=8916352;
#10;x=9016352;
#10;x=9116352;
#10;x=9216352;
#10;x=9316352;
#10;x=9416352;
#10;x=9516352;
#10;x=9616352;
#10;x=9716352;
#10;x=9816352;
#10;x=9916352;
#10;x=10016352;
#10;x=10116352;
#10;x=10216352;
#10;x=10316352;
#10;x=10416352;
#10;x=10516352;
#10;x=10616352;
#10;x=10716352;
#10;x=10816352;
#10;x=10916352;
#10;x=11016352;
#10;x=11116352;
#10;x=11216352;
#10;x=11316352;
#10;x=11416352;
#10;x=11516352;
#10;x=11616352;
#10;x=11716352;
#10;x=11816352;
#10;x=11916352;
#10;x=12016352;
#10;x=12116352;
#10;x=12216352;
#10;x=12316352;
#10;x=12416352;
#10;x=12516352;
#10;x=12616352;
#10;x=12716352;
#10;x=12816352;
#10;x=12916352;
#10;x=13016352;
#10;x=13116352;
#10;x=13216352;
#10;x=13316352;
#10;x=13416352;
#10;x=13516352;
#10;x=13616352;
#10;x=13716352;
#10;x=13816352;
#10;x=13916352;
#10;x=14016352;
#10;x=14116352;
#10;x=14216352;
#10;x=14316352;
#10;x=14416352;
#10;x=14516352;
#10;x=14616352;
#10;x=14716352;
#10;x=14816352;
#10;x=14916352;
#10;x=15016352;
#10;x=15116352;
#10;x=15216352;
#10;x=15316352;
#10;x=15416352;
#10;x=15516352;
#10;x=15616352;
#10;x=15716352;
#10;x=15816352;
#10;x=15916352;
#10;x=16016352;
#10;x=16116352;
#10;x=16216352;
#10;x=16316352;
#10;x=16416352;
#10;x=16516352;
#10;x=16616352;
#10;x=16716352;
#10;x=16816352;
#10;x=16916352;
#10;x=17016352;
#10;x=17116352;
#10;x=17216352;
#10;x=17316352;
#10;x=17416352;
#10;x=17516352;
#10;x=17616352;
#10;x=17716352;
#10;x=17816352;
#10;x=17916352;
#10;x=18016352;
#10;x=18116352;
#10;x=18216352;
#10;x=18316352;
#10;x=18416352;
#10;x=18516352;
#10;x=18616352;
#10;x=18716352;
#10;x=18816352;
#10;x=18916352;
#10;x=19016352;
#10;x=19116352;
#10;x=19216352;
#10;x=19316352;
#10;x=19416352;
#10;x=19516352;
#10;x=19616352;
#10;x=19716352;
#10;x=19816352;
#10;x=19916352;
#10;x=20016352;
#10;x=20116352;
#10;x=20216352;
#10;x=20316352;
#10;x=20416352;
#10;x=20516352;
#10;x=20616352;
#10;x=20716352;
#10;x=20816352;
#10;x=20916352;
#10;x=21016352;
#10;x=21116352;
#10;x=21216352;
#10;x=21316352;
#10;x=21416352;
#10;x=21516352;
#10;x=21616352;
#10;x=21716352;
#10;x=21816352;
#10;x=21916352;
#10;x=22016352;
#10;x=22116352;
#10;x=22216352;
#10;x=22316352;
#10;x=22416352;
#10;x=22516352;
#10;x=22616352;
#10;x=22716352;
#10;x=22816352;
#10;x=22916352;
#10;x=23016352;
#10;x=23116352;
#10;x=23216352;
#10;x=23316352;
#10;x=23416352;
#10;x=23516352;
#10;x=23616352;
#10;x=23716352;
#10;x=23816352;
#10;x=23916352;
#10;x=24016352;
#10;x=24116352;
#10;x=24216352;
#10;x=24316352;
#10;x=24416352;
#10;x=24516352;
#10;x=24616352;
#10;x=24716352;
#10;x=24816352;
#10;x=24916352;
#10;x=25016352;
#10;x=25116352;
#10;x=25216352;
#10;x=25316352;
#10;x=25416352;
#10;x=25516352;
#10;x=25616352;
#10;x=25716352;
#10;x=25816352;
#10;x=25916352;
#10;x=26016352;
#10;x=26116352;
#10;x=26216352;
#10;x=26316352;
#10;x=26416352;
#10;x=26516352;
#10;x=26616352;
#10;x=26716352;
#10;x=26816352;
#10;x=26916352;
#10;x=27016352;
#10;x=27116352;
#10;x=27216352;
#10;x=27316352;
#10;x=27416352;
#10;x=27516352;
#10;x=27616352;
#10;x=27716352;
#10;x=27816352;
#10;x=27916352;
#10;x=28016352;
#10;x=28116352;
#10;x=28216352;
#10;x=28316352;
#10;x=28416352;
#10;x=28516352;
#10;x=28616352;
#10;x=28716352;
#10;x=28816352;
#10;x=28916352;
#10;x=29016352;
#10;x=29116352;
#10;x=29216352;
#10;x=29316352;
#10;x=29416352;
#10;x=29516352;
#10;x=29616352;
#10;x=29716352;
#10;x=29816352;
#10;x=29916352;
#10;x=30016352;
#10;x=30116352;
#10;x=30216352;
#10;x=30316352;
#10;x=30416352;
#10;x=30516352;
#10;x=30616352;
#10;x=30716352;
#10;x=30816352;
#10;x=30916352;
#10;x=31016352;
#10;x=31116352;
#10;x=31216352;
#10;x=31316352;
#10;x=31416352;
#10;x=31516352;
#10;x=31616352;
#10;x=31716352;
#10;x=31816352;
#10;x=31916352;
#10;x=32016352;
#10;x=32116352;
#10;x=32216352;
#10;x=32316352;
#10;x=32416352;
#10;x=32516352;
#10;x=32616352;
#10;x=32716352;
#10;x=32816352;
#10;x=32916352;
#10;x=33016352;
#10;x=33116352;
#10;x=33216352;
#10;x=33316352;
#10;x=33416352;
#10;x=33516352;
#10;x=33616352;
#10;x=33716352;
#10;x=33816352;
#10;x=33916352;
#10;x=34016352;
#10;x=34116352;
#10;x=34216352;
#10;x=34316352;
#10;x=34416352;
#10;x=34516352;
#10;x=34616352;
#10;x=34716352;
#10;x=34816352;
#10;x=34916352;
#10;x=35016352;
#10;x=35116352;
#10;x=35216352;
#10;x=35316352;
#10;x=35416352;
#10;x=35516352;
#10;x=35616352;
#10;x=35716352;
#10;x=35816352;
#10;x=35916352;
#10;x=36016352;
#10;x=36116352;
#10;x=36216352;
#10;x=36316352;
#10;x=36416352;
#10;x=36516352;
#10;x=36616352;
#10;x=36716352;
#10;x=36816352;
#10;x=36916352;
#10;x=37016352;
#10;x=37116352;
#10;x=37216352;
#10;x=37316352;
#10;x=37416352;
#10;x=37516352;
#10;x=37616352;
#10;x=37716352;
#10;x=37816352;
#10;x=37916352;
#10;x=38016352;
#10;x=38116352;
#10;x=38216352;
#10;x=38316352;
#10;x=38416352;
#10;x=38516352;
#10;x=38616352;
#10;x=38716352;
#10;x=38816352;
#10;x=38916352;
#10;x=39016352;
#10;x=39116352;
#10;x=39216352;
#10;x=39316352;
#10;x=39416352;
#10;x=39516352;
#10;x=39616352;
#10;x=39716352;
#10;x=39816352;
#10;x=39916352;
#10;x=40016352;
#10;x=40116352;
#10;x=40216352;
#10;x=40316352;
#10;x=40416352;
#10;x=40516352;
#10;x=40616352;
#10;x=40716352;
#10;x=40816352;
#10;x=40916352;
#10;x=41016352;
#10;x=41116352;
#10;x=41216352;
#10;x=41316352;
#10;x=41416352;
#10;x=41516352;
#10;x=41616352;
#10;x=41716352;
#10;x=41816352;
#10;x=41916352;
#10;x=42016352;
#10;x=42116352;
#10;x=42216352;
#10;x=42316352;
#10;x=42416352;
#10;x=42516352;
#10;x=42616352;
#10;x=42716352;
#10;x=42816352;
#10;x=42916352;
#10;x=43016352;
#10;x=43116352;
#10;x=43216352;
#10;x=43316352;
#10;x=43416352;
#10;x=43516352;
#10;x=43616352;
#10;x=43716352;
#10;x=43816352;
#10;x=43916352;
#10;x=44016352;
#10;x=44116352;
#10;x=44216352;
#10;x=44316352;
#10;x=44416352;
#10;x=44516352;
#10;x=44616352;
#10;x=44716352;
#10;x=44816352;
#10;x=44916352;
#10;x=45016352;
#10;x=45116352;
#10;x=45216352;
#10;x=45316352;
#10;x=45416352;
#10;x=45516352;
#10;x=45616352;
#10;x=45716352;
#10;x=45816352;
#10;x=45916352;
#10;x=46016352;
#10;x=46116352;
#10;x=46216352;
#10;x=46316352;
#10;x=46416352;
#10;x=46516352;
#10;x=46616352;
#10;x=46716352;
#10;x=46816352;
#10;x=46916352;
#10;x=47016352;
#10;x=47116352;
#10;x=47216352;
#10;x=47316352;
#10;x=47416352;
#10;x=47516352;
#10;x=47616352;
#10;x=47716352;
#10;x=47816352;
#10;x=47916352;
#10;x=48016352;
#10;x=48116352;
#10;x=48216352;
#10;x=48316352;
#10;x=48416352;
#10;x=48516352;
#10;x=48616352;
#10;x=48716352;
#10;x=48816352;
#10;x=48916352;
#10;x=49016352;
#10;x=49116352;
#10;x=49216352;
#10;x=49316352;
#10;x=49416352;
#10;x=49516352;
#10;x=49616352;
#10;x=49716352;
#10;x=49816352;
#10;x=49916352;
#10;x=50016352;
#10;x=50116352;
#10;x=50216352;
#10;x=50316352;
#10;x=50416352;
#10;x=50516352;
#10;x=50616352;
#10;x=50716352;
#10;x=50816352;
#10;x=50916352;
#10;x=51016352;
#10;x=51116352;
#10;x=51216352;
#10;x=51316352;
#10;x=51416352;
#10;x=51516352;
#10;x=51616352;
#10;x=51716352;
#10;x=51816352;
#10;x=51916352;
#10;x=52016352;
#10;x=52116352;
#10;x=52216352;
#10;x=52316352;
#10;x=52416352;
#10;x=52516352;
#10;x=52616352;
#10;x=52716352;
#10;x=52816352;
#10;x=52916352;
#10;x=53016352;
#10;x=53116352;
#10;x=53216352;
#10;x=53316352;
#10;x=53416352;
#10;x=53516352;
#10;x=53616352;
#10;x=53716352;
#10;x=53816352;
#10;x=53916352;
#10;x=54016352;
#10;x=54116352;
#10;x=54216352;
#10;x=54316352;
#10;x=54416352;
#10;x=54516352;
#10;x=54616352;
#10;x=54716352;
#10;x=54816352;
#10;x=54916352;
#10;x=55016352;
#10;x=55116352;
#10;x=55216352;
#10;x=55316352;
#10;x=55416352;
#10;x=55516352;
#10;x=55616352;
#10;x=55716352;
#10;x=55816352;
#10;x=55916352;
#10;x=56016352;
#10;x=56116352;
#10;x=56216352;
#10;x=56316352;
#10;x=56416352;
#10;x=56516352;
#10;x=56616352;
#10;x=56716352;
#10;x=56816352;
#10;x=56916352;
#10;x=57016352;
#10;x=57116352;
#10;x=57216352;
#10;x=57316352;
#10;x=57416352;
#10;x=57516352;
#10;x=57616352;
#10;x=57716352;
#10;x=57816352;
#10;x=57916352;
#10;x=58016352;
#10;x=58116352;
#10;x=58216352;
#10;x=58316352;
#10;x=58416352;
#10;x=58516352;
#10;x=58616352;
#10;x=58716352;
#10;x=58816352;
#10;x=58916352;
#10;x=59016352;
#10;x=59116352;
#10;x=59216352;
#10;x=59316352;
#10;x=59416352;
#10;x=59516352;
#10;x=59616352;
#10;x=59716352;
#10;x=59816352;
#10;x=59916352;
#10;x=60016352;
#10;x=60116352;
#10;x=60216352;
#10;x=60316352;
#10;x=60416352;
#10;x=60516352;
#10;x=60616352;
#10;x=60716352;
#10;x=60816352;
#10;x=60916352;
#10;x=61016352;
#10;x=61116352;
#10;x=61216352;
#10;x=61316352;
#10;x=61416352;
#10;x=61516352;
#10;x=61616352;
#10;x=61716352;
#10;x=61816352;
#10;x=61916352;
#10;x=62016352;
#10;x=62116352;
#10;x=62216352;
#10;x=62316352;
#10;x=62416352;
#10;x=62516352;
#10;x=62616352;
#10;x=62716352;
#10;x=62816352;
#10;x=62916352;
#10;x=63016352;
#10;x=63116352;
#10;x=63216352;
#10;x=63316352;
#10;x=63416352;
#10;x=63516352;
#10;x=63616352;
#10;x=63716352;
#10;x=63816352;
#10;x=63916352;
#10;x=64016352;
#10;x=64116352;
#10;x=64216352;
#10;x=64316352;
#10;x=64416352;
#10;x=64516352;
#10;x=64616352;
#10;x=64716352;
#10;x=64816352;
#10;x=64916352;
#10;x=65016352;
#10;x=65116352;
#10;x=65216352;
#10;x=65316352;
#10;x=65416352;
#10;x=65516352;
#10;x=65616352;
#10;x=65716352;
#10;x=65816352;
#10;x=65916352;
#10;x=66016352;
#10;x=66116352;
#10;x=66216352;
#10;x=66316352;
#10;x=66416352;
#10;x=66516352;
#10;x=66616352;
#10;x=66716352;
#10;x=66816352;
#10;x=66916352;
#10;x=67016352;
#10;x=67116352;
#10;x=67216352;
#10;x=67316352;
#10;x=67416352;
#10;x=67516352;
#10;x=67616352;
#10;x=67716352;
#10;x=67816352;
#10;x=67916352;
#10;x=68016352;
#10;x=68116352;
#10;x=68216352;
#10;x=68316352;
#10;x=68416352;
#10;x=68516352;
#10;x=68616352;
#10;x=68716352;
#10;x=68816352;
#10;x=68916352;
#10;x=69016352;
#10;x=69116352;
#10;x=69216352;
#10;x=69316352;
#10;x=69416352;
#10;x=69516352;
#10;x=69616352;
#10;x=69716352;
#10;x=69816352;
#10;x=69916352;
#10;x=70016352;
#10;x=70116352;
#10;x=70216352;
#10;x=70316352;
#10;x=70416352;
#10;x=70516352;
#10;x=70616352;
#10;x=70716352;
#10;x=70816352;
#10;x=70916352;
#10;x=71016352;
#10;x=71116352;
#10;x=71216352;
#10;x=71316352;
#10;x=71416352;
#10;x=71516352;
#10;x=71616352;
#10;x=71716352;
#10;x=71816352;
#10;x=71916352;
#10;x=72016352;
#10;x=72116352;
#10;x=72216352;
#10;x=72316352;
#10;x=72416352;
#10;x=72516352;
#10;x=72616352;
#10;x=72716352;
#10;x=72816352;
#10;x=72916352;
#10;x=73016352;
#10;x=73116352;
#10;x=73216352;
#10;x=73316352;
#10;x=73416352;
#10;x=73516352;
#10;x=73616352;
#10;x=73716352;
#10;x=73816352;
#10;x=73916352;
#10;x=74016352;
#10;x=74116352;
#10;x=74216352;
#10;x=74316352;
#10;x=74416352;
#10;x=74516352;
#10;x=74616352;
#10;x=74716352;
#10;x=74816352;
#10;x=74916352;
#10;x=75016352;
#10;x=75116352;
#10;x=75216352;
#10;x=75316352;
#10;x=75416352;
#10;x=75516352;
#10;x=75616352;
#10;x=75716352;
#10;x=75816352;
#10;x=75916352;
#10;x=76016352;
#10;x=76116352;
#10;x=76216352;
#10;x=76316352;
#10;x=76416352;
#10;x=76516352;
#10;x=76616352;
#10;x=76716352;
#10;x=76816352;
#10;x=76916352;
#10;x=77016352;
#10;x=77116352;
#10;x=77216352;
#10;x=77316352;
#10;x=77416352;
#10;x=77516352;
#10;x=77616352;
#10;x=77716352;
#10;x=77816352;
#10;x=77916352;
#10;x=78016352;
#10;x=78116352;
#10;x=78216352;
#10;x=78316352;
#10;x=78416352;
#10;x=78516352;
#10;x=78616352;
#10;x=78716352;
#10;x=78816352;
#10;x=78916352;
#10;x=79016352;
#10;x=79116352;
#10;x=79216352;
#10;x=79316352;
#10;x=79416352;
#10;x=79516352;
#10;x=79616352;
#10;x=79716352;
#10;x=79816352;
#10;x=79916352;
#10;x=80016352;
#10;x=80116352;
#10;x=80216352;
#10;x=80316352;
#10;x=80416352;
#10;x=80516352;
#10;x=80616352;
#10;x=80716352;
#10;x=80816352;
#10;x=80916352;
#10;x=81016352;
#10;x=81116352;
#10;x=81216352;
#10;x=81316352;
#10;x=81416352;
#10;x=81516352;
#10;x=81616352;
#10;x=81716352;
#10;x=81816352;
#10;x=81916352;
#10;x=82016352;
#10;x=82116352;
#10;x=82216352;
#10;x=82316352;
#10;x=82416352;
#10;x=82516352;
#10;x=82616352;
#10;x=82716352;
#10;x=82816352;
#10;x=82916352;
#10;x=83016352;
#10;x=83116352;
#10;x=83216352;
#10;x=83316352;
#10;x=83416352;
#10;x=83516352;
#10;x=83616352;
#10;x=83716352;
#10;x=83816352;
#10;x=83916352;
#10;x=84016352;
#10;x=84116352;
#10;x=84216352;
#10;x=84316352;
#10;x=84416352;
#10;x=84516352;
#10;x=84616352;
#10;x=84716352;
#10;x=84816352;
#10;x=84916352;
#10;x=85016352;
#10;x=85116352;
#10;x=85216352;
#10;x=85316352;
#10;x=85416352;
#10;x=85516352;
#10;x=85616352;
#10;x=85716352;
#10;x=85816352;
#10;x=85916352;
#10;x=86016352;
#10;x=86116352;
#10;x=86216352;
#10;x=86316352;
#10;x=86416352;
#10;x=86516352;
#10;x=86616352;
#10;x=86716352;
#10;x=86816352;
#10;x=86916352;
#10;x=87016352;
#10;x=87116352;
#10;x=87216352;
#10;x=87316352;
#10;x=87416352;
#10;x=87516352;
#10;x=87616352;
#10;x=87716352;
#10;x=87816352;
#10;x=87916352;
#10;x=88016352;
#10;x=88116352;
#10;x=88216352;
#10;x=88316352;
#10;x=88416352;
#10;x=88516352;
#10;x=88616352;
#10;x=88716352;
#10;x=88816352;
#10;x=88916352;
#10;x=89016352;
#10;x=89116352;
#10;x=89216352;
#10;x=89316352;
#10;x=89416352;
#10;x=89516352;
#10;x=89616352;
#10;x=89716352;
#10;x=89816352;
#10;x=89916352;
#10;x=90016352;
#10;x=90116352;
#10;x=90216352;
#10;x=90316352;
#10;x=90416352;
#10;x=90516352;
#10;x=90616352;
#10;x=90716352;
#10;x=90816352;
#10;x=90916352;
#10;x=91016352;
#10;x=91116352;
#10;x=91216352;
#10;x=91316352;
#10;x=91416352;
#10;x=91516352;
#10;x=91616352;
#10;x=91716352;
#10;x=91816352;
#10;x=91916352;
#10;x=92016352;
#10;x=92116352;
#10;x=92216352;
#10;x=92316352;
#10;x=92416352;
#10;x=92516352;
#10;x=92616352;
#10;x=92716352;
#10;x=92816352;
#10;x=92916352;
#10;x=93016352;
#10;x=93116352;
#10;x=93216352;
#10;x=93316352;
#10;x=93416352;
#10;x=93516352;
#10;x=93616352;
#10;x=93716352;
#10;x=93816352;
#10;x=93916352;
#10;x=94016352;
#10;x=94116352;
#10;x=94216352;
#10;x=94316352;
#10;x=94416352;
#10;x=94516352;
#10;x=94616352;
#10;x=94716352;
#10;x=94816352;
#10;x=94916352;
#10;x=95016352;
#10;x=95116352;
#10;x=95216352;
#10;x=95316352;
#10;x=95416352;
#10;x=95516352;
#10;x=95616352;
#10;x=95716352;
#10;x=95816352;
#10;x=95916352;
#10;x=96016352;
#10;x=96116352;
#10;x=96216352;
#10;x=96316352;
#10;x=96416352;
#10;x=96516352;
#10;x=96616352;
#10;x=96716352;
#10;x=96816352;
#10;x=96916352;
#10;x=97016352;
#10;x=97116352;
#10;x=97216352;
#10;x=97316352;
#10;x=97416352;
#10;x=97516352;
#10;x=97616352;
#10;x=97716352;
#10;x=97816352;
#10;x=97916352;
#10;x=98016352;
#10;x=98116352;
#10;x=98216352;
#10;x=98316352;
#10;x=98416352;
#10;x=98516352;
#10;x=98616352;
#10;x=98716352;
#10;x=98816352;
#10;x=98916352;
#10;x=99016352;
#10;x=99116352;
#10;x=99216352;
#10;x=99316352;
#10;x=99416352;
#10;x=99516352;
#10;x=99616352;
#10;x=99716352;
#10;x=99816352;
#10;x=99916352;
#10;x=100016352;
#10;x=100116352;
#10;x=100216352;
#10;x=100316352;
#10;x=100416352;
#10;x=100516352;
#10;x=100616352;
#10;x=100716352;
#10;x=100816352;
#10;x=100916352;
#10;x=101016352;
#10;x=101116352;
#10;x=101216352;
#10;x=101316352;
#10;x=101416352;
#10;x=101516352;
#10;x=101616352;
#10;x=101716352;
#10;x=101816352;
#10;x=101916352;
#10;x=102016352;
#10;x=102116352;
#10;x=102216352;
#10;x=102316352;
#10;x=102416352;
#10;x=102516352;
#10;x=102616352;
#10;x=102716352;
#10;x=102816352;
#10;x=102916352;
#10;x=103016352;
#10;x=103116352;
#10;x=103216352;
#10;x=103316352;
#10;x=103416352;
#10;x=103516352;
#10;x=103616352;
#10;x=103716352;
#10;x=103816352;
#10;x=103916352;
#10;x=104016352;
#10;x=104116352;
#10;x=104216352;
#10;x=104316352;
#10;x=104416352;
#10;x=104516352;
#10;x=104616352;
#10;x=104716352;
#10;x=104816352;
#10;x=104916352;
#10;x=105016352;
#10;x=105116352;
#10;x=105216352;
#10;x=105316352;
#10;x=105416352;
#10;x=105516352;
#10;x=105616352;
#10;x=105716352;
#10;x=105816352;
#10;x=105916352;
#10;x=106016352;
#10;x=106116352;
#10;x=106216352;
#10;x=106316352;
#10;x=106416352;
#10;x=106516352;
#10;x=106616352;
#10;x=106716352;
#10;x=106816352;
#10;x=106916352;
#10;x=107016352;
#10;x=107116352;
#10;x=107216352;
#10;x=107316352;
#10;x=107416352;
#10;x=107516352;
#10;x=107616352;
#10;x=107716352;
#10;x=107816352;
#10;x=107916352;
#10;x=108016352;
#10;x=108116352;
#10;x=108216352;
#10;x=108316352;
#10;x=108416352;
#10;x=108516352;
#10;x=108616352;
#10;x=108716352;
#10;x=108816352;
#10;x=108916352;
#10;x=109016352;
#10;x=109116352;
#10;x=109216352;
#10;x=109316352;
#10;x=109416352;
#10;x=109516352;
#10;x=109616352;
#10;x=109716352;
#10;x=109816352;
#10;x=109916352;
#10;x=110016352;
#10;x=110116352;
#10;x=110216352;
#10;x=110316352;
#10;x=110416352;
#10;x=110516352;
#10;x=110616352;
#10;x=110716352;
#10;x=110816352;
#10;x=110916352;
#10;x=111016352;
#10;x=111116352;
#10;x=111216352;
#10;x=111316352;
#10;x=111416352;
#10;x=111516352;
#10;x=111616352;
#10;x=111716352;
#10;x=111816352;
#10;x=111916352;
#10;x=112016352;
#10;x=112116352;
#10;x=112216352;
#10;x=112316352;
#10;x=112416352;
#10;x=112516352;
#10;x=112616352;
#10;x=112716352;
#10;x=112816352;
#10;x=112916352;
#10;x=113016352;
#10;x=113116352;
#10;x=113216352;
#10;x=113316352;
#10;x=113416352;
#10;x=113516352;
#10;x=113616352;
#10;x=113716352;
#10;x=113816352;
#10;x=113916352;
#10;x=114016352;
#10;x=114116352;
#10;x=114216352;
#10;x=114316352;
#10;x=114416352;
#10;x=114516352;
#10;x=114616352;
#10;x=114716352;
#10;x=114816352;
#10;x=114916352;
#10;x=115016352;
#10;x=115116352;
#10;x=115216352;
#10;x=115316352;
#10;x=115416352;
#10;x=115516352;
#10;x=115616352;
#10;x=115716352;
#10;x=115816352;
#10;x=115916352;
#10;x=116016352;
#10;x=116116352;
#10;x=116216352;
#10;x=116316352;
#10;x=116416352;
#10;x=116516352;
#10;x=116616352;
#10;x=116716352;
#10;x=116816352;
#10;x=116916352;
#10;x=117016352;
#10;x=117116352;
#10;x=117216352;
#10;x=117316352;
#10;x=117416352;
#10;x=117516352;
#10;x=117616352;
#10;x=117716352;
#10;x=117816352;
#10;x=117916352;
#10;x=118016352;
#10;x=118116352;
#10;x=118216352;
#10;x=118316352;
#10;x=118416352;
#10;x=118516352;
#10;x=118616352;
#10;x=118716352;
#10;x=118816352;
#10;x=118916352;
#10;x=119016352;
#10;x=119116352;
#10;x=119216352;
#10;x=119316352;
#10;x=119416352;
#10;x=119516352;
#10;x=119616352;
#10;x=119716352;
#10;x=119816352;
#10;x=119916352;
#10;x=120016352;
#10;x=120116352;
#10;x=120216352;
#10;x=120316352;
#10;x=120416352;
#10;x=120516352;
#10;x=120616352;
#10;x=120716352;
#10;x=120816352;
#10;x=120916352;
#10;x=121016352;
#10;x=121116352;
#10;x=121216352;
#10;x=121316352;
#10;x=121416352;
#10;x=121516352;
#10;x=121616352;
#10;x=121716352;
#10;x=121816352;
#10;x=121916352;
#10;x=122016352;
#10;x=122116352;
#10;x=122216352;
#10;x=122316352;
#10;x=122416352;
#10;x=122516352;
#10;x=122616352;
#10;x=122716352;
#10;x=122816352;
#10;x=122916352;
#10;x=123016352;
#10;x=123116352;
#10;x=123216352;
#10;x=123316352;
#10;x=123416352;
#10;x=123516352;
#10;x=123616352;
#10;x=123716352;
#10;x=123816352;
#10;x=123916352;
#10;x=124016352;
#10;x=124116352;
#10;x=124216352;
#10;x=124316352;
#10;x=124416352;
#10;x=124516352;
#10;x=124616352;
#10;x=124716352;
#10;x=124816352;
#10;x=124916352;
#10;x=125016352;
#10;x=125116352;
#10;x=125216352;
#10;x=125316352;
#10;x=125416352;
#10;x=125516352;
#10;x=125616352;
#10;x=125716352;
#10;x=125816352;
#10;x=125916352;
#10;x=126016352;
#10;x=126116352;
#10;x=126216352;
#10;x=126316352;
#10;x=126416352;
#10;x=126516352;
#10;x=126616352;
#10;x=126716352;
#10;x=126816352;
#10;x=126916352;
#10;x=127016352;
#10;x=127116352;
#10;x=127216352;
#10;x=127316352;
#10;x=127416352;
#10;x=127516352;
#10;x=127616352;
#10;x=127716352;
#10;x=127816352;
#10;x=127916352;
#10;x=128016352;
#10;x=128116352;
#10;x=128216352;
#10;x=128316352;
#10;x=128416352;
#10;x=128516352;
#10;x=128616352;
#10;x=128716352;
#10;x=128816352;
#10;x=128916352;
#10;x=129016352;
#10;x=129116352;
#10;x=129216352;
#10;x=129316352;
#10;x=129416352;
#10;x=129516352;
#10;x=129616352;
#10;x=129716352;
#10;x=129816352;
#10;x=129916352;
#10;x=130016352;
#10;x=130116352;
#10;x=130216352;
#10;x=130316352;
#10;x=130416352;
#10;x=130516352;
#10;x=130616352;
#10;x=130716352;
#10;x=130816352;
#10;x=130916352;
#10;x=131016352;
#10;x=131116352;
#10;x=131216352;
#10;x=131316352;
#10;x=131416352;
#10;x=131516352;
#10;x=131616352;
#10;x=131716352;
#10;x=131816352;
#10;x=131916352;
#10;x=132016352;
#10;x=132116352;
#10;x=132216352;
#10;x=132316352;
#10;x=132416352;
#10;x=132516352;
#10;x=132616352;
#10;x=132716352;
#10;x=132816352;
#10;x=132916352;
#10;x=133016352;
#10;x=133116352;
#10;x=133216352;
#10;x=133316352;
#10;x=133416352;
#10;x=133516352;
#10;x=133616352;
#10;x=133716352;
#10;x=133816352;
#10;x=133916352;
#10;x=134016352;
#10;x=134116352;
#10;x=134216352;
#10;x=134316352;
#10;x=134416352;
#10;x=134516352;
#10;x=134616352;
#10;x=134716352;
#10;x=134816352;
#10;x=134916352;
#10;x=135016352;
#10;x=135116352;
#10;x=135216352;
#10;x=135316352;
#10;x=135416352;
#10;x=135516352;
#10;x=135616352;
#10;x=135716352;
#10;x=135816352;
#10;x=135916352;
#10;x=136016352;
#10;x=136116352;
#10;x=136216352;
#10;x=136316352;
#10;x=136416352;
#10;x=136516352;
#10;x=136616352;
#10;x=136716352;
#10;x=136816352;
#10;x=136916352;
#10;x=137016352;
#10;x=137116352;
#10;x=137216352;
#10;x=137316352;
#10;x=137416352;
#10;x=137516352;
#10;x=137616352;
#10;x=137716352;
#10;x=137816352;
#10;x=137916352;
#10;x=138016352;
#10;x=138116352;
#10;x=138216352;
#10;x=138316352;
#10;x=138416352;
#10;x=138516352;
#10;x=138616352;
#10;x=138716352;
#10;x=138816352;
#10;x=138916352;
#10;x=139016352;
#10;x=139116352;
#10;x=139216352;
#10;x=139316352;
#10;x=139416352;
#10;x=139516352;
#10;x=139616352;
#10;x=139716352;
#10;x=139816352;
#10;x=139916352;
#10;x=140016352;
#10;x=140116352;
#10;x=140216352;
#10;x=140316352;
#10;x=140416352;
#10;x=140516352;
#10;x=140616352;
#10;x=140716352;
#10;x=140816352;
#10;x=140916352;
#10;x=141016352;
#10;x=141116352;
#10;x=141216352;
#10;x=141316352;
#10;x=141416352;
#10;x=141516352;
#10;x=141616352;
#10;x=141716352;
#10;x=141816352;
#10;x=141916352;
#10;x=142016352;
#10;x=142116352;
#10;x=142216352;
#10;x=142316352;
#10;x=142416352;
#10;x=142516352;
#10;x=142616352;
#10;x=142716352;
#10;x=142816352;
#10;x=142916352;
#10;x=143016352;
#10;x=143116352;
#10;x=143216352;
#10;x=143316352;
#10;x=143416352;
#10;x=143516352;
#10;x=143616352;
#10;x=143716352;
#10;x=143816352;
#10;x=143916352;
#10;x=144016352;
#10;x=144116352;
#10;x=144216352;
#10;x=144316352;
#10;x=144416352;
#10;x=144516352;
#10;x=144616352;
#10;x=144716352;
#10;x=144816352;
#10;x=144916352;
#10;x=145016352;
#10;x=145116352;
#10;x=145216352;
#10;x=145316352;
#10;x=145416352;
#10;x=145516352;
#10;x=145616352;
#10;x=145716352;
#10;x=145816352;
#10;x=145916352;
#10;x=146016352;
#10;x=146116352;
#10;x=146216352;
#10;x=146316352;
#10;x=146416352;
#10;x=146516352;
#10;x=146616352;
#10;x=146716352;
#10;x=146816352;
#10;x=146916352;
#10;x=147016352;
#10;x=147116352;
#10;x=147216352;
#10;x=147316352;
#10;x=147416352;
#10;x=147516352;
#10;x=147616352;
#10;x=147716352;
#10;x=147816352;
#10;x=147916352;
#10;x=148016352;
#10;x=148116352;
#10;x=148216352;
#10;x=148316352;
#10;x=148416352;
#10;x=148516352;
#10;x=148616352;
#10;x=148716352;
#10;x=148816352;
#10;x=148916352;
#10;x=149016352;
#10;x=149116352;
#10;x=149216352;
#10;x=149316352;
#10;x=149416352;
#10;x=149516352;
#10;x=149616352;
#10;x=149716352;
#10;x=149816352;
#10;x=149916352;
#10;x=150016352;
#10;x=150116352;
#10;x=150216352;
#10;x=150316352;
#10;x=150416352;
#10;x=150516352;
#10;x=150616352;
#10;x=150716352;
#10;x=150816352;
#10;x=150916352;
#10;x=151016352;
#10;x=151116352;
#10;x=151216352;
#10;x=151316352;
#10;x=151416352;
#10;x=151516352;
#10;x=151616352;
#10;x=151716352;
#10;x=151816352;
#10;x=151916352;
#10;x=152016352;
#10;x=152116352;
#10;x=152216352;
#10;x=152316352;
#10;x=152416352;
#10;x=152516352;
#10;x=152616352;
#10;x=152716352;
#10;x=152816352;
#10;x=152916352;
#10;x=153016352;
#10;x=153116352;
#10;x=153216352;
#10;x=153316352;
#10;x=153416352;
#10;x=153516352;
#10;x=153616352;
#10;x=153716352;
#10;x=153816352;
#10;x=153916352;
#10;x=154016352;
#10;x=154116352;
#10;x=154216352;
#10;x=154316352;
#10;x=154416352;
#10;x=154516352;
#10;x=154616352;
#10;x=154716352;
#10;x=154816352;
#10;x=154916352;
#10;x=155016352;
#10;x=155116352;
#10;x=155216352;
#10;x=155316352;
#10;x=155416352;
#10;x=155516352;
#10;x=155616352;
#10;x=155716352;
#10;x=155816352;
#10;x=155916352;
#10;x=156016352;
#10;x=156116352;
#10;x=156216352;
#10;x=156316352;
#10;x=156416352;
#10;x=156516352;
#10;x=156616352;
#10;x=156716352;
#10;x=156816352;
#10;x=156916352;
#10;x=157016352;
#10;x=157116352;
#10;x=157216352;
#10;x=157316352;
#10;x=157416352;
#10;x=157516352;
#10;x=157616352;
#10;x=157716352;
#10;x=157816352;
#10;x=157916352;
#10;x=158016352;
#10;x=158116352;
#10;x=158216352;
#10;x=158316352;
#10;x=158416352;
#10;x=158516352;
#10;x=158616352;
#10;x=158716352;
#10;x=158816352;
#10;x=158916352;
#10;x=159016352;
#10;x=159116352;
#10;x=159216352;
#10;x=159316352;
#10;x=159416352;
#10;x=159516352;
#10;x=159616352;
#10;x=159716352;
#10;x=159816352;
#10;x=159916352;
#10;x=160016352;
#10;x=160116352;
#10;x=160216352;
#10;x=160316352;
#10;x=160416352;
#10;x=160516352;
#10;x=160616352;
#10;x=160716352;
#10;x=160816352;
#10;x=160916352;
#10;x=161016352;
#10;x=161116352;
#10;x=161216352;
#10;x=161316352;
#10;x=161416352;
#10;x=161516352;
#10;x=161616352;
#10;x=161716352;
#10;x=161816352;
#10;x=161916352;
#10;x=162016352;
#10;x=162116352;
#10;x=162216352;
#10;x=162316352;
#10;x=162416352;
#10;x=162516352;
#10;x=162616352;
#10;x=162716352;
#10;x=162816352;
#10;x=162916352;
#10;x=163016352;
#10;x=163116352;
#10;x=163216352;
#10;x=163316352;
#10;x=163416352;
#10;x=163516352;
#10;x=163616352;
#10;x=163716352;
#10;x=163816352;
#10;x=163916352;
#10;x=164016352;
#10;x=164116352;
#10;x=164216352;
#10;x=164316352;
#10;x=164416352;
#10;x=164516352;
#10;x=164616352;
#10;x=164716352;
#10;x=164816352;
#10;x=164916352;
#10;x=165016352;
#10;x=165116352;
#10;x=165216352;
#10;x=165316352;
#10;x=165416352;
#10;x=165516352;
#10;x=165616352;
#10;x=165716352;
#10;x=165816352;
#10;x=165916352;
#10;x=166016352;
#10;x=166116352;
#10;x=166216352;
#10;x=166316352;
#10;x=166416352;
#10;x=166516352;
#10;x=166616352;
#10;x=166716352;
#10;x=166816352;
#10;x=166916352;
#10;x=167016352;
#10;x=167116352;
#10;x=167216352;
#10;x=167316352;
#10;x=167416352;
#10;x=167516352;
#10;x=167616352;
#10;x=167716352;
#10;x=167816352;
#10;x=167916352;
#10;x=168016352;
#10;x=168116352;
#10;x=168216352;
#10;x=168316352;
#10;x=168416352;
#10;x=168516352;
#10;x=168616352;
#10;x=168716352;
#10;x=168816352;
#10;x=168916352;
#10;x=169016352;
#10;x=169116352;
#10;x=169216352;
#10;x=169316352;
#10;x=169416352;
#10;x=169516352;
#10;x=169616352;
#10;x=169716352;
#10;x=169816352;
#10;x=169916352;
#10;x=170016352;
#10;x=170116352;
#10;x=170216352;
#10;x=170316352;
#10;x=170416352;
#10;x=170516352;
#10;x=170616352;
#10;x=170716352;
#10;x=170816352;
#10;x=170916352;
#10;x=171016352;
#10;x=171116352;
#10;x=171216352;
#10;x=171316352;
#10;x=171416352;
#10;x=171516352;
#10;x=171616352;
#10;x=171716352;
#10;x=171816352;
#10;x=171916352;
#10;x=172016352;
#10;x=172116352;
#10;x=172216352;
#10;x=172316352;
#10;x=172416352;
#10;x=172516352;
#10;x=172616352;
#10;x=172716352;
#10;x=172816352;
#10;x=172916352;
#10;x=173016352;
#10;x=173116352;
#10;x=173216352;
#10;x=173316352;
#10;x=173416352;
#10;x=173516352;
#10;x=173616352;
#10;x=173716352;
#10;x=173816352;
#10;x=173916352;
#10;x=174016352;
#10;x=174116352;
#10;x=174216352;
#10;x=174316352;
#10;x=174416352;
#10;x=174516352;
#10;x=174616352;
#10;x=174716352;
#10;x=174816352;
#10;x=174916352;
#10;x=175016352;
#10;x=175116352;
#10;x=175216352;
#10;x=175316352;
#10;x=175416352;
#10;x=175516352;
#10;x=175616352;
#10;x=175716352;
#10;x=175816352;
#10;x=175916352;
#10;x=176016352;
#10;x=176116352;
#10;x=176216352;
#10;x=176316352;
#10;x=176416352;
#10;x=176516352;
#10;x=176616352;
#10;x=176716352;
#10;x=176816352;
#10;x=176916352;
#10;x=177016352;
#10;x=177116352;
#10;x=177216352;
#10;x=177316352;
#10;x=177416352;
#10;x=177516352;
#10;x=177616352;
#10;x=177716352;
#10;x=177816352;
#10;x=177916352;
#10;x=178016352;
#10;x=178116352;
#10;x=178216352;
#10;x=178316352;
#10;x=178416352;
#10;x=178516352;
#10;x=178616352;
#10;x=178716352;
#10;x=178816352;
#10;x=178916352;
#10;x=179016352;
#10;x=179116352;
#10;x=179216352;
#10;x=179316352;
#10;x=179416352;
#10;x=179516352;
#10;x=179616352;
#10;x=179716352;
#10;x=179816352;
#10;x=179916352;
#10;x=180016352;
#10;x=180116352;
#10;x=180216352;
#10;x=180316352;
#10;x=180416352;
#10;x=180516352;
#10;x=180616352;
#10;x=180716352;
#10;x=180816352;
#10;x=180916352;
#10;x=181016352;
#10;x=181116352;
#10;x=181216352;
#10;x=181316352;
#10;x=181416352;
#10;x=181516352;
#10;x=181616352;
#10;x=181716352;
#10;x=181816352;
#10;x=181916352;
#10;x=182016352;
#10;x=182116352;
#10;x=182216352;
#10;x=182316352;
#10;x=182416352;
#10;x=182516352;
#10;x=182616352;
#10;x=182716352;
#10;x=182816352;
#10;x=182916352;
#10;x=183016352;
#10;x=183116352;
#10;x=183216352;
#10;x=183316352;
#10;x=183416352;
#10;x=183516352;
#10;x=183616352;
#10;x=183716352;
#10;x=183816352;
#10;x=183916352;
#10;x=184016352;
#10;x=184116352;
#10;x=184216352;
#10;x=184316352;
#10;x=184416352;
#10;x=184516352;
#10;x=184616352;
#10;x=184716352;
#10;x=184816352;
#10;x=184916352;
#10;x=185016352;
#10;x=185116352;
#10;x=185216352;
#10;x=185316352;
#10;x=185416352;
#10;x=185516352;
#10;x=185616352;
#10;x=185716352;
#10;x=185816352;
#10;x=185916352;
#10;x=186016352;
#10;x=186116352;
#10;x=186216352;
#10;x=186316352;
#10;x=186416352;
#10;x=186516352;
#10;x=186616352;
#10;x=186716352;
#10;x=186816352;
#10;x=186916352;
#10;x=187016352;
#10;x=187116352;
#10;x=187216352;
#10;x=187316352;
#10;x=187416352;
#10;x=187516352;
#10;x=187616352;
#10;x=187716352;
#10;x=187816352;
#10;x=187916352;
#10;x=188016352;
#10;x=188116352;
#10;x=188216352;
#10;x=188316352;
#10;x=188416352;
#10;x=188516352;
#10;x=188616352;
#10;x=188716352;
#10;x=188816352;
#10;x=188916352;
#10;x=189016352;
#10;x=189116352;
#10;x=189216352;
#10;x=189316352;
#10;x=189416352;
#10;x=189516352;
#10;x=189616352;
#10;x=189716352;
#10;x=189816352;
#10;x=189916352;
#10;x=190016352;
#10;x=190116352;
#10;x=190216352;
#10;x=190316352;
#10;x=190416352;
#10;x=190516352;
#10;x=190616352;
#10;x=190716352;
#10;x=190816352;
#10;x=190916352;
#10;x=191016352;
#10;x=191116352;
#10;x=191216352;
#10;x=191316352;
#10;x=191416352;
#10;x=191516352;
#10;x=191616352;
#10;x=191716352;
#10;x=191816352;
#10;x=191916352;
#10;x=192016352;
#10;x=192116352;
#10;x=192216352;
#10;x=192316352;
#10;x=192416352;
#10;x=192516352;
#10;x=192616352;
#10;x=192716352;
#10;x=192816352;
#10;x=192916352;
#10;x=193016352;
#10;x=193116352;
#10;x=193216352;
#10;x=193316352;
#10;x=193416352;
#10;x=193516352;
#10;x=193616352;
#10;x=193716352;
#10;x=193816352;
#10;x=193916352;
#10;x=194016352;
#10;x=194116352;
#10;x=194216352;
#10;x=194316352;
#10;x=194416352;
#10;x=194516352;
#10;x=194616352;
#10;x=194716352;
#10;x=194816352;
#10;x=194916352;
#10;x=195016352;
#10;x=195116352;
#10;x=195216352;
#10;x=195316352;
#10;x=195416352;
#10;x=195516352;
#10;x=195616352;
#10;x=195716352;
#10;x=195816352;
#10;x=195916352;
#10;x=196016352;
#10;x=196116352;
#10;x=196216352;
#10;x=196316352;
#10;x=196416352;
#10;x=196516352;
#10;x=196616352;
#10;x=196716352;
#10;x=196816352;
#10;x=196916352;
#10;x=197016352;
#10;x=197116352;
#10;x=197216352;
#10;x=197316352;
#10;x=197416352;
#10;x=197516352;
#10;x=197616352;
#10;x=197716352;
#10;x=197816352;
#10;x=197916352;
#10;x=198016352;
#10;x=198116352;
#10;x=198216352;
#10;x=198316352;
#10;x=198416352;
#10;x=198516352;
#10;x=198616352;
#10;x=198716352;
#10;x=198816352;
#10;x=198916352;
#10;x=199016352;
#10;x=199116352;
#10;x=199216352;
#10;x=199316352;
#10;x=199416352;
#10;x=199516352;
#10;x=199616352;
#10;x=199716352;
#10;x=199816352;
#10;x=199916352;
#10;x=200016352;
#10;x=200116352;
#10;x=200216352;
#10;x=200316352;
#10;x=200416352;
#10;x=200516352;
#10;x=200616352;
#10;x=200716352;
#10;x=200816352;
#10;x=200916352;
#10;x=201016352;
#10;x=201116352;
#10;x=201216352;
#10;x=201316352;
#10;x=201416352;
#10;x=201516352;
#10;x=201616352;
#10;x=201716352;
#10;x=201816352;
#10;x=201916352;
#10;x=202016352;
#10;x=202116352;
#10;x=202216352;
#10;x=202316352;
#10;x=202416352;
#10;x=202516352;
#10;x=202616352;
#10;x=202716352;
#10;x=202816352;
#10;x=202916352;
#10;x=203016352;
#10;x=203116352;
#10;x=203216352;
#10;x=203316352;
#10;x=203416352;
#10;x=203516352;
#10;x=203616352;
#10;x=203716352;
#10;x=203816352;
#10;x=203916352;
#10;x=204016352;
#10;x=204116352;
#10;x=204216352;
#10;x=204316352;
#10;x=204416352;
#10;x=204516352;
#10;x=204616352;
#10;x=204716352;
#10;x=204816352;
#10;x=204916352;
#10;x=205016352;
#10;x=205116352;
#10;x=205216352;
#10;x=205316352;
#10;x=205416352;
#10;x=205516352;
#10;x=205616352;
#10;x=205716352;
#10;x=205816352;
#10;x=205916352;
#10;x=206016352;
#10;x=206116352;
#10;x=206216352;
#10;x=206316352;
#10;x=206416352;
#10;x=206516352;
#10;x=206616352;
#10;x=206716352;
#10;x=206816352;
#10;x=206916352;
#10;x=207016352;
#10;x=207116352;
#10;x=207216352;
#10;x=207316352;
#10;x=207416352;
#10;x=207516352;
#10;x=207616352;
#10;x=207716352;
#10;x=207816352;
#10;x=207916352;
#10;x=208016352;
#10;x=208116352;
#10;x=208216352;
#10;x=208316352;
#10;x=208416352;
#10;x=208516352;
#10;x=208616352;
#10;x=208716352;
#10;x=208816352;
#10;x=208916352;
#10;x=209016352;
#10;x=209116352;
#10;x=209216352;
#10;x=209316352;
#10;x=209416352;
#10;x=209516352;
#10;x=209616352;
#10;x=209716352;
#10;x=209816352;
#10;x=209916352;
#10;x=210016352;
#10;x=210116352;
#10;x=210216352;
#10;x=210316352;
#10;x=210416352;
#10;x=210516352;
#10;x=210616352;
#10;x=210716352;
#10;x=210816352;
#10;x=210916352;
#10;x=211016352;
#10;x=211116352;
#10;x=211216352;
#10;x=211316352;
#10;x=211416352;
#10;x=211516352;
#10;x=211616352;
#10;x=211716352;
#10;x=211816352;
#10;x=211916352;
#10;x=212016352;
#10;x=212116352;
#10;x=212216352;
#10;x=212316352;
#10;x=212416352;
#10;x=212516352;
#10;x=212616352;
#10;x=212716352;
#10;x=212816352;
#10;x=212916352;
#10;x=213016352;
#10;x=213116352;
#10;x=213216352;
#10;x=213316352;
#10;x=213416352;
#10;x=213516352;
#10;x=213616352;
#10;x=213716352;
#10;x=213816352;
#10;x=213916352;
#10;x=214016352;
#10;x=214116352;
#10;x=214216352;
#10;x=214316352;
#10;x=214416352;
#10;x=214516352;
#10;x=214616352;
#10;x=214716352;
#10;x=214816352;
#10;x=214916352;
#10;x=215016352;
#10;x=215116352;
#10;x=215216352;
#10;x=215316352;
#10;x=215416352;
#10;x=215516352;
#10;x=215616352;
#10;x=215716352;
#10;x=215816352;
#10;x=215916352;
#10;x=216016352;
#10;x=216116352;
#10;x=216216352;
#10;x=216316352;
#10;x=216416352;
#10;x=216516352;
#10;x=216616352;
#10;x=216716352;
#10;x=216816352;
#10;x=216916352;
#10;x=217016352;
#10;x=217116352;
#10;x=217216352;
#10;x=217316352;
#10;x=217416352;
#10;x=217516352;
#10;x=217616352;
#10;x=217716352;
#10;x=217816352;
#10;x=217916352;
#10;x=218016352;
#10;x=218116352;
#10;x=218216352;
#10;x=218316352;
#10;x=218416352;
#10;x=218516352;
#10;x=218616352;
#10;x=218716352;
#10;x=218816352;
#10;x=218916352;
#10;x=219016352;
#10;x=219116352;
#10;x=219216352;
#10;x=219316352;
#10;x=219416352;
#10;x=219516352;
#10;x=219616352;
#10;x=219716352;
#10;x=219816352;
#10;x=219916352;
#10;x=220016352;
#10;x=220116352;
#10;x=220216352;
#10;x=220316352;
#10;x=220416352;
#10;x=220516352;
#10;x=220616352;
#10;x=220716352;
#10;x=220816352;
#10;x=220916352;
#10;x=221016352;
#10;x=221116352;
#10;x=221216352;
#10;x=221316352;
#10;x=221416352;
#10;x=221516352;
#10;x=221616352;
#10;x=221716352;
#10;x=221816352;
#10;x=221916352;
#10;x=222016352;
#10;x=222116352;
#10;x=222216352;
#10;x=222316352;
#10;x=222416352;
#10;x=222516352;
#10;x=222616352;
#10;x=222716352;
#10;x=222816352;
#10;x=222916352;
#10;x=223016352;
#10;x=223116352;
#10;x=223216352;
#10;x=223316352;
#10;x=223416352;
#10;x=223516352;
#10;x=223616352;
#10;x=223716352;
#10;x=223816352;
#10;x=223916352;
#10;x=224016352;
#10;x=224116352;
#10;x=224216352;
#10;x=224316352;
#10;x=224416352;
#10;x=224516352;
#10;x=224616352;
#10;x=224716352;
#10;x=224816352;
#10;x=224916352;
#10;x=225016352;
#10;x=225116352;
#10;x=225216352;
#10;x=225316352;
#10;x=225416352;
#10;x=225516352;
#10;x=225616352;
#10;x=225716352;
#10;x=225816352;
#10;x=225916352;
#10;x=226016352;
#10;x=226116352;
#10;x=226216352;
#10;x=226316352;
#10;x=226416352;
#10;x=226516352;
#10;x=226616352;
#10;x=226716352;
#10;x=226816352;
#10;x=226916352;
#10;x=227016352;
#10;x=227116352;
#10;x=227216352;
#10;x=227316352;
#10;x=227416352;
#10;x=227516352;
#10;x=227616352;
#10;x=227716352;
#10;x=227816352;
#10;x=227916352;
#10;x=228016352;
#10;x=228116352;
#10;x=228216352;
#10;x=228316352;
#10;x=228416352;
#10;x=228516352;
#10;x=228616352;
#10;x=228716352;
#10;x=228816352;
#10;x=228916352;
#10;x=229016352;
#10;x=229116352;
#10;x=229216352;
#10;x=229316352;
#10;x=229416352;
#10;x=229516352;
#10;x=229616352;
#10;x=229716352;
#10;x=229816352;
#10;x=229916352;
#10;x=230016352;
#10;x=230116352;
#10;x=230216352;
#10;x=230316352;
#10;x=230416352;
#10;x=230516352;
#10;x=230616352;
#10;x=230716352;
#10;x=230816352;
#10;x=230916352;
#10;x=231016352;
#10;x=231116352;
#10;x=231216352;
#10;x=231316352;
#10;x=231416352;
#10;x=231516352;
#10;x=231616352;
#10;x=231716352;
#10;x=231816352;
#10;x=231916352;
#10;x=232016352;
#10;x=232116352;
#10;x=232216352;
#10;x=232316352;
#10;x=232416352;
#10;x=232516352;
#10;x=232616352;
#10;x=232716352;
#10;x=232816352;
#10;x=232916352;
#10;x=233016352;
#10;x=233116352;
#10;x=233216352;
#10;x=233316352;
#10;x=233416352;
#10;x=233516352;
#10;x=233616352;
#10;x=233716352;
#10;x=233816352;
#10;x=233916352;
#10;x=234016352;
#10;x=234116352;
#10;x=234216352;
#10;x=234316352;
#10;x=234416352;
#10;x=234516352;
#10;x=234616352;
#10;x=234716352;
#10;x=234816352;
#10;x=234916352;
#10;x=235016352;
#10;x=235116352;
#10;x=235216352;
#10;x=235316352;
#10;x=235416352;
#10;x=235516352;
#10;x=235616352;
#10;x=235716352;
#10;x=235816352;
#10;x=235916352;
#10;x=236016352;
#10;x=236116352;
#10;x=236216352;
#10;x=236316352;
#10;x=236416352;
#10;x=236516352;
#10;x=236616352;
#10;x=236716352;
#10;x=236816352;
#10;x=236916352;
#10;x=237016352;
#10;x=237116352;
#10;x=237216352;
#10;x=237316352;
#10;x=237416352;
#10;x=237516352;
#10;x=237616352;
#10;x=237716352;
#10;x=237816352;
#10;x=237916352;
#10;x=238016352;
#10;x=238116352;
#10;x=238216352;
#10;x=238316352;
#10;x=238416352;
#10;x=238516352;
#10;x=238616352;
#10;x=238716352;
#10;x=238816352;
#10;x=238916352;
#10;x=239016352;
#10;x=239116352;
#10;x=239216352;
#10;x=239316352;
#10;x=239416352;
#10;x=239516352;
#10;x=239616352;
#10;x=239716352;
#10;x=239816352;
#10;x=239916352;
#10;x=240016352;
#10;x=240116352;
#10;x=240216352;
#10;x=240316352;
#10;x=240416352;
#10;x=240516352;
#10;x=240616352;
#10;x=240716352;
#10;x=240816352;
#10;x=240916352;
#10;x=241016352;
#10;x=241116352;
#10;x=241216352;
#10;x=241316352;
#10;x=241416352;
#10;x=241516352;
#10;x=241616352;
#10;x=241716352;
#10;x=241816352;
#10;x=241916352;
#10;x=242016352;
#10;x=242116352;
#10;x=242216352;
#10;x=242316352;
#10;x=242416352;
#10;x=242516352;
#10;x=242616352;
#10;x=242716352;
#10;x=242816352;
#10;x=242916352;
#10;x=243016352;
#10;x=243116352;
#10;x=243216352;
#10;x=243316352;
#10;x=243416352;
#10;x=243516352;
#10;x=243616352;
#10;x=243716352;
#10;x=243816352;
#10;x=243916352;
#10;x=244016352;
#10;x=244116352;
#10;x=244216352;
#10;x=244316352;
#10;x=244416352;
#10;x=244516352;
#10;x=244616352;
#10;x=244716352;
#10;x=244816352;
#10;x=244916352;
#10;x=245016352;
#10;x=245116352;
#10;x=245216352;
#10;x=245316352;
#10;x=245416352;
#10;x=245516352;
#10;x=245616352;
#10;x=245716352;
#10;x=245816352;
#10;x=245916352;
#10;x=246016352;
#10;x=246116352;
#10;x=246216352;
#10;x=246316352;
#10;x=246416352;
#10;x=246516352;
#10;x=246616352;
#10;x=246716352;
#10;x=246816352;
#10;x=246916352;
#10;x=247016352;
#10;x=247116352;
#10;x=247216352;
#10;x=247316352;
#10;x=247416352;
#10;x=247516352;
#10;x=247616352;
#10;x=247716352;
#10;x=247816352;
#10;x=247916352;
#10;x=248016352;
#10;x=248116352;
#10;x=248216352;
#10;x=248316352;
#10;x=248416352;
#10;x=248516352;
#10;x=248616352;
#10;x=248716352;
#10;x=248816352;
#10;x=248916352;
#10;x=249016352;
#10;x=249116352;
#10;x=249216352;
#10;x=249316352;
#10;x=249416352;
#10;x=249516352;
#10;x=249616352;
#10;x=249716352;
#10;x=249816352;
#10;x=249916352;
#10;x=250016352;
#10;x=250116352;
#10;x=250216352;
#10;x=250316352;
#10;x=250416352;
#10;x=250516352;
#10;x=250616352;
#10;x=250716352;
#10;x=250816352;
#10;x=250916352;
#10;x=251016352;
#10;x=251116352;
#10;x=251216352;
#10;x=251316352;
#10;x=251416352;
#10;x=251516352;
#10;x=251616352;
#10;x=251716352;
#10;x=251816352;
#10;x=251916352;
#10;x=252016352;
#10;x=252116352;
#10;x=252216352;
#10;x=252316352;
#10;x=252416352;
#10;x=252516352;
#10;x=252616352;
#10;x=252716352;
#10;x=252816352;
#10;x=252916352;
#10;x=253016352;
#10;x=253116352;
#10;x=253216352;
#10;x=253316352;
#10;x=253416352;
#10;x=253516352;
#10;x=253616352;
#10;x=253716352;
#10;x=253816352;
#10;x=253916352;
#10;x=254016352;
#10;x=254116352;
#10;x=254216352;
#10;x=254316352;
#10;x=254416352;
#10;x=254516352;
#10;x=254616352;
#10;x=254716352;
#10;x=254816352;
#10;x=254916352;
#10;x=255016352;
#10;x=255116352;
#10;x=255216352;
#10;x=255316352;
#10;x=255416352;
#10;x=255516352;
#10;x=255616352;
#10;x=255716352;
#10;x=255816352;
#10;x=255916352;
#10;x=256016352;
#10;x=256116352;
#10;x=256216352;
#10;x=256316352;
#10;x=256416352;
#10;x=256516352;
#10;x=256616352;
#10;x=256716352;
#10;x=256816352;
#10;x=256916352;
#10;x=257016352;
#10;x=257116352;
#10;x=257216352;
#10;x=257316352;
#10;x=257416352;
#10;x=257516352;
#10;x=257616352;
#10;x=257716352;
#10;x=257816352;
#10;x=257916352;
#10;x=258016352;
#10;x=258116352;
#10;x=258216352;
#10;x=258316352;
#10;x=258416352;
#10;x=258516352;
#10;x=258616352;
#10;x=258716352;
#10;x=258816352;
#10;x=258916352;
#10;x=259016352;
#10;x=259116352;
#10;x=259216352;
#10;x=259316352;
#10;x=259416352;
#10;x=259516352;
#10;x=259616352;
#10;x=259716352;
#10;x=259816352;
#10;x=259916352;
#10;x=260016352;
#10;x=260116352;
#10;x=260216352;
#10;x=260316352;
#10;x=260416352;
#10;x=260516352;
#10;x=260616352;
#10;x=260716352;
#10;x=260816352;
#10;x=260916352;
#10;x=261016352;
#10;x=261116352;
#10;x=261216352;
#10;x=261316352;
#10;x=261416352;
#10;x=261516352;
#10;x=261616352;
#10;x=261716352;
#10;x=261816352;
#10;x=261916352;
#10;x=262016352;
#10;x=262116352;
#10;x=262216352;
#10;x=262316352;
#10;x=262416352;
#10;x=262516352;
#10;x=262616352;
#10;x=262716352;
#10;x=262816352;
#10;x=262916352;
#10;x=263016352;
#10;x=263116352;
#10;x=263216352;
#10;x=263316352;
#10;x=263416352;
#10;x=263516352;
#10;x=263616352;
#10;x=263716352;
#10;x=263816352;
#10;x=263916352;
#10;x=264016352;
#10;x=264116352;
#10;x=264216352;
#10;x=264316352;
#10;x=264416352;
#10;x=264516352;
#10;x=264616352;
#10;x=264716352;
#10;x=264816352;
#10;x=264916352;
#10;x=265016352;
#10;x=265116352;
#10;x=265216352;
#10;x=265316352;
#10;x=265416352;
#10;x=265516352;
#10;x=265616352;
#10;x=265716352;
#10;x=265816352;
#10;x=265916352;
#10;x=266016352;
#10;x=266116352;
#10;x=266216352;
#10;x=266316352;
#10;x=266416352;
#10;x=266516352;
#10;x=266616352;
#10;x=266716352;
#10;x=266816352;
#10;x=266916352;
#10;x=267016352;
#10;x=267116352;
#10;x=267216352;
#10;x=267316352;
#10;x=267416352;
#10;x=267516352;
#10;x=267616352;
#10;x=267716352;
#10;x=267816352;
#10;x=267916352;
#10;x=268016352;
#10;x=268116352;
#10;x=268216352;
#10;x=268316352;
#10;x=268416352;
#10;x=268516352;
#10;x=268616352;
#10;x=268716352;
#10;x=268816352;
#10;x=268916352;
#10;x=269016352;
#10;x=269116352;
#10;x=269216352;
#10;x=269316352;
#10;x=269416352;
#10;x=269516352;
#10;x=269616352;
#10;x=269716352;
#10;x=269816352;
#10;x=269916352;
#10;x=270016352;
#10;x=270116352;
#10;x=270216352;
#10;x=270316352;
#10;x=270416352;
#10;x=270516352;
#10;x=270616352;
#10;x=270716352;
#10;x=270816352;
#10;x=270916352;
#10;x=271016352;
#10;x=271116352;
#10;x=271216352;
#10;x=271316352;
#10;x=271416352;
#10;x=271516352;
#10;x=271616352;
#10;x=271716352;
#10;x=271816352;
#10;x=271916352;
#10;x=272016352;
#10;x=272116352;
#10;x=272216352;
#10;x=272316352;
#10;x=272416352;
#10;x=272516352;
#10;x=272616352;
#10;x=272716352;
#10;x=272816352;
#10;x=272916352;
#10;x=273016352;
#10;x=273116352;
#10;x=273216352;
#10;x=273316352;
#10;x=273416352;
#10;x=273516352;
#10;x=273616352;
#10;x=273716352;
#10;x=273816352;
#10;x=273916352;
#10;x=274016352;
#10;x=274116352;
#10;x=274216352;
#10;x=274316352;
#10;x=274416352;
#10;x=274516352;
#10;x=274616352;
#10;x=274716352;
#10;x=274816352;
#10;x=274916352;
#10;x=275016352;
#10;x=275116352;
#10;x=275216352;
#10;x=275316352;
#10;x=275416352;
#10;x=275516352;
#10;x=275616352;
#10;x=275716352;
#10;x=275816352;
#10;x=275916352;
#10;x=276016352;
#10;x=276116352;
#10;x=276216352;
#10;x=276316352;
#10;x=276416352;
#10;x=276516352;
#10;x=276616352;
#10;x=276716352;
#10;x=276816352;
#10;x=276916352;
#10;x=277016352;
#10;x=277116352;
#10;x=277216352;
#10;x=277316352;
#10;x=277416352;
#10;x=277516352;
#10;x=277616352;
#10;x=277716352;
#10;x=277816352;
#10;x=277916352;
#10;x=278016352;
#10;x=278116352;
#10;x=278216352;
#10;x=278316352;
#10;x=278416352;
#10;x=278516352;
#10;x=278616352;
#10;x=278716352;
#10;x=278816352;
#10;x=278916352;
#10;x=279016352;
#10;x=279116352;
#10;x=279216352;
#10;x=279316352;
#10;x=279416352;
#10;x=279516352;
#10;x=279616352;
#10;x=279716352;
#10;x=279816352;
#10;x=279916352;
#10;x=280016352;
#10;x=280116352;
#10;x=280216352;
#10;x=280316352;
#10;x=280416352;
#10;x=280516352;
#10;x=280616352;
#10;x=280716352;
#10;x=280816352;
#10;x=280916352;
#10;x=281016352;
#10;x=281116352;
#10;x=281216352;
#10;x=281316352;
#10;x=281416352;
#10;x=281516352;
#10;x=281616352;
#10;x=281716352;
#10;x=281816352;
#10;x=281916352;
#10;x=282016352;
#10;x=282116352;
#10;x=282216352;
#10;x=282316352;
#10;x=282416352;
#10;x=282516352;
#10;x=282616352;
#10;x=282716352;
#10;x=282816352;
#10;x=282916352;
#10;x=283016352;
#10;x=283116352;
#10;x=283216352;
#10;x=283316352;
#10;x=283416352;
#10;x=283516352;
#10;x=283616352;
#10;x=283716352;
#10;x=283816352;
#10;x=283916352;
#10;x=284016352;
#10;x=284116352;
#10;x=284216352;
#10;x=284316352;
#10;x=284416352;
#10;x=284516352;
#10;x=284616352;
#10;x=284716352;
#10;x=284816352;
#10;x=284916352;
#10;x=285016352;
#10;x=285116352;
#10;x=285216352;
#10;x=285316352;
#10;x=285416352;
#10;x=285516352;
#10;x=285616352;
#10;x=285716352;
#10;x=285816352;
#10;x=285916352;
#10;x=286016352;
#10;x=286116352;
#10;x=286216352;
#10;x=286316352;
#10;x=286416352;
#10;x=286516352;
#10;x=286616352;
#10;x=286716352;
#10;x=286816352;
#10;x=286916352;
#10;x=287016352;
#10;x=287116352;
#10;x=287216352;
#10;x=287316352;
#10;x=287416352;
#10;x=287516352;
#10;x=287616352;
#10;x=287716352;
#10;x=287816352;
#10;x=287916352;
#10;x=288016352;
#10;x=288116352;
#10;x=288216352;
#10;x=288316352;
#10;x=288416352;
#10;x=288516352;
#10;x=288616352;
#10;x=288716352;
#10;x=288816352;
#10;x=288916352;
#10;x=289016352;
#10;x=289116352;
#10;x=289216352;
#10;x=289316352;
#10;x=289416352;
#10;x=289516352;
#10;x=289616352;
#10;x=289716352;
#10;x=289816352;
#10;x=289916352;
#10;x=290016352;
#10;x=290116352;
#10;x=290216352;
#10;x=290316352;
#10;x=290416352;
#10;x=290516352;
#10;x=290616352;
#10;x=290716352;
#10;x=290816352;
#10;x=290916352;
#10;x=291016352;
#10;x=291116352;
#10;x=291216352;
#10;x=291316352;
#10;x=291416352;
#10;x=291516352;
#10;x=291616352;
#10;x=291716352;
#10;x=291816352;
#10;x=291916352;
#10;x=292016352;
#10;x=292116352;
#10;x=292216352;
#10;x=292316352;
#10;x=292416352;
#10;x=292516352;
#10;x=292616352;
#10;x=292716352;
#10;x=292816352;
#10;x=292916352;
#10;x=293016352;
#10;x=293116352;
#10;x=293216352;
#10;x=293316352;
#10;x=293416352;
#10;x=293516352;
#10;x=293616352;
#10;x=293716352;
#10;x=293816352;
#10;x=293916352;
#10;x=294016352;
#10;x=294116352;
#10;x=294216352;
#10;x=294316352;
#10;x=294416352;
#10;x=294516352;
#10;x=294616352;
#10;x=294716352;
#10;x=294816352;
#10;x=294916352;
#10;x=295016352;
#10;x=295116352;
#10;x=295216352;
#10;x=295316352;
#10;x=295416352;
#10;x=295516352;
#10;x=295616352;
#10;x=295716352;
#10;x=295816352;
#10;x=295916352;
#10;x=296016352;
#10;x=296116352;
#10;x=296216352;
#10;x=296316352;
#10;x=296416352;
#10;x=296516352;
#10;x=296616352;
#10;x=296716352;
#10;x=296816352;
#10;x=296916352;
#10;x=297016352;
#10;x=297116352;
#10;x=297216352;
#10;x=297316352;
#10;x=297416352;
#10;x=297516352;
#10;x=297616352;
#10;x=297716352;
#10;x=297816352;
#10;x=297916352;
#10;x=298016352;
#10;x=298116352;
#10;x=298216352;
#10;x=298316352;
#10;x=298416352;
#10;x=298516352;
#10;x=298616352;
#10;x=298716352;
#10;x=298816352;
#10;x=298916352;
#10;x=299016352;
#10;x=299116352;
#10;x=299216352;
#10;x=299316352;
#10;x=299416352;
#10;x=299516352;
#10;x=299616352;
#10;x=299716352;
#10;x=299816352;
#10;x=299916352;
#10;x=300016352;
#10;x=300116352;
#10;x=300216352;
#10;x=300316352;
#10;x=300416352;
#10;x=300516352;
#10;x=300616352;
#10;x=300716352;
#10;x=300816352;
#10;x=300916352;
#10;x=301016352;
#10;x=301116352;
#10;x=301216352;
#10;x=301316352;
#10;x=301416352;
#10;x=301516352;
#10;x=301616352;
#10;x=301716352;
#10;x=301816352;
#10;x=301916352;
#10;x=302016352;
#10;x=302116352;
#10;x=302216352;
#10;x=302316352;
#10;x=302416352;
#10;x=302516352;
#10;x=302616352;
#10;x=302716352;
#10;x=302816352;
#10;x=302916352;
#10;x=303016352;
#10;x=303116352;
#10;x=303216352;
#10;x=303316352;
#10;x=303416352;
#10;x=303516352;
#10;x=303616352;
#10;x=303716352;
#10;x=303816352;
#10;x=303916352;
#10;x=304016352;
#10;x=304116352;
#10;x=304216352;
#10;x=304316352;
#10;x=304416352;
#10;x=304516352;
#10;x=304616352;
#10;x=304716352;
#10;x=304816352;
#10;x=304916352;
#10;x=305016352;
#10;x=305116352;
#10;x=305216352;
#10;x=305316352;
#10;x=305416352;
#10;x=305516352;
#10;x=305616352;
#10;x=305716352;
#10;x=305816352;
#10;x=305916352;
#10;x=306016352;
#10;x=306116352;
#10;x=306216352;
#10;x=306316352;
#10;x=306416352;
#10;x=306516352;
#10;x=306616352;
#10;x=306716352;
#10;x=306816352;
#10;x=306916352;
#10;x=307016352;
#10;x=307116352;
#10;x=307216352;
#10;x=307316352;
#10;x=307416352;
#10;x=307516352;
#10;x=307616352;
#10;x=307716352;
#10;x=307816352;
#10;x=307916352;
#10;x=308016352;
#10;x=308116352;
#10;x=308216352;
#10;x=308316352;
#10;x=308416352;
#10;x=308516352;
#10;x=308616352;
#10;x=308716352;
#10;x=308816352;
#10;x=308916352;
#10;x=309016352;
#10;x=309116352;
#10;x=309216352;
#10;x=309316352;
#10;x=309416352;
#10;x=309516352;
#10;x=309616352;
#10;x=309716352;
#10;x=309816352;
#10;x=309916352;
#10;x=310016352;
#10;x=310116352;
#10;x=310216352;
#10;x=310316352;
#10;x=310416352;
#10;x=310516352;
#10;x=310616352;
#10;x=310716352;
#10;x=310816352;
#10;x=310916352;
#10;x=311016352;
#10;x=311116352;
#10;x=311216352;
#10;x=311316352;
#10;x=311416352;
#10;x=311516352;
#10;x=311616352;
#10;x=311716352;
#10;x=311816352;
#10;x=311916352;
#10;x=312016352;
#10;x=312116352;
#10;x=312216352;
#10;x=312316352;
#10;x=312416352;
#10;x=312516352;
#10;x=312616352;
#10;x=312716352;
#10;x=312816352;
#10;x=312916352;
#10;x=313016352;
#10;x=313116352;
#10;x=313216352;
#10;x=313316352;
#10;x=313416352;
#10;x=313516352;
#10;x=313616352;
#10;x=313716352;
#10;x=313816352;
#10;x=313916352;
#10;x=314016352;
#10;x=314116352;
#10;x=314216352;
#10;x=314316352;
#10;x=314416352;
#10;x=314516352;
#10;x=314616352;
#10;x=314716352;
#10;x=314816352;
#10;x=314916352;
#10;x=315016352;
#10;x=315116352;
#10;x=315216352;
#10;x=315316352;
#10;x=315416352;
#10;x=315516352;
#10;x=315616352;
#10;x=315716352;
#10;x=315816352;
#10;x=315916352;
#10;x=316016352;
#10;x=316116352;
#10;x=316216352;
#10;x=316316352;
#10;x=316416352;
#10;x=316516352;
#10;x=316616352;
#10;x=316716352;
#10;x=316816352;
#10;x=316916352;
#10;x=317016352;
#10;x=317116352;
#10;x=317216352;
#10;x=317316352;
#10;x=317416352;
#10;x=317516352;
#10;x=317616352;
#10;x=317716352;
#10;x=317816352;
#10;x=317916352;
#10;x=318016352;
#10;x=318116352;
#10;x=318216352;
#10;x=318316352;
#10;x=318416352;
#10;x=318516352;
#10;x=318616352;
#10;x=318716352;
#10;x=318816352;
#10;x=318916352;
#10;x=319016352;
#10;x=319116352;
#10;x=319216352;
#10;x=319316352;
#10;x=319416352;
#10;x=319516352;
#10;x=319616352;
#10;x=319716352;
#10;x=319816352;
#10;x=319916352;
#10;x=320016352;
#10;x=320116352;
#10;x=320216352;
#10;x=320316352;
#10;x=320416352;
#10;x=320516352;
#10;x=320616352;
#10;x=320716352;
#10;x=320816352;
#10;x=320916352;
#10;x=321016352;
#10;x=321116352;
#10;x=321216352;
#10;x=321316352;
#10;x=321416352;
#10;x=321516352;
#10;x=321616352;
#10;x=321716352;
#10;x=321816352;
#10;x=321916352;
#10;x=322016352;
#10;x=322116352;
#10;x=322216352;
#10;x=322316352;
#10;x=322416352;
#10;x=322516352;
#10;x=322616352;
#10;x=322716352;
#10;x=322816352;
#10;x=322916352;
#10;x=323016352;
#10;x=323116352;
#10;x=323216352;
#10;x=323316352;
#10;x=323416352;
#10;x=323516352;
#10;x=323616352;
#10;x=323716352;
#10;x=323816352;
#10;x=323916352;
#10;x=324016352;
#10;x=324116352;
#10;x=324216352;
#10;x=324316352;
#10;x=324416352;
#10;x=324516352;
#10;x=324616352;
#10;x=324716352;
#10;x=324816352;
#10;x=324916352;
#10;x=325016352;
#10;x=325116352;
#10;x=325216352;
#10;x=325316352;
#10;x=325416352;
#10;x=325516352;
#10;x=325616352;
#10;x=325716352;
#10;x=325816352;
#10;x=325916352;
#10;x=326016352;
#10;x=326116352;
#10;x=326216352;
#10;x=326316352;
#10;x=326416352;
#10;x=326516352;
#10;x=326616352;
#10;x=326716352;
#10;x=326816352;
#10;x=326916352;
#10;x=327016352;
#10;x=327116352;
#10;x=327216352;
#10;x=327316352;
#10;x=327416352;
#10;x=327516352;
#10;x=327616352;
#10;x=327716352;
#10;x=327816352;
#10;x=327916352;
#10;x=328016352;
#10;x=328116352;
#10;x=328216352;
#10;x=328316352;
#10;x=328416352;
#10;x=328516352;
#10;x=328616352;
#10;x=328716352;
#10;x=328816352;
#10;x=328916352;
#10;x=329016352;
#10;x=329116352;
#10;x=329216352;
#10;x=329316352;
#10;x=329416352;
#10;x=329516352;
#10;x=329616352;
#10;x=329716352;
#10;x=329816352;
#10;x=329916352;
#10;x=330016352;
#10;x=330116352;
#10;x=330216352;
#10;x=330316352;
#10;x=330416352;
#10;x=330516352;
#10;x=330616352;
#10;x=330716352;
#10;x=330816352;
#10;x=330916352;
#10;x=331016352;
#10;x=331116352;
#10;x=331216352;
#10;x=331316352;
#10;x=331416352;
#10;x=331516352;
#10;x=331616352;
#10;x=331716352;
#10;x=331816352;
#10;x=331916352;
#10;x=332016352;
#10;x=332116352;
#10;x=332216352;
#10;x=332316352;
#10;x=332416352;
#10;x=332516352;
#10;x=332616352;
#10;x=332716352;
#10;x=332816352;
#10;x=332916352;
#10;x=333016352;
#10;x=333116352;
#10;x=333216352;
#10;x=333316352;
#10;x=333416352;
#10;x=333516352;
#10;x=333616352;
#10;x=333716352;
#10;x=333816352;
#10;x=333916352;
#10;x=334016352;
#10;x=334116352;
#10;x=334216352;
#10;x=334316352;
#10;x=334416352;
#10;x=334516352;
#10;x=334616352;
#10;x=334716352;
#10;x=334816352;
#10;x=334916352;
#10;x=335016352;
#10;x=335116352;
#10;x=335216352;
#10;x=335316352;
#10;x=335416352;
#10;x=335516352;
#10;x=335616352;
#10;x=335716352;
#10;x=335816352;
#10;x=335916352;
#10;x=336016352;
#10;x=336116352;
#10;x=336216352;
#10;x=336316352;
#10;x=336416352;
#10;x=336516352;
#10;x=336616352;
#10;x=336716352;
#10;x=336816352;
#10;x=336916352;
#10;x=337016352;
#10;x=337116352;
#10;x=337216352;
#10;x=337316352;
#10;x=337416352;
#10;x=337516352;
#10;x=337616352;
#10;x=337716352;
#10;x=337816352;
#10;x=337916352;
#10;x=338016352;
#10;x=338116352;
#10;x=338216352;
#10;x=338316352;
#10;x=338416352;
#10;x=338516352;
#10;x=338616352;
#10;x=338716352;
#10;x=338816352;
#10;x=338916352;
#10;x=339016352;
#10;x=339116352;
#10;x=339216352;
#10;x=339316352;
#10;x=339416352;
#10;x=339516352;
#10;x=339616352;
#10;x=339716352;
#10;x=339816352;
#10;x=339916352;
#10;x=340016352;
#10;x=340116352;
#10;x=340216352;
#10;x=340316352;
#10;x=340416352;
#10;x=340516352;
#10;x=340616352;
#10;x=340716352;
#10;x=340816352;
#10;x=340916352;
#10;x=341016352;
#10;x=341116352;
#10;x=341216352;
#10;x=341316352;
#10;x=341416352;
#10;x=341516352;
#10;x=341616352;
#10;x=341716352;
#10;x=341816352;
#10;x=341916352;
#10;x=342016352;
#10;x=342116352;
#10;x=342216352;
#10;x=342316352;
#10;x=342416352;
#10;x=342516352;
#10;x=342616352;
#10;x=342716352;
#10;x=342816352;
#10;x=342916352;
#10;x=343016352;
#10;x=343116352;
#10;x=343216352;
#10;x=343316352;
#10;x=343416352;
#10;x=343516352;
#10;x=343616352;
#10;x=343716352;
#10;x=343816352;
#10;x=343916352;
#10;x=344016352;
#10;x=344116352;
#10;x=344216352;
#10;x=344316352;
#10;x=344416352;
#10;x=344516352;
#10;x=344616352;
#10;x=344716352;
#10;x=344816352;
#10;x=344916352;
#10;x=345016352;
#10;x=345116352;
#10;x=345216352;
#10;x=345316352;
#10;x=345416352;
#10;x=345516352;
#10;x=345616352;
#10;x=345716352;
#10;x=345816352;
#10;x=345916352;
#10;x=346016352;
#10;x=346116352;
#10;x=346216352;
#10;x=346316352;
#10;x=346416352;
#10;x=346516352;
#10;x=346616352;
#10;x=346716352;
#10;x=346816352;
#10;x=346916352;
#10;x=347016352;
#10;x=347116352;
#10;x=347216352;
#10;x=347316352;
#10;x=347416352;
#10;x=347516352;
#10;x=347616352;
#10;x=347716352;
#10;x=347816352;
#10;x=347916352;
#10;x=348016352;
#10;x=348116352;
#10;x=348216352;
#10;x=348316352;
#10;x=348416352;
#10;x=348516352;
#10;x=348616352;
#10;x=348716352;
#10;x=348816352;
#10;x=348916352;
#10;x=349016352;
#10;x=349116352;
#10;x=349216352;
#10;x=349316352;
#10;x=349416352;
#10;x=349516352;
#10;x=349616352;
#10;x=349716352;
#10;x=349816352;
#10;x=349916352;
#10;x=350016352;
#10;x=350116352;
#10;x=350216352;
#10;x=350316352;
#10;x=350416352;
#10;x=350516352;
#10;x=350616352;
#10;x=350716352;
#10;x=350816352;
#10;x=350916352;
#10;x=351016352;
#10;x=351116352;
#10;x=351216352;
#10;x=351316352;
#10;x=351416352;
#10;x=351516352;
#10;x=351616352;
#10;x=351716352;
#10;x=351816352;
#10;x=351916352;
#10;x=352016352;
#10;x=352116352;
#10;x=352216352;
#10;x=352316352;
#10;x=352416352;
#10;x=352516352;
#10;x=352616352;
#10;x=352716352;
#10;x=352816352;
#10;x=352916352;
#10;x=353016352;
#10;x=353116352;
#10;x=353216352;
#10;x=353316352;
#10;x=353416352;
#10;x=353516352;
#10;x=353616352;
#10;x=353716352;
#10;x=353816352;
#10;x=353916352;
#10;x=354016352;
#10;x=354116352;
#10;x=354216352;
#10;x=354316352;
#10;x=354416352;
#10;x=354516352;
#10;x=354616352;
#10;x=354716352;
#10;x=354816352;
#10;x=354916352;
#10;x=355016352;
#10;x=355116352;
#10;x=355216352;
#10;x=355316352;
#10;x=355416352;
#10;x=355516352;
#10;x=355616352;
#10;x=355716352;
#10;x=355816352;
#10;x=355916352;
#10;x=356016352;
#10;x=356116352;
#10;x=356216352;
#10;x=356316352;
#10;x=356416352;
#10;x=356516352;
#10;x=356616352;
#10;x=356716352;
#10;x=356816352;
#10;x=356916352;
#10;x=357016352;
#10;x=357116352;
#10;x=357216352;
#10;x=357316352;
#10;x=357416352;
#10;x=357516352;
#10;x=357616352;
#10;x=357716352;
#10;x=357816352;
#10;x=357916352;
#10;x=358016352;
#10;x=358116352;
#10;x=358216352;
#10;x=358316352;
#10;x=358416352;
#10;x=358516352;
#10;x=358616352;
#10;x=358716352;
#10;x=358816352;
#10;x=358916352;
#10;x=359016352;
#10;x=359116352;
#10;x=359216352;
#10;x=359316352;
#10;x=359416352;
#10;x=359516352;
#10;x=359616352;
#10;x=359716352;
#10;x=359816352;
#10;x=359916352;
#10;x=360016352;
#10;x=360116352;
#10;x=360216352;
#10;x=360316352;
#10;x=360416352;
#10;x=360516352;
#10;x=360616352;
#10;x=360716352;
#10;x=360816352;
#10;x=360916352;
#10;x=361016352;
#10;x=361116352;
#10;x=361216352;
#10;x=361316352;
#10;x=361416352;
#10;x=361516352;
#10;x=361616352;
#10;x=361716352;
#10;x=361816352;
#10;x=361916352;
#10;x=362016352;
#10;x=362116352;
#10;x=362216352;
#10;x=362316352;
#10;x=362416352;
#10;x=362516352;
#10;x=362616352;
#10;x=362716352;
#10;x=362816352;
#10;x=362916352;
#10;x=363016352;
#10;x=363116352;
#10;x=363216352;
#10;x=363316352;
#10;x=363416352;
#10;x=363516352;
#10;x=363616352;
#10;x=363716352;
#10;x=363816352;
#10;x=363916352;
#10;x=364016352;
#10;x=364116352;
#10;x=364216352;
#10;x=364316352;
#10;x=364416352;
#10;x=364516352;
#10;x=364616352;
#10;x=364716352;
#10;x=364816352;
#10;x=364916352;
#10;x=365016352;
#10;x=365116352;
#10;x=365216352;
#10;x=365316352;
#10;x=365416352;
#10;x=365516352;
#10;x=365616352;
#10;x=365716352;
#10;x=365816352;
#10;x=365916352;
#10;x=366016352;
#10;x=366116352;
#10;x=366216352;
#10;x=366316352;
#10;x=366416352;
#10;x=366516352;
#10;x=366616352;
#10;x=366716352;
#10;x=366816352;
#10;x=366916352;
#10;x=367016352;
#10;x=367116352;
#10;x=367216352;
#10;x=367316352;
#10;x=367416352;
#10;x=367516352;
#10;x=367616352;
#10;x=367716352;
#10;x=367816352;
#10;x=367916352;
#10;x=368016352;
#10;x=368116352;
#10;x=368216352;
#10;x=368316352;
#10;x=368416352;
#10;x=368516352;
#10;x=368616352;
#10;x=368716352;
#10;x=368816352;
#10;x=368916352;
#10;x=369016352;
#10;x=369116352;
#10;x=369216352;
#10;x=369316352;
#10;x=369416352;
#10;x=369516352;
#10;x=369616352;
#10;x=369716352;
#10;x=369816352;
#10;x=369916352;
#10;x=370016352;
#10;x=370116352;
#10;x=370216352;
#10;x=370316352;
#10;x=370416352;
#10;x=370516352;
#10;x=370616352;
#10;x=370716352;
#10;x=370816352;
#10;x=370916352;
#10;x=371016352;
#10;x=371116352;
#10;x=371216352;
#10;x=371316352;
#10;x=371416352;
#10;x=371516352;
#10;x=371616352;
#10;x=371716352;
#10;x=371816352;
#10;x=371916352;
#10;x=372016352;
#10;x=372116352;
#10;x=372216352;
#10;x=372316352;
#10;x=372416352;
#10;x=372516352;
#10;x=372616352;
#10;x=372716352;
#10;x=372816352;
#10;x=372916352;
#10;x=373016352;
#10;x=373116352;
#10;x=373216352;
#10;x=373316352;
#10;x=373416352;
#10;x=373516352;
#10;x=373616352;
#10;x=373716352;
#10;x=373816352;
#10;x=373916352;
#10;x=374016352;
#10;x=374116352;
#10;x=374216352;
#10;x=374316352;
#10;x=374416352;
#10;x=374516352;
#10;x=374616352;
#10;x=374716352;
#10;x=374816352;
#10;x=374916352;
#10;x=375016352;
#10;x=375116352;
#10;x=375216352;
#10;x=375316352;
#10;x=375416352;
#10;x=375516352;
#10;x=375616352;
#10;x=375716352;
#10;x=375816352;
#10;x=375916352;
#10;x=376016352;
#10;x=376116352;
#10;x=376216352;
#10;x=376316352;
#10;x=376416352;
#10;x=376516352;
#10;x=376616352;
#10;x=376716352;
#10;x=376816352;
#10;x=376916352;
#10;x=377016352;
#10;x=377116352;
#10;x=377216352;
#10;x=377316352;
#10;x=377416352;
#10;x=377516352;
#10;x=377616352;
#10;x=377716352;
#10;x=377816352;
#10;x=377916352;
#10;x=378016352;
#10;x=378116352;
#10;x=378216352;
#10;x=378316352;
#10;x=378416352;
#10;x=378516352;
#10;x=378616352;
#10;x=378716352;
#10;x=378816352;
#10;x=378916352;
#10;x=379016352;
#10;x=379116352;
#10;x=379216352;
#10;x=379316352;
#10;x=379416352;
#10;x=379516352;
#10;x=379616352;
#10;x=379716352;
#10;x=379816352;
#10;x=379916352;
#10;x=380016352;
#10;x=380116352;
#10;x=380216352;
#10;x=380316352;
#10;x=380416352;
#10;x=380516352;
#10;x=380616352;
#10;x=380716352;
#10;x=380816352;
#10;x=380916352;
#10;x=381016352;
#10;x=381116352;
#10;x=381216352;
#10;x=381316352;
#10;x=381416352;
#10;x=381516352;
#10;x=381616352;
#10;x=381716352;
#10;x=381816352;
#10;x=381916352;
#10;x=382016352;
#10;x=382116352;
#10;x=382216352;
#10;x=382316352;
#10;x=382416352;
#10;x=382516352;
#10;x=382616352;
#10;x=382716352;
#10;x=382816352;
#10;x=382916352;
#10;x=383016352;
#10;x=383116352;
#10;x=383216352;
#10;x=383316352;
#10;x=383416352;
#10;x=383516352;
#10;x=383616352;
#10;x=383716352;
#10;x=383816352;
#10;x=383916352;
#10;x=384016352;
#10;x=384116352;
#10;x=384216352;
#10;x=384316352;
#10;x=384416352;
#10;x=384516352;
#10;x=384616352;
#10;x=384716352;
#10;x=384816352;
#10;x=384916352;
#10;x=385016352;
#10;x=385116352;
#10;x=385216352;
#10;x=385316352;
#10;x=385416352;
#10;x=385516352;
#10;x=385616352;
#10;x=385716352;
#10;x=385816352;
#10;x=385916352;
#10;x=386016352;
#10;x=386116352;
#10;x=386216352;
#10;x=386316352;
#10;x=386416352;
#10;x=386516352;
#10;x=386616352;
#10;x=386716352;
#10;x=386816352;
#10;x=386916352;
#10;x=387016352;
#10;x=387116352;
#10;x=387216352;
#10;x=387316352;
#10;x=387416352;
#10;x=387516352;
#10;x=387616352;
#10;x=387716352;
#10;x=387816352;
#10;x=387916352;
#10;x=388016352;
#10;x=388116352;
#10;x=388216352;
#10;x=388316352;
#10;x=388416352;
#10;x=388516352;
#10;x=388616352;
#10;x=388716352;
#10;x=388816352;
#10;x=388916352;
#10;x=389016352;
#10;x=389116352;
#10;x=389216352;
#10;x=389316352;
#10;x=389416352;
#10;x=389516352;
#10;x=389616352;
#10;x=389716352;
#10;x=389816352;
#10;x=389916352;
#10;x=390016352;
#10;x=390116352;
#10;x=390216352;
#10;x=390316352;
#10;x=390416352;
#10;x=390516352;
#10;x=390616352;
#10;x=390716352;
#10;x=390816352;
#10;x=390916352;
#10;x=391016352;
#10;x=391116352;
#10;x=391216352;
#10;x=391316352;
#10;x=391416352;
#10;x=391516352;
#10;x=391616352;
#10;x=391716352;
#10;x=391816352;
#10;x=391916352;
#10;x=392016352;
#10;x=392116352;
#10;x=392216352;
#10;x=392316352;
#10;x=392416352;
#10;x=392516352;
#10;x=392616352;
#10;x=392716352;
#10;x=392816352;
#10;x=392916352;
#10;x=393016352;
#10;x=393116352;
#10;x=393216352;
#10;x=393316352;
#10;x=393416352;
#10;x=393516352;
#10;x=393616352;
#10;x=393716352;
#10;x=393816352;
#10;x=393916352;
#10;x=394016352;
#10;x=394116352;
#10;x=394216352;
#10;x=394316352;
#10;x=394416352;
#10;x=394516352;
#10;x=394616352;
#10;x=394716352;
#10;x=394816352;
#10;x=394916352;
#10;x=395016352;
#10;x=395116352;
#10;x=395216352;
#10;x=395316352;
#10;x=395416352;
#10;x=395516352;
#10;x=395616352;
#10;x=395716352;
#10;x=395816352;
#10;x=395916352;
#10;x=396016352;
#10;x=396116352;
#10;x=396216352;
#10;x=396316352;
#10;x=396416352;
#10;x=396516352;
#10;x=396616352;
#10;x=396716352;
#10;x=396816352;
#10;x=396916352;
#10;x=397016352;
#10;x=397116352;
#10;x=397216352;
#10;x=397316352;
#10;x=397416352;
#10;x=397516352;
#10;x=397616352;
#10;x=397716352;
#10;x=397816352;
#10;x=397916352;
#10;x=398016352;
#10;x=398116352;
#10;x=398216352;
#10;x=398316352;
#10;x=398416352;
#10;x=398516352;
#10;x=398616352;
#10;x=398716352;
#10;x=398816352;
#10;x=398916352;
#10;x=399016352;
#10;x=399116352;
#10;x=399216352;
#10;x=399316352;
#10;x=399416352;
#10;x=399516352;
#10;x=399616352;
#10;x=399716352;
#10;x=399816352;
#10;x=399916352;
#10;x=400016352;
#10;x=400116352;
#10;x=400216352;
#10;x=400316352;
#10;x=400416352;
#10;x=400516352;
#10;x=400616352;
#10;x=400716352;
#10;x=400816352;
#10;x=400916352;
#10;x=401016352;
#10;x=401116352;
#10;x=401216352;
#10;x=401316352;
#10;x=401416352;
#10;x=401516352;
#10;x=401616352;
#10;x=401716352;
#10;x=401816352;
#10;x=401916352;
#10;x=402016352;
#10;x=402116352;
#10;x=402216352;
#10;x=402316352;
#10;x=402416352;
#10;x=402516352;
#10;x=402616352;
#10;x=402716352;
#10;x=402816352;
#10;x=402916352;
#10;x=403016352;
#10;x=403116352;
#10;x=403216352;
#10;x=403316352;
#10;x=403416352;
#10;x=403516352;
#10;x=403616352;
#10;x=403716352;
#10;x=403816352;
#10;x=403916352;
#10;x=404016352;
#10;x=404116352;
#10;x=404216352;
#10;x=404316352;
#10;x=404416352;
#10;x=404516352;
#10;x=404616352;
#10;x=404716352;
#10;x=404816352;
#10;x=404916352;
#10;x=405016352;
#10;x=405116352;
#10;x=405216352;
#10;x=405316352;
#10;x=405416352;
#10;x=405516352;
#10;x=405616352;
#10;x=405716352;
#10;x=405816352;
#10;x=405916352;
#10;x=406016352;
#10;x=406116352;
#10;x=406216352;
#10;x=406316352;
#10;x=406416352;
#10;x=406516352;
#10;x=406616352;
#10;x=406716352;
#10;x=406816352;
#10;x=406916352;
#10;x=407016352;
#10;x=407116352;
#10;x=407216352;
#10;x=407316352;
#10;x=407416352;
#10;x=407516352;
#10;x=407616352;
#10;x=407716352;
#10;x=407816352;
#10;x=407916352;
#10;x=408016352;
#10;x=408116352;
#10;x=408216352;
#10;x=408316352;
#10;x=408416352;
#10;x=408516352;
#10;x=408616352;
#10;x=408716352;
#10;x=408816352;
#10;x=408916352;
#10;x=409016352;
#10;x=409116352;
#10;x=409216352;
#10;x=409316352;
#10;x=409416352;
#10;x=409516352;
#10;x=409616352;
#10;x=409716352;
#10;x=409816352;
#10;x=409916352;
#10;x=410016352;
#10;x=410116352;
#10;x=410216352;
#10;x=410316352;
#10;x=410416352;
#10;x=410516352;
#10;x=410616352;
#10;x=410716352;
#10;x=410816352;
#10;x=410916352;
#10;x=411016352;
#10;x=411116352;
#10;x=411216352;
#10;x=411316352;
#10;x=411416352;
#10;x=411516352;
#10;x=411616352;
#10;x=411716352;
#10;x=411816352;
#10;x=411916352;
#10;x=412016352;
#10;x=412116352;
#10;x=412216352;
#10;x=412316352;
#10;x=412416352;
#10;x=412516352;
#10;x=412616352;
#10;x=412716352;
#10;x=412816352;
#10;x=412916352;
#10;x=413016352;
#10;x=413116352;
#10;x=413216352;
#10;x=413316352;
#10;x=413416352;
#10;x=413516352;
#10;x=413616352;
#10;x=413716352;
#10;x=413816352;
#10;x=413916352;
#10;x=414016352;
#10;x=414116352;
#10;x=414216352;
#10;x=414316352;
#10;x=414416352;
#10;x=414516352;
#10;x=414616352;
#10;x=414716352;
#10;x=414816352;
#10;x=414916352;
#10;x=415016352;
#10;x=415116352;
#10;x=415216352;
#10;x=415316352;
#10;x=415416352;
#10;x=415516352;
#10;x=415616352;
#10;x=415716352;
#10;x=415816352;
#10;x=415916352;
#10;x=416016352;
#10;x=416116352;
#10;x=416216352;
#10;x=416316352;
#10;x=416416352;
#10;x=416516352;
#10;x=416616352;
#10;x=416716352;
#10;x=416816352;
#10;x=416916352;
#10;x=417016352;
#10;x=417116352;
#10;x=417216352;
#10;x=417316352;
#10;x=417416352;
#10;x=417516352;
#10;x=417616352;
#10;x=417716352;
#10;x=417816352;
#10;x=417916352;
#10;x=418016352;
#10;x=418116352;
#10;x=418216352;
#10;x=418316352;
#10;x=418416352;
#10;x=418516352;
#10;x=418616352;
#10;x=418716352;
#10;x=418816352;
#10;x=418916352;
#10;x=419016352;
#10;x=419116352;
#10;x=419216352;
#10;x=419316352;
#10;x=419416352;
#10;x=419516352;
#10;x=419616352;
#10;x=419716352;
#10;x=419816352;
#10;x=419916352;
#10;x=420016352;
#10;x=420116352;
#10;x=420216352;
#10;x=420316352;
#10;x=420416352;
#10;x=420516352;
#10;x=420616352;
#10;x=420716352;
#10;x=420816352;
#10;x=420916352;
#10;x=421016352;
#10;x=421116352;
#10;x=421216352;
#10;x=421316352;
#10;x=421416352;
#10;x=421516352;
#10;x=421616352;
#10;x=421716352;
#10;x=421816352;
#10;x=421916352;
#10;x=422016352;
#10;x=422116352;
#10;x=422216352;
#10;x=422316352;
#10;x=422416352;
#10;x=422516352;
#10;x=422616352;
#10;x=422716352;
#10;x=422816352;
#10;x=422916352;
#10;x=423016352;
#10;x=423116352;
#10;x=423216352;
#10;x=423316352;
#10;x=423416352;
#10;x=423516352;
#10;x=423616352;
#10;x=423716352;
#10;x=423816352;
#10;x=423916352;
#10;x=424016352;
#10;x=424116352;
#10;x=424216352;
#10;x=424316352;
#10;x=424416352;
#10;x=424516352;
#10;x=424616352;
#10;x=424716352;
#10;x=424816352;
#10;x=424916352;
#10;x=425016352;
#10;x=425116352;
#10;x=425216352;
#10;x=425316352;
#10;x=425416352;
#10;x=425516352;
#10;x=425616352;
#10;x=425716352;
#10;x=425816352;
#10;x=425916352;
#10;x=426016352;
#10;x=426116352;
#10;x=426216352;
#10;x=426316352;
#10;x=426416352;
#10;x=426516352;
#10;x=426616352;
#10;x=426716352;
#10;x=426816352;
#10;x=426916352;
#10;x=427016352;
#10;x=427116352;
#10;x=427216352;
#10;x=427316352;
#10;x=427416352;
#10;x=427516352;
#10;x=427616352;
#10;x=427716352;
#10;x=427816352;
#10;x=427916352;
#10;x=428016352;
#10;x=428116352;
#10;x=428216352;
#10;x=428316352;
#10;x=428416352;
#10;x=428516352;
#10;x=428616352;
#10;x=428716352;
#10;x=428816352;
#10;x=428916352;
#10;x=429016352;
#10;x=429116352;
#10;x=429216352;
#10;x=429316352;
#10;x=429416352;
#10;x=429516352;
#10;x=429616352;
#10;x=429716352;
#10;x=429816352;
#10;x=429916352;
#10;x=430016352;
#10;x=430116352;
#10;x=430216352;
#10;x=430316352;
#10;x=430416352;
#10;x=430516352;
#10;x=430616352;
#10;x=430716352;
#10;x=430816352;
#10;x=430916352;
#10;x=431016352;
#10;x=431116352;
#10;x=431216352;
#10;x=431316352;
#10;x=431416352;
#10;x=431516352;
#10;x=431616352;
#10;x=431716352;
#10;x=431816352;
#10;x=431916352;
#10;x=432016352;
#10;x=432116352;
#10;x=432216352;
#10;x=432316352;
#10;x=432416352;
#10;x=432516352;
#10;x=432616352;
#10;x=432716352;
#10;x=432816352;
#10;x=432916352;
#10;x=433016352;
#10;x=433116352;
#10;x=433216352;
#10;x=433316352;
#10;x=433416352;
#10;x=433516352;
#10;x=433616352;
#10;x=433716352;
#10;x=433816352;
#10;x=433916352;
#10;x=434016352;
#10;x=434116352;
#10;x=434216352;
#10;x=434316352;
#10;x=434416352;
#10;x=434516352;
#10;x=434616352;
#10;x=434716352;
#10;x=434816352;
#10;x=434916352;
#10;x=435016352;
#10;x=435116352;
#10;x=435216352;
#10;x=435316352;
#10;x=435416352;
#10;x=435516352;
#10;x=435616352;
#10;x=435716352;
#10;x=435816352;
#10;x=435916352;
#10;x=436016352;
#10;x=436116352;
#10;x=436216352;
#10;x=436316352;
#10;x=436416352;
#10;x=436516352;
#10;x=436616352;
#10;x=436716352;
#10;x=436816352;
#10;x=436916352;
#10;x=437016352;
#10;x=437116352;
#10;x=437216352;
#10;x=437316352;
#10;x=437416352;
#10;x=437516352;
#10;x=437616352;
#10;x=437716352;
#10;x=437816352;
#10;x=437916352;
#10;x=438016352;
#10;x=438116352;
#10;x=438216352;
#10;x=438316352;
#10;x=438416352;
#10;x=438516352;
#10;x=438616352;
#10;x=438716352;
#10;x=438816352;
#10;x=438916352;
#10;x=439016352;
#10;x=439116352;
#10;x=439216352;
#10;x=439316352;
#10;x=439416352;
#10;x=439516352;
#10;x=439616352;
#10;x=439716352;
#10;x=439816352;
#10;x=439916352;
#10;x=440016352;
#10;x=440116352;
#10;x=440216352;
#10;x=440316352;
#10;x=440416352;
#10;x=440516352;
#10;x=440616352;
#10;x=440716352;
#10;x=440816352;
#10;x=440916352;
#10;x=441016352;
#10;x=441116352;
#10;x=441216352;
#10;x=441316352;
#10;x=441416352;
#10;x=441516352;
#10;x=441616352;
#10;x=441716352;
#10;x=441816352;
#10;x=441916352;
#10;x=442016352;
#10;x=442116352;
#10;x=442216352;
#10;x=442316352;
#10;x=442416352;
#10;x=442516352;
#10;x=442616352;
#10;x=442716352;
#10;x=442816352;
#10;x=442916352;
#10;x=443016352;
#10;x=443116352;
#10;x=443216352;
#10;x=443316352;
#10;x=443416352;
#10;x=443516352;
#10;x=443616352;
#10;x=443716352;
#10;x=443816352;
#10;x=443916352;
#10;x=444016352;
#10;x=444116352;
#10;x=444216352;
#10;x=444316352;
#10;x=444416352;
#10;x=444516352;
#10;x=444616352;
#10;x=444716352;
#10;x=444816352;
#10;x=444916352;
#10;x=445016352;
#10;x=445116352;
#10;x=445216352;
#10;x=445316352;
#10;x=445416352;
#10;x=445516352;
#10;x=445616352;
#10;x=445716352;
#10;x=445816352;
#10;x=445916352;
#10;x=446016352;
#10;x=446116352;
#10;x=446216352;
#10;x=446316352;
#10;x=446416352;
#10;x=446516352;
#10;x=446616352;
#10;x=446716352;
#10;x=446816352;
#10;x=446916352;
#10;x=447016352;
#10;x=447116352;
#10;x=447216352;
#10;x=447316352;
#10;x=447416352;
#10;x=447516352;
#10;x=447616352;
#10;x=447716352;
#10;x=447816352;
#10;x=447916352;
#10;x=448016352;
#10;x=448116352;
#10;x=448216352;
#10;x=448316352;
#10;x=448416352;
#10;x=448516352;
#10;x=448616352;
#10;x=448716352;
#10;x=448816352;
#10;x=448916352;
#10;x=449016352;
#10;x=449116352;
#10;x=449216352;
#10;x=449316352;
#10;x=449416352;
#10;x=449516352;
#10;x=449616352;
#10;x=449716352;
#10;x=449816352;
#10;x=449916352;
#10;x=450016352;
#10;x=450116352;
#10;x=450216352;
#10;x=450316352;
#10;x=450416352;
#10;x=450516352;
#10;x=450616352;
#10;x=450716352;
#10;x=450816352;
#10;x=450916352;
#10;x=451016352;
#10;x=451116352;
#10;x=451216352;
#10;x=451316352;
#10;x=451416352;
#10;x=451516352;
#10;x=451616352;
#10;x=451716352;
#10;x=451816352;
#10;x=451916352;
#10;x=452016352;
#10;x=452116352;
#10;x=452216352;
#10;x=452316352;
#10;x=452416352;
#10;x=452516352;
#10;x=452616352;
#10;x=452716352;
#10;x=452816352;
#10;x=452916352;
#10;x=453016352;
#10;x=453116352;
#10;x=453216352;
#10;x=453316352;
#10;x=453416352;
#10;x=453516352;
#10;x=453616352;
#10;x=453716352;
#10;x=453816352;
#10;x=453916352;
#10;x=454016352;
#10;x=454116352;
#10;x=454216352;
#10;x=454316352;
#10;x=454416352;
#10;x=454516352;
#10;x=454616352;
#10;x=454716352;
#10;x=454816352;
#10;x=454916352;
#10;x=455016352;
#10;x=455116352;
#10;x=455216352;
#10;x=455316352;
#10;x=455416352;
#10;x=455516352;
#10;x=455616352;
#10;x=455716352;
#10;x=455816352;
#10;x=455916352;
#10;x=456016352;
#10;x=456116352;
#10;x=456216352;
#10;x=456316352;
#10;x=456416352;
#10;x=456516352;
#10;x=456616352;
#10;x=456716352;
#10;x=456816352;
#10;x=456916352;
#10;x=457016352;
#10;x=457116352;
#10;x=457216352;
#10;x=457316352;
#10;x=457416352;
#10;x=457516352;
#10;x=457616352;
#10;x=457716352;
#10;x=457816352;
#10;x=457916352;
#10;x=458016352;
#10;x=458116352;
#10;x=458216352;
#10;x=458316352;
#10;x=458416352;
#10;x=458516352;
#10;x=458616352;
#10;x=458716352;
#10;x=458816352;
#10;x=458916352;
#10;x=459016352;
#10;x=459116352;
#10;x=459216352;
#10;x=459316352;
#10;x=459416352;
#10;x=459516352;
#10;x=459616352;
#10;x=459716352;
#10;x=459816352;
#10;x=459916352;
#10;x=460016352;
#10;x=460116352;
#10;x=460216352;
#10;x=460316352;
#10;x=460416352;
#10;x=460516352;
#10;x=460616352;
#10;x=460716352;
#10;x=460816352;
#10;x=460916352;
#10;x=461016352;
#10;x=461116352;
#10;x=461216352;
#10;x=461316352;
#10;x=461416352;
#10;x=461516352;
#10;x=461616352;
#10;x=461716352;
#10;x=461816352;
#10;x=461916352;
#10;x=462016352;
#10;x=462116352;
#10;x=462216352;
#10;x=462316352;
#10;x=462416352;
#10;x=462516352;
#10;x=462616352;
#10;x=462716352;
#10;x=462816352;
#10;x=462916352;
#10;x=463016352;
#10;x=463116352;
#10;x=463216352;
#10;x=463316352;
#10;x=463416352;
#10;x=463516352;
#10;x=463616352;
#10;x=463716352;
#10;x=463816352;
#10;x=463916352;
#10;x=464016352;
#10;x=464116352;
#10;x=464216352;
#10;x=464316352;
#10;x=464416352;
#10;x=464516352;
#10;x=464616352;
#10;x=464716352;
#10;x=464816352;
#10;x=464916352;
#10;x=465016352;
#10;x=465116352;
#10;x=465216352;
#10;x=465316352;
#10;x=465416352;
#10;x=465516352;
#10;x=465616352;
#10;x=465716352;
#10;x=465816352;
#10;x=465916352;
#10;x=466016352;
#10;x=466116352;
#10;x=466216352;
#10;x=466316352;
#10;x=466416352;
#10;x=466516352;
#10;x=466616352;
#10;x=466716352;
#10;x=466816352;
#10;x=466916352;
#10;x=467016352;
#10;x=467116352;
#10;x=467216352;
#10;x=467316352;
#10;x=467416352;
#10;x=467516352;
#10;x=467616352;
#10;x=467716352;
#10;x=467816352;
#10;x=467916352;
#10;x=468016352;
#10;x=468116352;
#10;x=468216352;
#10;x=468316352;
#10;x=468416352;
#10;x=468516352;
#10;x=468616352;
#10;x=468716352;
#10;x=468816352;
#10;x=468916352;
#10;x=469016352;
#10;x=469116352;
#10;x=469216352;
#10;x=469316352;
#10;x=469416352;
#10;x=469516352;
#10;x=469616352;
#10;x=469716352;
#10;x=469816352;
#10;x=469916352;
#10;x=470016352;
#10;x=470116352;
#10;x=470216352;
#10;x=470316352;
#10;x=470416352;
#10;x=470516352;
#10;x=470616352;
#10;x=470716352;
#10;x=470816352;
#10;x=470916352;
#10;x=471016352;
#10;x=471116352;
#10;x=471216352;
#10;x=471316352;
#10;x=471416352;
#10;x=471516352;
#10;x=471616352;
#10;x=471716352;
#10;x=471816352;
#10;x=471916352;
#10;x=472016352;
#10;x=472116352;
#10;x=472216352;
#10;x=472316352;
#10;x=472416352;
#10;x=472516352;
#10;x=472616352;
#10;x=472716352;
#10;x=472816352;
#10;x=472916352;
#10;x=473016352;
#10;x=473116352;
#10;x=473216352;
#10;x=473316352;
#10;x=473416352;
#10;x=473516352;
#10;x=473616352;
#10;x=473716352;
#10;x=473816352;
#10;x=473916352;
#10;x=474016352;
#10;x=474116352;
#10;x=474216352;
#10;x=474316352;
#10;x=474416352;
#10;x=474516352;
#10;x=474616352;
#10;x=474716352;
#10;x=474816352;
#10;x=474916352;
#10;x=475016352;
#10;x=475116352;
#10;x=475216352;
#10;x=475316352;
#10;x=475416352;
#10;x=475516352;
#10;x=475616352;
#10;x=475716352;
#10;x=475816352;
#10;x=475916352;
#10;x=476016352;
#10;x=476116352;
#10;x=476216352;
#10;x=476316352;
#10;x=476416352;
#10;x=476516352;
#10;x=476616352;
#10;x=476716352;
#10;x=476816352;
#10;x=476916352;
#10;x=477016352;
#10;x=477116352;
#10;x=477216352;
#10;x=477316352;
#10;x=477416352;
#10;x=477516352;
#10;x=477616352;
#10;x=477716352;
#10;x=477816352;
#10;x=477916352;
#10;x=478016352;
#10;x=478116352;
#10;x=478216352;
#10;x=478316352;
#10;x=478416352;
#10;x=478516352;
#10;x=478616352;
#10;x=478716352;
#10;x=478816352;
#10;x=478916352;
#10;x=479016352;
#10;x=479116352;
#10;x=479216352;
#10;x=479316352;
#10;x=479416352;
#10;x=479516352;
#10;x=479616352;
#10;x=479716352;
#10;x=479816352;
#10;x=479916352;
#10;x=480016352;
#10;x=480116352;
#10;x=480216352;
#10;x=480316352;
#10;x=480416352;
#10;x=480516352;
#10;x=480616352;
#10;x=480716352;
#10;x=480816352;
#10;x=480916352;
#10;x=481016352;
#10;x=481116352;
#10;x=481216352;
#10;x=481316352;
#10;x=481416352;
#10;x=481516352;
#10;x=481616352;
#10;x=481716352;
#10;x=481816352;
#10;x=481916352;
#10;x=482016352;
#10;x=482116352;
#10;x=482216352;
#10;x=482316352;
#10;x=482416352;
#10;x=482516352;
#10;x=482616352;
#10;x=482716352;
#10;x=482816352;
#10;x=482916352;
#10;x=483016352;
#10;x=483116352;
#10;x=483216352;
#10;x=483316352;
#10;x=483416352;
#10;x=483516352;
#10;x=483616352;
#10;x=483716352;
#10;x=483816352;
#10;x=483916352;
#10;x=484016352;
#10;x=484116352;
#10;x=484216352;
#10;x=484316352;
#10;x=484416352;
#10;x=484516352;
#10;x=484616352;
#10;x=484716352;
#10;x=484816352;
#10;x=484916352;
#10;x=485016352;
#10;x=485116352;
#10;x=485216352;
#10;x=485316352;
#10;x=485416352;
#10;x=485516352;
#10;x=485616352;
#10;x=485716352;
#10;x=485816352;
#10;x=485916352;
#10;x=486016352;
#10;x=486116352;
#10;x=486216352;
#10;x=486316352;
#10;x=486416352;
#10;x=486516352;
#10;x=486616352;
#10;x=486716352;
#10;x=486816352;
#10;x=486916352;
#10;x=487016352;
#10;x=487116352;
#10;x=487216352;
#10;x=487316352;
#10;x=487416352;
#10;x=487516352;
#10;x=487616352;
#10;x=487716352;
#10;x=487816352;
#10;x=487916352;
#10;x=488016352;
#10;x=488116352;
#10;x=488216352;
#10;x=488316352;
#10;x=488416352;
#10;x=488516352;
#10;x=488616352;
#10;x=488716352;
#10;x=488816352;
#10;x=488916352;
#10;x=489016352;
#10;x=489116352;
#10;x=489216352;
#10;x=489316352;
#10;x=489416352;
#10;x=489516352;
#10;x=489616352;
#10;x=489716352;
#10;x=489816352;
#10;x=489916352;
#10;x=490016352;
#10;x=490116352;
#10;x=490216352;
#10;x=490316352;
#10;x=490416352;
#10;x=490516352;
#10;x=490616352;
#10;x=490716352;
#10;x=490816352;
#10;x=490916352;
#10;x=491016352;
#10;x=491116352;
#10;x=491216352;
#10;x=491316352;
#10;x=491416352;
#10;x=491516352;
#10;x=491616352;
#10;x=491716352;
#10;x=491816352;
#10;x=491916352;
#10;x=492016352;
#10;x=492116352;
#10;x=492216352;
#10;x=492316352;
#10;x=492416352;
#10;x=492516352;
#10;x=492616352;
#10;x=492716352;
#10;x=492816352;
#10;x=492916352;
#10;x=493016352;
#10;x=493116352;
#10;x=493216352;
#10;x=493316352;
#10;x=493416352;
#10;x=493516352;
#10;x=493616352;
#10;x=493716352;
#10;x=493816352;
#10;x=493916352;
#10;x=494016352;
#10;x=494116352;
#10;x=494216352;
#10;x=494316352;
#10;x=494416352;
#10;x=494516352;
#10;x=494616352;
#10;x=494716352;
#10;x=494816352;
#10;x=494916352;
#10;x=495016352;
#10;x=495116352;
#10;x=495216352;
#10;x=495316352;
#10;x=495416352;
#10;x=495516352;
#10;x=495616352;
#10;x=495716352;
#10;x=495816352;
#10;x=495916352;
#10;x=496016352;
#10;x=496116352;
#10;x=496216352;
#10;x=496316352;
#10;x=496416352;
#10;x=496516352;
#10;x=496616352;
#10;x=496716352;
#10;x=496816352;
#10;x=496916352;
#10;x=497016352;
#10;x=497116352;
#10;x=497216352;
#10;x=497316352;
#10;x=497416352;
#10;x=497516352;
#10;x=497616352;
#10;x=497716352;
#10;x=497816352;
#10;x=497916352;
#10;x=498016352;
#10;x=498116352;
#10;x=498216352;
#10;x=498316352;
#10;x=498416352;
#10;x=498516352;
#10;x=498616352;
#10;x=498716352;
#10;x=498816352;
#10;x=498916352;
#10;x=499016352;
#10;x=499116352;
#10;x=499216352;
#10;x=499316352;
#10;x=499416352;
#10;x=499516352;
#10;x=499616352;
#10;x=499716352;
#10;x=499816352;
#10;x=499916352;
#10;x=500016352;
#10;x=500116352;
#10;x=500216352;
#10;x=500316352;
#10;x=500416352;
#10;x=500516352;
#10;x=500616352;
#10;x=500716352;
#10;x=500816352;
#10;x=500916352;
#10;x=501016352;
#10;x=501116352;
#10;x=501216352;
#10;x=501316352;
#10;x=501416352;
#10;x=501516352;
#10;x=501616352;
#10;x=501716352;
#10;x=501816352;
#10;x=501916352;
#10;x=502016352;
#10;x=502116352;
#10;x=502216352;
#10;x=502316352;
#10;x=502416352;
#10;x=502516352;
#10;x=502616352;
#10;x=502716352;
#10;x=502816352;
#10;x=502916352;
#10;x=503016352;
#10;x=503116352;
#10;x=503216352;
#10;x=503316352;
#10;x=503416352;
#10;x=503516352;
#10;x=503616352;
#10;x=503716352;
#10;x=503816352;
#10;x=503916352;
#10;x=504016352;
#10;x=504116352;
#10;x=504216352;
#10;x=504316352;
#10;x=504416352;
#10;x=504516352;
#10;x=504616352;
#10;x=504716352;
#10;x=504816352;
#10;x=504916352;
#10;x=505016352;
#10;x=505116352;
#10;x=505216352;
#10;x=505316352;
#10;x=505416352;
#10;x=505516352;
#10;x=505616352;
#10;x=505716352;
#10;x=505816352;
#10;x=505916352;
#10;x=506016352;
#10;x=506116352;
#10;x=506216352;
#10;x=506316352;
#10;x=506416352;
#10;x=506516352;
#10;x=506616352;
#10;x=506716352;
#10;x=506816352;
#10;x=506916352;
#10;x=507016352;
#10;x=507116352;
#10;x=507216352;
#10;x=507316352;
#10;x=507416352;
#10;x=507516352;
#10;x=507616352;
#10;x=507716352;
#10;x=507816352;
#10;x=507916352;
#10;x=508016352;
#10;x=508116352;
#10;x=508216352;
#10;x=508316352;
#10;x=508416352;
#10;x=508516352;
#10;x=508616352;
#10;x=508716352;
#10;x=508816352;
#10;x=508916352;
#10;x=509016352;
#10;x=509116352;
#10;x=509216352;
#10;x=509316352;
#10;x=509416352;
#10;x=509516352;
#10;x=509616352;
#10;x=509716352;
#10;x=509816352;
#10;x=509916352;
#10;x=510016352;
#10;x=510116352;
#10;x=510216352;
#10;x=510316352;
#10;x=510416352;
#10;x=510516352;
#10;x=510616352;
#10;x=510716352;
#10;x=510816352;
#10;x=510916352;
#10;x=511016352;
#10;x=511116352;
#10;x=511216352;
#10;x=511316352;
#10;x=511416352;
#10;x=511516352;
#10;x=511616352;
#10;x=511716352;
#10;x=511816352;
#10;x=511916352;
#10;x=512016352;
#10;x=512116352;
#10;x=512216352;
#10;x=512316352;
#10;x=512416352;
#10;x=512516352;
#10;x=512616352;
#10;x=512716352;
#10;x=512816352;
#10;x=512916352;
#10;x=513016352;
#10;x=513116352;
#10;x=513216352;
#10;x=513316352;
#10;x=513416352;
#10;x=513516352;
#10;x=513616352;
#10;x=513716352;
#10;x=513816352;
#10;x=513916352;
#10;x=514016352;
#10;x=514116352;
#10;x=514216352;
#10;x=514316352;
#10;x=514416352;
#10;x=514516352;
#10;x=514616352;
#10;x=514716352;
#10;x=514816352;
#10;x=514916352;
#10;x=515016352;
#10;x=515116352;
#10;x=515216352;
#10;x=515316352;
#10;x=515416352;
#10;x=515516352;
#10;x=515616352;
#10;x=515716352;
#10;x=515816352;
#10;x=515916352;
#10;x=516016352;
#10;x=516116352;
#10;x=516216352;
#10;x=516316352;
#10;x=516416352;
#10;x=516516352;
#10;x=516616352;
#10;x=516716352;
#10;x=516816352;
#10;x=516916352;
#10;x=517016352;
#10;x=517116352;
#10;x=517216352;
#10;x=517316352;
#10;x=517416352;
#10;x=517516352;
#10;x=517616352;
#10;x=517716352;
#10;x=517816352;
#10;x=517916352;
#10;x=518016352;
#10;x=518116352;
#10;x=518216352;
#10;x=518316352;
#10;x=518416352;
#10;x=518516352;
#10;x=518616352;
#10;x=518716352;
#10;x=518816352;
#10;x=518916352;
#10;x=519016352;
#10;x=519116352;
#10;x=519216352;
#10;x=519316352;
#10;x=519416352;
#10;x=519516352;
#10;x=519616352;
#10;x=519716352;
#10;x=519816352;
#10;x=519916352;
#10;x=520016352;
#10;x=520116352;
#10;x=520216352;
#10;x=520316352;
#10;x=520416352;
#10;x=520516352;
#10;x=520616352;
#10;x=520716352;
#10;x=520816352;
#10;x=520916352;
#10;x=521016352;
#10;x=521116352;
#10;x=521216352;
#10;x=521316352;
#10;x=521416352;
#10;x=521516352;
#10;x=521616352;
#10;x=521716352;
#10;x=521816352;
#10;x=521916352;
#10;x=522016352;
#10;x=522116352;
#10;x=522216352;
#10;x=522316352;
#10;x=522416352;
#10;x=522516352;
#10;x=522616352;
#10;x=522716352;
#10;x=522816352;
#10;x=522916352;
#10;x=523016352;
#10;x=523116352;
#10;x=523216352;
#10;x=523316352;
#10;x=523416352;
#10;x=523516352;
#10;x=523616352;
#10;x=523716352;
#10;x=523816352;
#10;x=523916352;
#10;x=524016352;
#10;x=524116352;
#10;x=524216352;
#10;x=524316352;
#10;x=524416352;
#10;x=524516352;
#10;x=524616352;
#10;x=524716352;
#10;x=524816352;
#10;x=524916352;
#10;x=525016352;
#10;x=525116352;
#10;x=525216352;
#10;x=525316352;
#10;x=525416352;
#10;x=525516352;
#10;x=525616352;
#10;x=525716352;
#10;x=525816352;
#10;x=525916352;
#10;x=526016352;
#10;x=526116352;
#10;x=526216352;
#10;x=526316352;
#10;x=526416352;
#10;x=526516352;
#10;x=526616352;
#10;x=526716352;
#10;x=526816352;
#10;x=526916352;
#10;x=527016352;
#10;x=527116352;
#10;x=527216352;
#10;x=527316352;
#10;x=527416352;
#10;x=527516352;
#10;x=527616352;
#10;x=527716352;
#10;x=527816352;
#10;x=527916352;
#10;x=528016352;
#10;x=528116352;
#10;x=528216352;
#10;x=528316352;
#10;x=528416352;
#10;x=528516352;
#10;x=528616352;
#10;x=528716352;
#10;x=528816352;
#10;x=528916352;
#10;x=529016352;
#10;x=529116352;
#10;x=529216352;
#10;x=529316352;
#10;x=529416352;
#10;x=529516352;
#10;x=529616352;
#10;x=529716352;
#10;x=529816352;
#10;x=529916352;
#10;x=530016352;
#10;x=530116352;
#10;x=530216352;
#10;x=530316352;
#10;x=530416352;
#10;x=530516352;
#10;x=530616352;
#10;x=530716352;
#10;x=530816352;
#10;x=530916352;
#10;x=531016352;
#10;x=531116352;
#10;x=531216352;
#10;x=531316352;
#10;x=531416352;
#10;x=531516352;
#10;x=531616352;
#10;x=531716352;
#10;x=531816352;
#10;x=531916352;
#10;x=532016352;
#10;x=532116352;
#10;x=532216352;
#10;x=532316352;
#10;x=532416352;
#10;x=532516352;
#10;x=532616352;
#10;x=532716352;
#10;x=532816352;
#10;x=532916352;
#10;x=533016352;
#10;x=533116352;
#10;x=533216352;
#10;x=533316352;
#10;x=533416352;
#10;x=533516352;
#10;x=533616352;
#10;x=533716352;
#10;x=533816352;
#10;x=533916352;
#10;x=534016352;
#10;x=534116352;
#10;x=534216352;
#10;x=534316352;
#10;x=534416352;
#10;x=534516352;
#10;x=534616352;
#10;x=534716352;
#10;x=534816352;
#10;x=534916352;
#10;x=535016352;
#10;x=535116352;
#10;x=535216352;
#10;x=535316352;
#10;x=535416352;
#10;x=535516352;
#10;x=535616352;
#10;x=535716352;
#10;x=535816352;
#10;x=535916352;
#10;x=536016352;
#10;x=536116352;
#10;x=536216352;
#10;x=536316352;
#10;x=536416352;
#10;x=536516352;
#10;x=536616352;
#10;x=536716352;
#10;x=536816352;
#10;x=536916352;
#10;x=537016352;
#10;x=537116352;
#10;x=537216352;
#10;x=537316352;
#10;x=537416352;
#10;x=537516352;
#10;x=537616352;
#10;x=537716352;
#10;x=537816352;
#10;x=537916352;
#10;x=538016352;
#10;x=538116352;
#10;x=538216352;
#10;x=538316352;
#10;x=538416352;
#10;x=538516352;
#10;x=538616352;
#10;x=538716352;
#10;x=538816352;
#10;x=538916352;
#10;x=539016352;
#10;x=539116352;
#10;x=539216352;
#10;x=539316352;
#10;x=539416352;
#10;x=539516352;
#10;x=539616352;
#10;x=539716352;
#10;x=539816352;
#10;x=539916352;
#10;x=540016352;
#10;x=540116352;
#10;x=540216352;
#10;x=540316352;
#10;x=540416352;
#10;x=540516352;
#10;x=540616352;
#10;x=540716352;
#10;x=540816352;
#10;x=540916352;
#10;x=541016352;
#10;x=541116352;
#10;x=541216352;
#10;x=541316352;
#10;x=541416352;
#10;x=541516352;
#10;x=541616352;
#10;x=541716352;
#10;x=541816352;
#10;x=541916352;
#10;x=542016352;
#10;x=542116352;
#10;x=542216352;
#10;x=542316352;
#10;x=542416352;
#10;x=542516352;
#10;x=542616352;
#10;x=542716352;
#10;x=542816352;
#10;x=542916352;
#10;x=543016352;
#10;x=543116352;
#10;x=543216352;
#10;x=543316352;
#10;x=543416352;
#10;x=543516352;
#10;x=543616352;
#10;x=543716352;
#10;x=543816352;
#10;x=543916352;
#10;x=544016352;
#10;x=544116352;
#10;x=544216352;
#10;x=544316352;
#10;x=544416352;
#10;x=544516352;
#10;x=544616352;
#10;x=544716352;
#10;x=544816352;
#10;x=544916352;
#10;x=545016352;
#10;x=545116352;
#10;x=545216352;
#10;x=545316352;
#10;x=545416352;
#10;x=545516352;
#10;x=545616352;
#10;x=545716352;
#10;x=545816352;
#10;x=545916352;
#10;x=546016352;
#10;x=546116352;
#10;x=546216352;
#10;x=546316352;
#10;x=546416352;
#10;x=546516352;
#10;x=546616352;
#10;x=546716352;
#10;x=546816352;
#10;x=546916352;
#10;x=547016352;
#10;x=547116352;
#10;x=547216352;
#10;x=547316352;
#10;x=547416352;
#10;x=547516352;
#10;x=547616352;
#10;x=547716352;
#10;x=547816352;
#10;x=547916352;
#10;x=548016352;
#10;x=548116352;
#10;x=548216352;
#10;x=548316352;
#10;x=548416352;
#10;x=548516352;
#10;x=548616352;
#10;x=548716352;
#10;x=548816352;
#10;x=548916352;
#10;x=549016352;
#10;x=549116352;
#10;x=549216352;
#10;x=549316352;
#10;x=549416352;
#10;x=549516352;
#10;x=549616352;
#10;x=549716352;
#10;x=549816352;
#10;x=549916352;
#10;x=550016352;
#10;x=550116352;
#10;x=550216352;
#10;x=550316352;
#10;x=550416352;
#10;x=550516352;
#10;x=550616352;
#10;x=550716352;
#10;x=550816352;
#10;x=550916352;
#10;x=551016352;
#10;x=551116352;
#10;x=551216352;
#10;x=551316352;
#10;x=551416352;
#10;x=551516352;
#10;x=551616352;
#10;x=551716352;
#10;x=551816352;
#10;x=551916352;
#10;x=552016352;
#10;x=552116352;
#10;x=552216352;
#10;x=552316352;
#10;x=552416352;
#10;x=552516352;
#10;x=552616352;
#10;x=552716352;
#10;x=552816352;
#10;x=552916352;
#10;x=553016352;
#10;x=553116352;
#10;x=553216352;
#10;x=553316352;
#10;x=553416352;
#10;x=553516352;
#10;x=553616352;
#10;x=553716352;
#10;x=553816352;
#10;x=553916352;
#10;x=554016352;
#10;x=554116352;
#10;x=554216352;
#10;x=554316352;
#10;x=554416352;
#10;x=554516352;
#10;x=554616352;
#10;x=554716352;
#10;x=554816352;
#10;x=554916352;
#10;x=555016352;
#10;x=555116352;
#10;x=555216352;
#10;x=555316352;
#10;x=555416352;
#10;x=555516352;
#10;x=555616352;
#10;x=555716352;
#10;x=555816352;
#10;x=555916352;
#10;x=556016352;
#10;x=556116352;
#10;x=556216352;
#10;x=556316352;
#10;x=556416352;
#10;x=556516352;
#10;x=556616352;
#10;x=556716352;
#10;x=556816352;
#10;x=556916352;
#10;x=557016352;
#10;x=557116352;
#10;x=557216352;
#10;x=557316352;
#10;x=557416352;
#10;x=557516352;
#10;x=557616352;
#10;x=557716352;
#10;x=557816352;
#10;x=557916352;
#10;x=558016352;
#10;x=558116352;
#10;x=558216352;
#10;x=558316352;
#10;x=558416352;
#10;x=558516352;
#10;x=558616352;
#10;x=558716352;
#10;x=558816352;
#10;x=558916352;
#10;x=559016352;
#10;x=559116352;
#10;x=559216352;
#10;x=559316352;
#10;x=559416352;
#10;x=559516352;
#10;x=559616352;
#10;x=559716352;
#10;x=559816352;
#10;x=559916352;
#10;x=560016352;
#10;x=560116352;
#10;x=560216352;
#10;x=560316352;
#10;x=560416352;
#10;x=560516352;
#10;x=560616352;
#10;x=560716352;
#10;x=560816352;
#10;x=560916352;
#10;x=561016352;
#10;x=561116352;
#10;x=561216352;
#10;x=561316352;
#10;x=561416352;
#10;x=561516352;
#10;x=561616352;
#10;x=561716352;
#10;x=561816352;
#10;x=561916352;
#10;x=562016352;
#10;x=562116352;
#10;x=562216352;
#10;x=562316352;
#10;x=562416352;
#10;x=562516352;
#10;x=562616352;
#10;x=562716352;
#10;x=562816352;
#10;x=562916352;
#10;x=563016352;
#10;x=563116352;
#10;x=563216352;
#10;x=563316352;
#10;x=563416352;
#10;x=563516352;
#10;x=563616352;
#10;x=563716352;
#10;x=563816352;
#10;x=563916352;
#10;x=564016352;
#10;x=564116352;
#10;x=564216352;
#10;x=564316352;
#10;x=564416352;
#10;x=564516352;
#10;x=564616352;
#10;x=564716352;
#10;x=564816352;
#10;x=564916352;
#10;x=565016352;
#10;x=565116352;
#10;x=565216352;
#10;x=565316352;
#10;x=565416352;
#10;x=565516352;
#10;x=565616352;
#10;x=565716352;
#10;x=565816352;
#10;x=565916352;
#10;x=566016352;
#10;x=566116352;
#10;x=566216352;
#10;x=566316352;
#10;x=566416352;
#10;x=566516352;
#10;x=566616352;
#10;x=566716352;
#10;x=566816352;
#10;x=566916352;
#10;x=567016352;
#10;x=567116352;
#10;x=567216352;
#10;x=567316352;
#10;x=567416352;
#10;x=567516352;
#10;x=567616352;
#10;x=567716352;
#10;x=567816352;
#10;x=567916352;
#10;x=568016352;
#10;x=568116352;
#10;x=568216352;
#10;x=568316352;
#10;x=568416352;
#10;x=568516352;
#10;x=568616352;
#10;x=568716352;
#10;x=568816352;
#10;x=568916352;
#10;x=569016352;
#10;x=569116352;
#10;x=569216352;
#10;x=569316352;
#10;x=569416352;
#10;x=569516352;
#10;x=569616352;
#10;x=569716352;
#10;x=569816352;
#10;x=569916352;
#10;x=570016352;
#10;x=570116352;
#10;x=570216352;
#10;x=570316352;
#10;x=570416352;
#10;x=570516352;
#10;x=570616352;
#10;x=570716352;
#10;x=570816352;
#10;x=570916352;
#10;x=571016352;
#10;x=571116352;
#10;x=571216352;
#10;x=571316352;
#10;x=571416352;
#10;x=571516352;
#10;x=571616352;
#10;x=571716352;
#10;x=571816352;
#10;x=571916352;
#10;x=572016352;
#10;x=572116352;
#10;x=572216352;
#10;x=572316352;
#10;x=572416352;
#10;x=572516352;
#10;x=572616352;
#10;x=572716352;
#10;x=572816352;
#10;x=572916352;
#10;x=573016352;
#10;x=573116352;
#10;x=573216352;
#10;x=573316352;
#10;x=573416352;
#10;x=573516352;
#10;x=573616352;
#10;x=573716352;
#10;x=573816352;
#10;x=573916352;
#10;x=574016352;
#10;x=574116352;
#10;x=574216352;
#10;x=574316352;
#10;x=574416352;
#10;x=574516352;
#10;x=574616352;
#10;x=574716352;
#10;x=574816352;
#10;x=574916352;
#10;x=575016352;
#10;x=575116352;
#10;x=575216352;
#10;x=575316352;
#10;x=575416352;
#10;x=575516352;
#10;x=575616352;
#10;x=575716352;
#10;x=575816352;
#10;x=575916352;
#10;x=576016352;
#10;x=576116352;
#10;x=576216352;
#10;x=576316352;
#10;x=576416352;
#10;x=576516352;
#10;x=576616352;
#10;x=576716352;
#10;x=576816352;
#10;x=576916352;
#10;x=577016352;
#10;x=577116352;
#10;x=577216352;
#10;x=577316352;
#10;x=577416352;
#10;x=577516352;
#10;x=577616352;
#10;x=577716352;
#10;x=577816352;
#10;x=577916352;
#10;x=578016352;
#10;x=578116352;
#10;x=578216352;
#10;x=578316352;
#10;x=578416352;
#10;x=578516352;
#10;x=578616352;
#10;x=578716352;
#10;x=578816352;
#10;x=578916352;
#10;x=579016352;
#10;x=579116352;
#10;x=579216352;
#10;x=579316352;
#10;x=579416352;
#10;x=579516352;
#10;x=579616352;
#10;x=579716352;
#10;x=579816352;
#10;x=579916352;
#10;x=580016352;
#10;x=580116352;
#10;x=580216352;
#10;x=580316352;
#10;x=580416352;
#10;x=580516352;
#10;x=580616352;
#10;x=580716352;
#10;x=580816352;
#10;x=580916352;
#10;x=581016352;
#10;x=581116352;
#10;x=581216352;
#10;x=581316352;
#10;x=581416352;
#10;x=581516352;
#10;x=581616352;
#10;x=581716352;
#10;x=581816352;
#10;x=581916352;
#10;x=582016352;
#10;x=582116352;
#10;x=582216352;
#10;x=582316352;
#10;x=582416352;
#10;x=582516352;
#10;x=582616352;
#10;x=582716352;
#10;x=582816352;
#10;x=582916352;
#10;x=583016352;
#10;x=583116352;
#10;x=583216352;
#10;x=583316352;
#10;x=583416352;
#10;x=583516352;
#10;x=583616352;
#10;x=583716352;
#10;x=583816352;
#10;x=583916352;
#10;x=584016352;
#10;x=584116352;
#10;x=584216352;
#10;x=584316352;
#10;x=584416352;
#10;x=584516352;
#10;x=584616352;
#10;x=584716352;
#10;x=584816352;
#10;x=584916352;
#10;x=585016352;
#10;x=585116352;
#10;x=585216352;
#10;x=585316352;
#10;x=585416352;
#10;x=585516352;
#10;x=585616352;
#10;x=585716352;
#10;x=585816352;
#10;x=585916352;
#10;x=586016352;
#10;x=586116352;
#10;x=586216352;
#10;x=586316352;
#10;x=586416352;
#10;x=586516352;
#10;x=586616352;
#10;x=586716352;
#10;x=586816352;
#10;x=586916352;
#10;x=587016352;
#10;x=587116352;
#10;x=587216352;
#10;x=587316352;
#10;x=587416352;
#10;x=587516352;
#10;x=587616352;
#10;x=587716352;
#10;x=587816352;
#10;x=587916352;
#10;x=588016352;
#10;x=588116352;
#10;x=588216352;
#10;x=588316352;
#10;x=588416352;
#10;x=588516352;
#10;x=588616352;
#10;x=588716352;
#10;x=588816352;
#10;x=588916352;
#10;x=589016352;
#10;x=589116352;
#10;x=589216352;
#10;x=589316352;
#10;x=589416352;
#10;x=589516352;
#10;x=589616352;
#10;x=589716352;
#10;x=589816352;
#10;x=589916352;
#10;x=590016352;
#10;x=590116352;
#10;x=590216352;
#10;x=590316352;
#10;x=590416352;
#10;x=590516352;
#10;x=590616352;
#10;x=590716352;
#10;x=590816352;
#10;x=590916352;
#10;x=591016352;
#10;x=591116352;
#10;x=591216352;
#10;x=591316352;
#10;x=591416352;
#10;x=591516352;
#10;x=591616352;
#10;x=591716352;
#10;x=591816352;
#10;x=591916352;
#10;x=592016352;
#10;x=592116352;
#10;x=592216352;
#10;x=592316352;
#10;x=592416352;
#10;x=592516352;
#10;x=592616352;
#10;x=592716352;
#10;x=592816352;
#10;x=592916352;
#10;x=593016352;
#10;x=593116352;
#10;x=593216352;
#10;x=593316352;
#10;x=593416352;
#10;x=593516352;
#10;x=593616352;
#10;x=593716352;
#10;x=593816352;
#10;x=593916352;
#10;x=594016352;
#10;x=594116352;
#10;x=594216352;
#10;x=594316352;
#10;x=594416352;
#10;x=594516352;
#10;x=594616352;
#10;x=594716352;
#10;x=594816352;
#10;x=594916352;
#10;x=595016352;
#10;x=595116352;
#10;x=595216352;
#10;x=595316352;
#10;x=595416352;
#10;x=595516352;
#10;x=595616352;
#10;x=595716352;
#10;x=595816352;
#10;x=595916352;
#10;x=596016352;
#10;x=596116352;
#10;x=596216352;
#10;x=596316352;
#10;x=596416352;
#10;x=596516352;
#10;x=596616352;
#10;x=596716352;
#10;x=596816352;
#10;x=596916352;
#10;x=597016352;
#10;x=597116352;
#10;x=597216352;
#10;x=597316352;
#10;x=597416352;
#10;x=597516352;
#10;x=597616352;
#10;x=597716352;
#10;x=597816352;
#10;x=597916352;
#10;x=598016352;
#10;x=598116352;
#10;x=598216352;
#10;x=598316352;
#10;x=598416352;
#10;x=598516352;
#10;x=598616352;
#10;x=598716352;
#10;x=598816352;
#10;x=598916352;
#10;x=599016352;
#10;x=599116352;
#10;x=599216352;
#10;x=599316352;
#10;x=599416352;
#10;x=599516352;
#10;x=599616352;
#10;x=599716352;
#10;x=599816352;
#10;x=599916352;
#10;x=600016352;
#10;x=600116352;
#10;x=600216352;
#10;x=600316352;
#10;x=600416352;
#10;x=600516352;
#10;x=600616352;
#10;x=600716352;
#10;x=600816352;
#10;x=600916352;
#10;x=601016352;
#10;x=601116352;
#10;x=601216352;
#10;x=601316352;
#10;x=601416352;
#10;x=601516352;
#10;x=601616352;
#10;x=601716352;
#10;x=601816352;
#10;x=601916352;
#10;x=602016352;
#10;x=602116352;
#10;x=602216352;
#10;x=602316352;
#10;x=602416352;
#10;x=602516352;
#10;x=602616352;
#10;x=602716352;
#10;x=602816352;
#10;x=602916352;
#10;x=603016352;
#10;x=603116352;
#10;x=603216352;
#10;x=603316352;
#10;x=603416352;
#10;x=603516352;
#10;x=603616352;
#10;x=603716352;
#10;x=603816352;
#10;x=603916352;
#10;x=604016352;
#10;x=604116352;
#10;x=604216352;
#10;x=604316352;
#10;x=604416352;
#10;x=604516352;
#10;x=604616352;
#10;x=604716352;
#10;x=604816352;
#10;x=604916352;
#10;x=605016352;
#10;x=605116352;
#10;x=605216352;
#10;x=605316352;
#10;x=605416352;
#10;x=605516352;
#10;x=605616352;
#10;x=605716352;
#10;x=605816352;
#10;x=605916352;
#10;x=606016352;
#10;x=606116352;
#10;x=606216352;
#10;x=606316352;
#10;x=606416352;
#10;x=606516352;
#10;x=606616352;
#10;x=606716352;
#10;x=606816352;
#10;x=606916352;
#10;x=607016352;
#10;x=607116352;
#10;x=607216352;
#10;x=607316352;
#10;x=607416352;
#10;x=607516352;
#10;x=607616352;
#10;x=607716352;
#10;x=607816352;
#10;x=607916352;
#10;x=608016352;
#10;x=608116352;
#10;x=608216352;
#10;x=608316352;
#10;x=608416352;
#10;x=608516352;
#10;x=608616352;
#10;x=608716352;
#10;x=608816352;
#10;x=608916352;
#10;x=609016352;
#10;x=609116352;
#10;x=609216352;
#10;x=609316352;
#10;x=609416352;
#10;x=609516352;
#10;x=609616352;
#10;x=609716352;
#10;x=609816352;
#10;x=609916352;
#10;x=610016352;
#10;x=610116352;
#10;x=610216352;
#10;x=610316352;
#10;x=610416352;
#10;x=610516352;
#10;x=610616352;
#10;x=610716352;
#10;x=610816352;
#10;x=610916352;
#10;x=611016352;
#10;x=611116352;
#10;x=611216352;
#10;x=611316352;
#10;x=611416352;
#10;x=611516352;
#10;x=611616352;
#10;x=611716352;
#10;x=611816352;
#10;x=611916352;
#10;x=612016352;
#10;x=612116352;
#10;x=612216352;
#10;x=612316352;
#10;x=612416352;
#10;x=612516352;
#10;x=612616352;
#10;x=612716352;
#10;x=612816352;
#10;x=612916352;
#10;x=613016352;
#10;x=613116352;
#10;x=613216352;
#10;x=613316352;
#10;x=613416352;
#10;x=613516352;
#10;x=613616352;
#10;x=613716352;
#10;x=613816352;
#10;x=613916352;
#10;x=614016352;
#10;x=614116352;
#10;x=614216352;
#10;x=614316352;
#10;x=614416352;
#10;x=614516352;
#10;x=614616352;
#10;x=614716352;
#10;x=614816352;
#10;x=614916352;
#10;x=615016352;
#10;x=615116352;
#10;x=615216352;
#10;x=615316352;
#10;x=615416352;
#10;x=615516352;
#10;x=615616352;
#10;x=615716352;
#10;x=615816352;
#10;x=615916352;
#10;x=616016352;
#10;x=616116352;
#10;x=616216352;
#10;x=616316352;
#10;x=616416352;
#10;x=616516352;
#10;x=616616352;
#10;x=616716352;
#10;x=616816352;
#10;x=616916352;
#10;x=617016352;
#10;x=617116352;
#10;x=617216352;
#10;x=617316352;
#10;x=617416352;
#10;x=617516352;
#10;x=617616352;
#10;x=617716352;
#10;x=617816352;
#10;x=617916352;
#10;x=618016352;
#10;x=618116352;
#10;x=618216352;
#10;x=618316352;
#10;x=618416352;
#10;x=618516352;
#10;x=618616352;
#10;x=618716352;
#10;x=618816352;
#10;x=618916352;
#10;x=619016352;
#10;x=619116352;
#10;x=619216352;
#10;x=619316352;
#10;x=619416352;
#10;x=619516352;
#10;x=619616352;
#10;x=619716352;
#10;x=619816352;
#10;x=619916352;
#10;x=620016352;
#10;x=620116352;
#10;x=620216352;
#10;x=620316352;
#10;x=620416352;
#10;x=620516352;
#10;x=620616352;
#10;x=620716352;
#10;x=620816352;
#10;x=620916352;
#10;x=621016352;
#10;x=621116352;
#10;x=621216352;
#10;x=621316352;
#10;x=621416352;
#10;x=621516352;
#10;x=621616352;
#10;x=621716352;
#10;x=621816352;
#10;x=621916352;
#10;x=622016352;
#10;x=622116352;
#10;x=622216352;
#10;x=622316352;
#10;x=622416352;
#10;x=622516352;
#10;x=622616352;
#10;x=622716352;
#10;x=622816352;
#10;x=622916352;
#10;x=623016352;
#10;x=623116352;
#10;x=623216352;
#10;x=623316352;
#10;x=623416352;
#10;x=623516352;
#10;x=623616352;
#10;x=623716352;
#10;x=623816352;
#10;x=623916352;
#10;x=624016352;
#10;x=624116352;
#10;x=624216352;
#10;x=624316352;
#10;x=624416352;
#10;x=624516352;
#10;x=624616352;
#10;x=624716352;
#10;x=624816352;
#10;x=624916352;
#10;x=625016352;
#10;x=625116352;
#10;x=625216352;
#10;x=625316352;
#10;x=625416352;
#10;x=625516352;
#10;x=625616352;
#10;x=625716352;
#10;x=625816352;
#10;x=625916352;
#10;x=626016352;
#10;x=626116352;
#10;x=626216352;
#10;x=626316352;
#10;x=626416352;
#10;x=626516352;
#10;x=626616352;
#10;x=626716352;
#10;x=626816352;
#10;x=626916352;
#10;x=627016352;
#10;x=627116352;
#10;x=627216352;
#10;x=627316352;
#10;x=627416352;
#10;x=627516352;
#10;x=627616352;
#10;x=627716352;
#10;x=627816352;
#10;x=627916352;
#10;x=628016352;
#10;x=628116352;
#10;x=628216352;
#10;x=628316352;
#10;x=628416352;
#10;x=628516352;
#10;x=628616352;
#10;x=628716352;
#10;x=628816352;
#10;x=628916352;
#10;x=629016352;
#10;x=629116352;
#10;x=629216352;
#10;x=629316352;
#10;x=629416352;
#10;x=629516352;
#10;x=629616352;
#10;x=629716352;
#10;x=629816352;
#10;x=629916352;
#10;x=630016352;
#10;x=630116352;
#10;x=630216352;
#10;x=630316352;
#10;x=630416352;
#10;x=630516352;
#10;x=630616352;
#10;x=630716352;
#10;x=630816352;
#10;x=630916352;
#10;x=631016352;
#10;x=631116352;
#10;x=631216352;
#10;x=631316352;
#10;x=631416352;
#10;x=631516352;
#10;x=631616352;
#10;x=631716352;
#10;x=631816352;
#10;x=631916352;
#10;x=632016352;
#10;x=632116352;
#10;x=632216352;
#10;x=632316352;
#10;x=632416352;
#10;x=632516352;
#10;x=632616352;
#10;x=632716352;
#10;x=632816352;
#10;x=632916352;
#10;x=633016352;
#10;x=633116352;
#10;x=633216352;
#10;x=633316352;
#10;x=633416352;
#10;x=633516352;
#10;x=633616352;
#10;x=633716352;
#10;x=633816352;
#10;x=633916352;
#10;x=634016352;
#10;x=634116352;
#10;x=634216352;
#10;x=634316352;
#10;x=634416352;
#10;x=634516352;
#10;x=634616352;
#10;x=634716352;
#10;x=634816352;
#10;x=634916352;
#10;x=635016352;
#10;x=635116352;
#10;x=635216352;
#10;x=635316352;
#10;x=635416352;
#10;x=635516352;
#10;x=635616352;
#10;x=635716352;
#10;x=635816352;
#10;x=635916352;
#10;x=636016352;
#10;x=636116352;
#10;x=636216352;
#10;x=636316352;
#10;x=636416352;
#10;x=636516352;
#10;x=636616352;
#10;x=636716352;
#10;x=636816352;
#10;x=636916352;
#10;x=637016352;
#10;x=637116352;
#10;x=637216352;
#10;x=637316352;
#10;x=637416352;
#10;x=637516352;
#10;x=637616352;
#10;x=637716352;
#10;x=637816352;
#10;x=637916352;
#10;x=638016352;
#10;x=638116352;
#10;x=638216352;
#10;x=638316352;
#10;x=638416352;
#10;x=638516352;
#10;x=638616352;
#10;x=638716352;
#10;x=638816352;
#10;x=638916352;
#10;x=639016352;
#10;x=639116352;
#10;x=639216352;
#10;x=639316352;
#10;x=639416352;
#10;x=639516352;
#10;x=639616352;
#10;x=639716352;
#10;x=639816352;
#10;x=639916352;
#10;x=640016352;
#10;x=640116352;
#10;x=640216352;
#10;x=640316352;
#10;x=640416352;
#10;x=640516352;
#10;x=640616352;
#10;x=640716352;
#10;x=640816352;
#10;x=640916352;
#10;x=641016352;
#10;x=641116352;
#10;x=641216352;
#10;x=641316352;
#10;x=641416352;
#10;x=641516352;
#10;x=641616352;
#10;x=641716352;
#10;x=641816352;
#10;x=641916352;
#10;x=642016352;
#10;x=642116352;
#10;x=642216352;
#10;x=642316352;
#10;x=642416352;
#10;x=642516352;
#10;x=642616352;
#10;x=642716352;
#10;x=642816352;
#10;x=642916352;
#10;x=643016352;
#10;x=643116352;
#10;x=643216352;
#10;x=643316352;
#10;x=643416352;
#10;x=643516352;
#10;x=643616352;
#10;x=643716352;
#10;x=643816352;
#10;x=643916352;
#10;x=644016352;
#10;x=644116352;
#10;x=644216352;
#10;x=644316352;
#10;x=644416352;
#10;x=644516352;
#10;x=644616352;
#10;x=644716352;
#10;x=644816352;
#10;x=644916352;
#10;x=645016352;
#10;x=645116352;
#10;x=645216352;
#10;x=645316352;
#10;x=645416352;
#10;x=645516352;
#10;x=645616352;
#10;x=645716352;
#10;x=645816352;
#10;x=645916352;
#10;x=646016352;
#10;x=646116352;
#10;x=646216352;
#10;x=646316352;
#10;x=646416352;
#10;x=646516352;
#10;x=646616352;
#10;x=646716352;
#10;x=646816352;
#10;x=646916352;
#10;x=647016352;
#10;x=647116352;
#10;x=647216352;
#10;x=647316352;
#10;x=647416352;
#10;x=647516352;
#10;x=647616352;
#10;x=647716352;
#10;x=647816352;
#10;x=647916352;
#10;x=648016352;
#10;x=648116352;
#10;x=648216352;
#10;x=648316352;
#10;x=648416352;
#10;x=648516352;
#10;x=648616352;
#10;x=648716352;
#10;x=648816352;
#10;x=648916352;
#10;x=649016352;
#10;x=649116352;
#10;x=649216352;
#10;x=649316352;
#10;x=649416352;
#10;x=649516352;
#10;x=649616352;
#10;x=649716352;
#10;x=649816352;
#10;x=649916352;
#10;x=650016352;
#10;x=650116352;
#10;x=650216352;
#10;x=650316352;
#10;x=650416352;
#10;x=650516352;
#10;x=650616352;
#10;x=650716352;
#10;x=650816352;
#10;x=650916352;
#10;x=651016352;
#10;x=651116352;
#10;x=651216352;
#10;x=651316352;
#10;x=651416352;
#10;x=651516352;
#10;x=651616352;
#10;x=651716352;
#10;x=651816352;
#10;x=651916352;
#10;x=652016352;
#10;x=652116352;
#10;x=652216352;
#10;x=652316352;
#10;x=652416352;
#10;x=652516352;
#10;x=652616352;
#10;x=652716352;
#10;x=652816352;
#10;x=652916352;
#10;x=653016352;
#10;x=653116352;
#10;x=653216352;
#10;x=653316352;
#10;x=653416352;
#10;x=653516352;
#10;x=653616352;
#10;x=653716352;
#10;x=653816352;
#10;x=653916352;
#10;x=654016352;
#10;x=654116352;
#10;x=654216352;
#10;x=654316352;
#10;x=654416352;
#10;x=654516352;
#10;x=654616352;
#10;x=654716352;
#10;x=654816352;
#10;x=654916352;
#10;x=655016352;
#10;x=655116352;
#10;x=655216352;
#10;x=655316352;
#10;x=655416352;
#10;x=655516352;
#10;x=655616352;
#10;x=655716352;
#10;x=655816352;
#10;x=655916352;
#10;x=656016352;
#10;x=656116352;
#10;x=656216352;
#10;x=656316352;
#10;x=656416352;
#10;x=656516352;
#10;x=656616352;
#10;x=656716352;
#10;x=656816352;
#10;x=656916352;
#10;x=657016352;
#10;x=657116352;
#10;x=657216352;
#10;x=657316352;
#10;x=657416352;
#10;x=657516352;
#10;x=657616352;
#10;x=657716352;
#10;x=657816352;
#10;x=657916352;
#10;x=658016352;
#10;x=658116352;
#10;x=658216352;
#10;x=658316352;
#10;x=658416352;
#10;x=658516352;
#10;x=658616352;
#10;x=658716352;
#10;x=658816352;
#10;x=658916352;
#10;x=659016352;
#10;x=659116352;
#10;x=659216352;
#10;x=659316352;
#10;x=659416352;
#10;x=659516352;
#10;x=659616352;
#10;x=659716352;
#10;x=659816352;
#10;x=659916352;
#10;x=660016352;
#10;x=660116352;
#10;x=660216352;
#10;x=660316352;
#10;x=660416352;
#10;x=660516352;
#10;x=660616352;
#10;x=660716352;
#10;x=660816352;
#10;x=660916352;
#10;x=661016352;
#10;x=661116352;
#10;x=661216352;
#10;x=661316352;
#10;x=661416352;
#10;x=661516352;
#10;x=661616352;
#10;x=661716352;
#10;x=661816352;
#10;x=661916352;
#10;x=662016352;
#10;x=662116352;
#10;x=662216352;
#10;x=662316352;
#10;x=662416352;
#10;x=662516352;
#10;x=662616352;
#10;x=662716352;
#10;x=662816352;
#10;x=662916352;
#10;x=663016352;
#10;x=663116352;
#10;x=663216352;
#10;x=663316352;
#10;x=663416352;
#10;x=663516352;
#10;x=663616352;
#10;x=663716352;
#10;x=663816352;
#10;x=663916352;
#10;x=664016352;
#10;x=664116352;
#10;x=664216352;
#10;x=664316352;
#10;x=664416352;
#10;x=664516352;
#10;x=664616352;
#10;x=664716352;
#10;x=664816352;
#10;x=664916352;
#10;x=665016352;
#10;x=665116352;
#10;x=665216352;
#10;x=665316352;
#10;x=665416352;
#10;x=665516352;
#10;x=665616352;
#10;x=665716352;
#10;x=665816352;
#10;x=665916352;
#10;x=666016352;
#10;x=666116352;
#10;x=666216352;
#10;x=666316352;
#10;x=666416352;
#10;x=666516352;
#10;x=666616352;
#10;x=666716352;
#10;x=666816352;
#10;x=666916352;
#10;x=667016352;
#10;x=667116352;
#10;x=667216352;
#10;x=667316352;
#10;x=667416352;
#10;x=667516352;
#10;x=667616352;
#10;x=667716352;
#10;x=667816352;
#10;x=667916352;
#10;x=668016352;
#10;x=668116352;
#10;x=668216352;
#10;x=668316352;
#10;x=668416352;
#10;x=668516352;
#10;x=668616352;
#10;x=668716352;
#10;x=668816352;
#10;x=668916352;
#10;x=669016352;
#10;x=669116352;
#10;x=669216352;
#10;x=669316352;
#10;x=669416352;
#10;x=669516352;
#10;x=669616352;
#10;x=669716352;
#10;x=669816352;
#10;x=669916352;
#10;x=670016352;
#10;x=670116352;
#10;x=670216352;
#10;x=670316352;
#10;x=670416352;
#10;x=670516352;
#10;x=670616352;
#10;x=670716352;
#10;x=670816352;
#10;x=670916352;
#10;x=671016352;
#10;x=671116352;
#10;x=671216352;
#10;x=671316352;
#10;x=671416352;
#10;x=671516352;
#10;x=671616352;
#10;x=671716352;
#10;x=671816352;
#10;x=671916352;
#10;x=672016352;
#10;x=672116352;
#10;x=672216352;
#10;x=672316352;
#10;x=672416352;
#10;x=672516352;
#10;x=672616352;
#10;x=672716352;
#10;x=672816352;
#10;x=672916352;
#10;x=673016352;
#10;x=673116352;
#10;x=673216352;
#10;x=673316352;
#10;x=673416352;
#10;x=673516352;
#10;x=673616352;
#10;x=673716352;
#10;x=673816352;
#10;x=673916352;
#10;x=674016352;
#10;x=674116352;
#10;x=674216352;
#10;x=674316352;
#10;x=674416352;
#10;x=674516352;
#10;x=674616352;
#10;x=674716352;
#10;x=674816352;
#10;x=674916352;
#10;x=675016352;
#10;x=675116352;
#10;x=675216352;
#10;x=675316352;
#10;x=675416352;
#10;x=675516352;
#10;x=675616352;
#10;x=675716352;
#10;x=675816352;
#10;x=675916352;
#10;x=676016352;
#10;x=676116352;
#10;x=676216352;
#10;x=676316352;
#10;x=676416352;
#10;x=676516352;
#10;x=676616352;
#10;x=676716352;
#10;x=676816352;
#10;x=676916352;
#10;x=677016352;
#10;x=677116352;
#10;x=677216352;
#10;x=677316352;
#10;x=677416352;
#10;x=677516352;
#10;x=677616352;
#10;x=677716352;
#10;x=677816352;
#10;x=677916352;
#10;x=678016352;
#10;x=678116352;
#10;x=678216352;
#10;x=678316352;
#10;x=678416352;
#10;x=678516352;
#10;x=678616352;
#10;x=678716352;
#10;x=678816352;
#10;x=678916352;
#10;x=679016352;
#10;x=679116352;
#10;x=679216352;
#10;x=679316352;
#10;x=679416352;
#10;x=679516352;
#10;x=679616352;
#10;x=679716352;
#10;x=679816352;
#10;x=679916352;
#10;x=680016352;
#10;x=680116352;
#10;x=680216352;
#10;x=680316352;
#10;x=680416352;
#10;x=680516352;
#10;x=680616352;
#10;x=680716352;
#10;x=680816352;
#10;x=680916352;
#10;x=681016352;
#10;x=681116352;
#10;x=681216352;
#10;x=681316352;
#10;x=681416352;
#10;x=681516352;
#10;x=681616352;
#10;x=681716352;
#10;x=681816352;
#10;x=681916352;
#10;x=682016352;
#10;x=682116352;
#10;x=682216352;
#10;x=682316352;
#10;x=682416352;
#10;x=682516352;
#10;x=682616352;
#10;x=682716352;
#10;x=682816352;
#10;x=682916352;
#10;x=683016352;
#10;x=683116352;
#10;x=683216352;
#10;x=683316352;
#10;x=683416352;
#10;x=683516352;
#10;x=683616352;
#10;x=683716352;
#10;x=683816352;
#10;x=683916352;
#10;x=684016352;
#10;x=684116352;
#10;x=684216352;
#10;x=684316352;
#10;x=684416352;
#10;x=684516352;
#10;x=684616352;
#10;x=684716352;
#10;x=684816352;
#10;x=684916352;
#10;x=685016352;
#10;x=685116352;
#10;x=685216352;
#10;x=685316352;
#10;x=685416352;
#10;x=685516352;
#10;x=685616352;
#10;x=685716352;
#10;x=685816352;
#10;x=685916352;
#10;x=686016352;
#10;x=686116352;
#10;x=686216352;
#10;x=686316352;
#10;x=686416352;
#10;x=686516352;
#10;x=686616352;
#10;x=686716352;
#10;x=686816352;
#10;x=686916352;
#10;x=687016352;
#10;x=687116352;
#10;x=687216352;
#10;x=687316352;
#10;x=687416352;
#10;x=687516352;
#10;x=687616352;
#10;x=687716352;
#10;x=687816352;
#10;x=687916352;
#10;x=688016352;
#10;x=688116352;
#10;x=688216352;
#10;x=688316352;
#10;x=688416352;
#10;x=688516352;
#10;x=688616352;
#10;x=688716352;
#10;x=688816352;
#10;x=688916352;
#10;x=689016352;
#10;x=689116352;
#10;x=689216352;
#10;x=689316352;
#10;x=689416352;
#10;x=689516352;
#10;x=689616352;
#10;x=689716352;
#10;x=689816352;
#10;x=689916352;
#10;x=690016352;
#10;x=690116352;
#10;x=690216352;
#10;x=690316352;
#10;x=690416352;
#10;x=690516352;
#10;x=690616352;
#10;x=690716352;
#10;x=690816352;
#10;x=690916352;
#10;x=691016352;
#10;x=691116352;
#10;x=691216352;
#10;x=691316352;
#10;x=691416352;
#10;x=691516352;
#10;x=691616352;
#10;x=691716352;
#10;x=691816352;
#10;x=691916352;
#10;x=692016352;
#10;x=692116352;
#10;x=692216352;
#10;x=692316352;
#10;x=692416352;
#10;x=692516352;
#10;x=692616352;
#10;x=692716352;
#10;x=692816352;
#10;x=692916352;
#10;x=693016352;
#10;x=693116352;
#10;x=693216352;
#10;x=693316352;
#10;x=693416352;
#10;x=693516352;
#10;x=693616352;
#10;x=693716352;
#10;x=693816352;
#10;x=693916352;
#10;x=694016352;
#10;x=694116352;
#10;x=694216352;
#10;x=694316352;
#10;x=694416352;
#10;x=694516352;
#10;x=694616352;
#10;x=694716352;
#10;x=694816352;
#10;x=694916352;
#10;x=695016352;
#10;x=695116352;
#10;x=695216352;
#10;x=695316352;
#10;x=695416352;
#10;x=695516352;
#10;x=695616352;
#10;x=695716352;
#10;x=695816352;
#10;x=695916352;
#10;x=696016352;
#10;x=696116352;
#10;x=696216352;
#10;x=696316352;
#10;x=696416352;
#10;x=696516352;
#10;x=696616352;
#10;x=696716352;
#10;x=696816352;
#10;x=696916352;
#10;x=697016352;
#10;x=697116352;
#10;x=697216352;
#10;x=697316352;
#10;x=697416352;
#10;x=697516352;
#10;x=697616352;
#10;x=697716352;
#10;x=697816352;
#10;x=697916352;
#10;x=698016352;
#10;x=698116352;
#10;x=698216352;
#10;x=698316352;
#10;x=698416352;
#10;x=698516352;
#10;x=698616352;
#10;x=698716352;
#10;x=698816352;
#10;x=698916352;
#10;x=699016352;
#10;x=699116352;
#10;x=699216352;
#10;x=699316352;
#10;x=699416352;
#10;x=699516352;
#10;x=699616352;
#10;x=699716352;
#10;x=699816352;
#10;x=699916352;
#10;x=700016352;
#10;x=700116352;
#10;x=700216352;
#10;x=700316352;
#10;x=700416352;
#10;x=700516352;
#10;x=700616352;
#10;x=700716352;
#10;x=700816352;
#10;x=700916352;
#10;x=701016352;
#10;x=701116352;
#10;x=701216352;
#10;x=701316352;
#10;x=701416352;
#10;x=701516352;
#10;x=701616352;
#10;x=701716352;
#10;x=701816352;
#10;x=701916352;
#10;x=702016352;
#10;x=702116352;
#10;x=702216352;
#10;x=702316352;
#10;x=702416352;
#10;x=702516352;
#10;x=702616352;
#10;x=702716352;
#10;x=702816352;
#10;x=702916352;
#10;x=703016352;
#10;x=703116352;
#10;x=703216352;
#10;x=703316352;
#10;x=703416352;
#10;x=703516352;
#10;x=703616352;
#10;x=703716352;
#10;x=703816352;
#10;x=703916352;
#10;x=704016352;
#10;x=704116352;
#10;x=704216352;
#10;x=704316352;
#10;x=704416352;
#10;x=704516352;
#10;x=704616352;
#10;x=704716352;
#10;x=704816352;
#10;x=704916352;
#10;x=705016352;
#10;x=705116352;
#10;x=705216352;
#10;x=705316352;
#10;x=705416352;
#10;x=705516352;
#10;x=705616352;
#10;x=705716352;
#10;x=705816352;
#10;x=705916352;
#10;x=706016352;
#10;x=706116352;
#10;x=706216352;
#10;x=706316352;
#10;x=706416352;
#10;x=706516352;
#10;x=706616352;
#10;x=706716352;
#10;x=706816352;
#10;x=706916352;
#10;x=707016352;
#10;x=707116352;
#10;x=707216352;
#10;x=707316352;
#10;x=707416352;
#10;x=707516352;
#10;x=707616352;
#10;x=707716352;
#10;x=707816352;
#10;x=707916352;
#10;x=708016352;
#10;x=708116352;
#10;x=708216352;
#10;x=708316352;
#10;x=708416352;
#10;x=708516352;
#10;x=708616352;
#10;x=708716352;
#10;x=708816352;
#10;x=708916352;
#10;x=709016352;
#10;x=709116352;
#10;x=709216352;
#10;x=709316352;
#10;x=709416352;
#10;x=709516352;
#10;x=709616352;
#10;x=709716352;
#10;x=709816352;
#10;x=709916352;
#10;x=710016352;
#10;x=710116352;
#10;x=710216352;
#10;x=710316352;
#10;x=710416352;
#10;x=710516352;
#10;x=710616352;
#10;x=710716352;
#10;x=710816352;
#10;x=710916352;
#10;x=711016352;
#10;x=711116352;
#10;x=711216352;
#10;x=711316352;
#10;x=711416352;
#10;x=711516352;
#10;x=711616352;
#10;x=711716352;
#10;x=711816352;
#10;x=711916352;
#10;x=712016352;
#10;x=712116352;
#10;x=712216352;
#10;x=712316352;
#10;x=712416352;
#10;x=712516352;
#10;x=712616352;
#10;x=712716352;
#10;x=712816352;
#10;x=712916352;
#10;x=713016352;
#10;x=713116352;
#10;x=713216352;
#10;x=713316352;
#10;x=713416352;
#10;x=713516352;
#10;x=713616352;
#10;x=713716352;
#10;x=713816352;
#10;x=713916352;
#10;x=714016352;
#10;x=714116352;
#10;x=714216352;
#10;x=714316352;
#10;x=714416352;
#10;x=714516352;
#10;x=714616352;
#10;x=714716352;
#10;x=714816352;
#10;x=714916352;
#10;x=715016352;
#10;x=715116352;
#10;x=715216352;
#10;x=715316352;
#10;x=715416352;
#10;x=715516352;
#10;x=715616352;
#10;x=715716352;
#10;x=715816352;
#10;x=715916352;
#10;x=716016352;
#10;x=716116352;
#10;x=716216352;
#10;x=716316352;
#10;x=716416352;
#10;x=716516352;
#10;x=716616352;
#10;x=716716352;
#10;x=716816352;
#10;x=716916352;
#10;x=717016352;
#10;x=717116352;
#10;x=717216352;
#10;x=717316352;
#10;x=717416352;
#10;x=717516352;
#10;x=717616352;
#10;x=717716352;
#10;x=717816352;
#10;x=717916352;
#10;x=718016352;
#10;x=718116352;
#10;x=718216352;
#10;x=718316352;
#10;x=718416352;
#10;x=718516352;
#10;x=718616352;
#10;x=718716352;
#10;x=718816352;
#10;x=718916352;
#10;x=719016352;
#10;x=719116352;
#10;x=719216352;
#10;x=719316352;
#10;x=719416352;
#10;x=719516352;
#10;x=719616352;
#10;x=719716352;
#10;x=719816352;
#10;x=719916352;
#10;x=720016352;
#10;x=720116352;
#10;x=720216352;
#10;x=720316352;
#10;x=720416352;
#10;x=720516352;
#10;x=720616352;
#10;x=720716352;
#10;x=720816352;
#10;x=720916352;
#10;x=721016352;
#10;x=721116352;
#10;x=721216352;
#10;x=721316352;
#10;x=721416352;
#10;x=721516352;
#10;x=721616352;
#10;x=721716352;
#10;x=721816352;
#10;x=721916352;
#10;x=722016352;
#10;x=722116352;
#10;x=722216352;
#10;x=722316352;
#10;x=722416352;
#10;x=722516352;
#10;x=722616352;
#10;x=722716352;
#10;x=722816352;
#10;x=722916352;
#10;x=723016352;
#10;x=723116352;
#10;x=723216352;
#10;x=723316352;
#10;x=723416352;
#10;x=723516352;
#10;x=723616352;
#10;x=723716352;
#10;x=723816352;
#10;x=723916352;
#10;x=724016352;
#10;x=724116352;
#10;x=724216352;
#10;x=724316352;
#10;x=724416352;
#10;x=724516352;
#10;x=724616352;
#10;x=724716352;
#10;x=724816352;
#10;x=724916352;
#10;x=725016352;
#10;x=725116352;
#10;x=725216352;
#10;x=725316352;
#10;x=725416352;
#10;x=725516352;
#10;x=725616352;
#10;x=725716352;
#10;x=725816352;
#10;x=725916352;
#10;x=726016352;
#10;x=726116352;
#10;x=726216352;
#10;x=726316352;
#10;x=726416352;
#10;x=726516352;
#10;x=726616352;
#10;x=726716352;
#10;x=726816352;
#10;x=726916352;
#10;x=727016352;
#10;x=727116352;
#10;x=727216352;
#10;x=727316352;
#10;x=727416352;
#10;x=727516352;
#10;x=727616352;
#10;x=727716352;
#10;x=727816352;
#10;x=727916352;
#10;x=728016352;
#10;x=728116352;
#10;x=728216352;
#10;x=728316352;
#10;x=728416352;
#10;x=728516352;
#10;x=728616352;
#10;x=728716352;
#10;x=728816352;
#10;x=728916352;
#10;x=729016352;
#10;x=729116352;
#10;x=729216352;
#10;x=729316352;
#10;x=729416352;
#10;x=729516352;
#10;x=729616352;
#10;x=729716352;
#10;x=729816352;
#10;x=729916352;
#10;x=730016352;
#10;x=730116352;
#10;x=730216352;
#10;x=730316352;
#10;x=730416352;
#10;x=730516352;
#10;x=730616352;
#10;x=730716352;
#10;x=730816352;
#10;x=730916352;
#10;x=731016352;
#10;x=731116352;
#10;x=731216352;
#10;x=731316352;
#10;x=731416352;
#10;x=731516352;
#10;x=731616352;
#10;x=731716352;
#10;x=731816352;
#10;x=731916352;
#10;x=732016352;
#10;x=732116352;
#10;x=732216352;
#10;x=732316352;
#10;x=732416352;
#10;x=732516352;
#10;x=732616352;
#10;x=732716352;
#10;x=732816352;
#10;x=732916352;
#10;x=733016352;
#10;x=733116352;
#10;x=733216352;
#10;x=733316352;
#10;x=733416352;
#10;x=733516352;
#10;x=733616352;
#10;x=733716352;
#10;x=733816352;
#10;x=733916352;
#10;x=734016352;
#10;x=734116352;
#10;x=734216352;
#10;x=734316352;
#10;x=734416352;
#10;x=734516352;
#10;x=734616352;
#10;x=734716352;
#10;x=734816352;
#10;x=734916352;
#10;x=735016352;
#10;x=735116352;
#10;x=735216352;
#10;x=735316352;
#10;x=735416352;
#10;x=735516352;
#10;x=735616352;
#10;x=735716352;
#10;x=735816352;
#10;x=735916352;
#10;x=736016352;
#10;x=736116352;
#10;x=736216352;
#10;x=736316352;
#10;x=736416352;
#10;x=736516352;
#10;x=736616352;
#10;x=736716352;
#10;x=736816352;
#10;x=736916352;
#10;x=737016352;
#10;x=737116352;
#10;x=737216352;
#10;x=737316352;
#10;x=737416352;
#10;x=737516352;
#10;x=737616352;
#10;x=737716352;
#10;x=737816352;
#10;x=737916352;
#10;x=738016352;
#10;x=738116352;
#10;x=738216352;
#10;x=738316352;
#10;x=738416352;
#10;x=738516352;
#10;x=738616352;
#10;x=738716352;
#10;x=738816352;
#10;x=738916352;
#10;x=739016352;
#10;x=739116352;
#10;x=739216352;
#10;x=739316352;
#10;x=739416352;
#10;x=739516352;
#10;x=739616352;
#10;x=739716352;
#10;x=739816352;
#10;x=739916352;
#10;x=740016352;
#10;x=740116352;
#10;x=740216352;
#10;x=740316352;
#10;x=740416352;
#10;x=740516352;
#10;x=740616352;
#10;x=740716352;
#10;x=740816352;
#10;x=740916352;
#10;x=741016352;
#10;x=741116352;
#10;x=741216352;
#10;x=741316352;
#10;x=741416352;
#10;x=741516352;
#10;x=741616352;
#10;x=741716352;
#10;x=741816352;
#10;x=741916352;
#10;x=742016352;
#10;x=742116352;
#10;x=742216352;
#10;x=742316352;
#10;x=742416352;
#10;x=742516352;
#10;x=742616352;
#10;x=742716352;
#10;x=742816352;
#10;x=742916352;
#10;x=743016352;
#10;x=743116352;
#10;x=743216352;
#10;x=743316352;
#10;x=743416352;
#10;x=743516352;
#10;x=743616352;
#10;x=743716352;
#10;x=743816352;
#10;x=743916352;
#10;x=744016352;
#10;x=744116352;
#10;x=744216352;
#10;x=744316352;
#10;x=744416352;
#10;x=744516352;
#10;x=744616352;
#10;x=744716352;
#10;x=744816352;
#10;x=744916352;
#10;x=745016352;
#10;x=745116352;
#10;x=745216352;
#10;x=745316352;
#10;x=745416352;
#10;x=745516352;
#10;x=745616352;
#10;x=745716352;
#10;x=745816352;
#10;x=745916352;
#10;x=746016352;
#10;x=746116352;
#10;x=746216352;
#10;x=746316352;
#10;x=746416352;
#10;x=746516352;
#10;x=746616352;
#10;x=746716352;
#10;x=746816352;
#10;x=746916352;
#10;x=747016352;
#10;x=747116352;
#10;x=747216352;
#10;x=747316352;
#10;x=747416352;
#10;x=747516352;
#10;x=747616352;
#10;x=747716352;
#10;x=747816352;
#10;x=747916352;
#10;x=748016352;
#10;x=748116352;
#10;x=748216352;
#10;x=748316352;
#10;x=748416352;
#10;x=748516352;
#10;x=748616352;
#10;x=748716352;
#10;x=748816352;
#10;x=748916352;
#10;x=749016352;
#10;x=749116352;
#10;x=749216352;
#10;x=749316352;
#10;x=749416352;
#10;x=749516352;
#10;x=749616352;
#10;x=749716352;
#10;x=749816352;
#10;x=749916352;
#10;x=750016352;
#10;x=750116352;
#10;x=750216352;
#10;x=750316352;
#10;x=750416352;
#10;x=750516352;
#10;x=750616352;
#10;x=750716352;
#10;x=750816352;
#10;x=750916352;
#10;x=751016352;
#10;x=751116352;
#10;x=751216352;
#10;x=751316352;
#10;x=751416352;
#10;x=751516352;
#10;x=751616352;
#10;x=751716352;
#10;x=751816352;
#10;x=751916352;
#10;x=752016352;
#10;x=752116352;
#10;x=752216352;
#10;x=752316352;
#10;x=752416352;
#10;x=752516352;
#10;x=752616352;
#10;x=752716352;
#10;x=752816352;
#10;x=752916352;
#10;x=753016352;
#10;x=753116352;
#10;x=753216352;
#10;x=753316352;
#10;x=753416352;
#10;x=753516352;
#10;x=753616352;
#10;x=753716352;
#10;x=753816352;
#10;x=753916352;
#10;x=754016352;
#10;x=754116352;
#10;x=754216352;
#10;x=754316352;
#10;x=754416352;
#10;x=754516352;
#10;x=754616352;
#10;x=754716352;
#10;x=754816352;
#10;x=754916352;
#10;x=755016352;
#10;x=755116352;
#10;x=755216352;
#10;x=755316352;
#10;x=755416352;
#10;x=755516352;
#10;x=755616352;
#10;x=755716352;
#10;x=755816352;
#10;x=755916352;
#10;x=756016352;
#10;x=756116352;
#10;x=756216352;
#10;x=756316352;
#10;x=756416352;
#10;x=756516352;
#10;x=756616352;
#10;x=756716352;
#10;x=756816352;
#10;x=756916352;
#10;x=757016352;
#10;x=757116352;
#10;x=757216352;
#10;x=757316352;
#10;x=757416352;
#10;x=757516352;
#10;x=757616352;
#10;x=757716352;
#10;x=757816352;
#10;x=757916352;
#10;x=758016352;
#10;x=758116352;
#10;x=758216352;
#10;x=758316352;
#10;x=758416352;
#10;x=758516352;
#10;x=758616352;
#10;x=758716352;
#10;x=758816352;
#10;x=758916352;
#10;x=759016352;
#10;x=759116352;
#10;x=759216352;
#10;x=759316352;
#10;x=759416352;
#10;x=759516352;
#10;x=759616352;
#10;x=759716352;
#10;x=759816352;
#10;x=759916352;
#10;x=760016352;
#10;x=760116352;
#10;x=760216352;
#10;x=760316352;
#10;x=760416352;
#10;x=760516352;
#10;x=760616352;
#10;x=760716352;
#10;x=760816352;
#10;x=760916352;
#10;x=761016352;
#10;x=761116352;
#10;x=761216352;
#10;x=761316352;
#10;x=761416352;
#10;x=761516352;
#10;x=761616352;
#10;x=761716352;
#10;x=761816352;
#10;x=761916352;
#10;x=762016352;
#10;x=762116352;
#10;x=762216352;
#10;x=762316352;
#10;x=762416352;
#10;x=762516352;
#10;x=762616352;
#10;x=762716352;
#10;x=762816352;
#10;x=762916352;
#10;x=763016352;
#10;x=763116352;
#10;x=763216352;
#10;x=763316352;
#10;x=763416352;
#10;x=763516352;
#10;x=763616352;
#10;x=763716352;
#10;x=763816352;
#10;x=763916352;
#10;x=764016352;
#10;x=764116352;
#10;x=764216352;
#10;x=764316352;
#10;x=764416352;
#10;x=764516352;
#10;x=764616352;
#10;x=764716352;
#10;x=764816352;
#10;x=764916352;
#10;x=765016352;
#10;x=765116352;
#10;x=765216352;
#10;x=765316352;
#10;x=765416352;
#10;x=765516352;
#10;x=765616352;
#10;x=765716352;
#10;x=765816352;
#10;x=765916352;
#10;x=766016352;
#10;x=766116352;
#10;x=766216352;
#10;x=766316352;
#10;x=766416352;
#10;x=766516352;
#10;x=766616352;
#10;x=766716352;
#10;x=766816352;
#10;x=766916352;
#10;x=767016352;
#10;x=767116352;
#10;x=767216352;
#10;x=767316352;
#10;x=767416352;
#10;x=767516352;
#10;x=767616352;
#10;x=767716352;
#10;x=767816352;
#10;x=767916352;
#10;x=768016352;
#10;x=768116352;
#10;x=768216352;
#10;x=768316352;
#10;x=768416352;
#10;x=768516352;
#10;x=768616352;
#10;x=768716352;
#10;x=768816352;
#10;x=768916352;
#10;x=769016352;
#10;x=769116352;
#10;x=769216352;
#10;x=769316352;
#10;x=769416352;
#10;x=769516352;
#10;x=769616352;
#10;x=769716352;
#10;x=769816352;
#10;x=769916352;
#10;x=770016352;
#10;x=770116352;
#10;x=770216352;
#10;x=770316352;
#10;x=770416352;
#10;x=770516352;
#10;x=770616352;
#10;x=770716352;
#10;x=770816352;
#10;x=770916352;
#10;x=771016352;
#10;x=771116352;
#10;x=771216352;
#10;x=771316352;
#10;x=771416352;
#10;x=771516352;
#10;x=771616352;
#10;x=771716352;
#10;x=771816352;
#10;x=771916352;
#10;x=772016352;
#10;x=772116352;
#10;x=772216352;
#10;x=772316352;
#10;x=772416352;
#10;x=772516352;
#10;x=772616352;
#10;x=772716352;
#10;x=772816352;
#10;x=772916352;
#10;x=773016352;
#10;x=773116352;
#10;x=773216352;
#10;x=773316352;
#10;x=773416352;
#10;x=773516352;
#10;x=773616352;
#10;x=773716352;
#10;x=773816352;
#10;x=773916352;
#10;x=774016352;
#10;x=774116352;
#10;x=774216352;
#10;x=774316352;
#10;x=774416352;
#10;x=774516352;
#10;x=774616352;
#10;x=774716352;
#10;x=774816352;
#10;x=774916352;
#10;x=775016352;
#10;x=775116352;
#10;x=775216352;
#10;x=775316352;
#10;x=775416352;
#10;x=775516352;
#10;x=775616352;
#10;x=775716352;
#10;x=775816352;
#10;x=775916352;
#10;x=776016352;
#10;x=776116352;
#10;x=776216352;
#10;x=776316352;
#10;x=776416352;
#10;x=776516352;
#10;x=776616352;
#10;x=776716352;
#10;x=776816352;
#10;x=776916352;
#10;x=777016352;
#10;x=777116352;
#10;x=777216352;
#10;x=777316352;
#10;x=777416352;
#10;x=777516352;
#10;x=777616352;
#10;x=777716352;
#10;x=777816352;
#10;x=777916352;
#10;x=778016352;
#10;x=778116352;
#10;x=778216352;
#10;x=778316352;
#10;x=778416352;
#10;x=778516352;
#10;x=778616352;
#10;x=778716352;
#10;x=778816352;
#10;x=778916352;
#10;x=779016352;
#10;x=779116352;
#10;x=779216352;
#10;x=779316352;
#10;x=779416352;
#10;x=779516352;
#10;x=779616352;
#10;x=779716352;
#10;x=779816352;
#10;x=779916352;
#10;x=780016352;
#10;x=780116352;
#10;x=780216352;
#10;x=780316352;
#10;x=780416352;
#10;x=780516352;
#10;x=780616352;
#10;x=780716352;
#10;x=780816352;
#10;x=780916352;
#10;x=781016352;
#10;x=781116352;
#10;x=781216352;
#10;x=781316352;
#10;x=781416352;
#10;x=781516352;
#10;x=781616352;
#10;x=781716352;
#10;x=781816352;
#10;x=781916352;
#10;x=782016352;
#10;x=782116352;
#10;x=782216352;
#10;x=782316352;
#10;x=782416352;
#10;x=782516352;
#10;x=782616352;
#10;x=782716352;
#10;x=782816352;
#10;x=782916352;
#10;x=783016352;
#10;x=783116352;
#10;x=783216352;
#10;x=783316352;
#10;x=783416352;
#10;x=783516352;
#10;x=783616352;
#10;x=783716352;
#10;x=783816352;
#10;x=783916352;
#10;x=784016352;
#10;x=784116352;
#10;x=784216352;
#10;x=784316352;
#10;x=784416352;
#10;x=784516352;
#10;x=784616352;
#10;x=784716352;
#10;x=784816352;
#10;x=784916352;
#10;x=785016352;
#10;x=785116352;
#10;x=785216352;
#10;x=785316352;
#10;x=785416352;
#10;x=785516352;
#10;x=785616352;
#10;x=785716352;
#10;x=785816352;
#10;x=785916352;
#10;x=786016352;
#10;x=786116352;
#10;x=786216352;
#10;x=786316352;
#10;x=786416352;
#10;x=786516352;
#10;x=786616352;
#10;x=786716352;
#10;x=786816352;
#10;x=786916352;
#10;x=787016352;
#10;x=787116352;
#10;x=787216352;
#10;x=787316352;
#10;x=787416352;
#10;x=787516352;
#10;x=787616352;
#10;x=787716352;
#10;x=787816352;
#10;x=787916352;
#10;x=788016352;
#10;x=788116352;
#10;x=788216352;
#10;x=788316352;
#10;x=788416352;
#10;x=788516352;
#10;x=788616352;
#10;x=788716352;
#10;x=788816352;
#10;x=788916352;
#10;x=789016352;
#10;x=789116352;
#10;x=789216352;
#10;x=789316352;
#10;x=789416352;
#10;x=789516352;
#10;x=789616352;
#10;x=789716352;
#10;x=789816352;
#10;x=789916352;
#10;x=790016352;
#10;x=790116352;
#10;x=790216352;
#10;x=790316352;
#10;x=790416352;
#10;x=790516352;
#10;x=790616352;
#10;x=790716352;
#10;x=790816352;
#10;x=790916352;
#10;x=791016352;
#10;x=791116352;
#10;x=791216352;
#10;x=791316352;
#10;x=791416352;
#10;x=791516352;
#10;x=791616352;
#10;x=791716352;
#10;x=791816352;
#10;x=791916352;
#10;x=792016352;
#10;x=792116352;
#10;x=792216352;
#10;x=792316352;
#10;x=792416352;
#10;x=792516352;
#10;x=792616352;
#10;x=792716352;
#10;x=792816352;
#10;x=792916352;
#10;x=793016352;
#10;x=793116352;
#10;x=793216352;
#10;x=793316352;
#10;x=793416352;
#10;x=793516352;
#10;x=793616352;
#10;x=793716352;
#10;x=793816352;
#10;x=793916352;
#10;x=794016352;
#10;x=794116352;
#10;x=794216352;
#10;x=794316352;
#10;x=794416352;
#10;x=794516352;
#10;x=794616352;
#10;x=794716352;
#10;x=794816352;
#10;x=794916352;
#10;x=795016352;
#10;x=795116352;
#10;x=795216352;
#10;x=795316352;
#10;x=795416352;
#10;x=795516352;
#10;x=795616352;
#10;x=795716352;
#10;x=795816352;
#10;x=795916352;
#10;x=796016352;
#10;x=796116352;
#10;x=796216352;
#10;x=796316352;
#10;x=796416352;
#10;x=796516352;
#10;x=796616352;
#10;x=796716352;
#10;x=796816352;
#10;x=796916352;
#10;x=797016352;
#10;x=797116352;
#10;x=797216352;
#10;x=797316352;
#10;x=797416352;
#10;x=797516352;
#10;x=797616352;
#10;x=797716352;
#10;x=797816352;
#10;x=797916352;
#10;x=798016352;
#10;x=798116352;
#10;x=798216352;
#10;x=798316352;
#10;x=798416352;
#10;x=798516352;
#10;x=798616352;
#10;x=798716352;
#10;x=798816352;
#10;x=798916352;
#10;x=799016352;
#10;x=799116352;
#10;x=799216352;
#10;x=799316352;
#10;x=799416352;
#10;x=799516352;
#10;x=799616352;
#10;x=799716352;
#10;x=799816352;
#10;x=799916352;
#10;x=800016352;
#10;x=800116352;
#10;x=800216352;
#10;x=800316352;
#10;x=800416352;
#10;x=800516352;
#10;x=800616352;
#10;x=800716352;
#10;x=800816352;
#10;x=800916352;
#10;x=801016352;
#10;x=801116352;
#10;x=801216352;
#10;x=801316352;
#10;x=801416352;
#10;x=801516352;
#10;x=801616352;
#10;x=801716352;
#10;x=801816352;
#10;x=801916352;
#10;x=802016352;
#10;x=802116352;
#10;x=802216352;
#10;x=802316352;
#10;x=802416352;
#10;x=802516352;
#10;x=802616352;
#10;x=802716352;
#10;x=802816352;
#10;x=802916352;
#10;x=803016352;
#10;x=803116352;
#10;x=803216352;
#10;x=803316352;
#10;x=803416352;
#10;x=803516352;
#10;x=803616352;
#10;x=803716352;
#10;x=803816352;
#10;x=803916352;
#10;x=804016352;
#10;x=804116352;
#10;x=804216352;
#10;x=804316352;
#10;x=804416352;
#10;x=804516352;
#10;x=804616352;
#10;x=804716352;
#10;x=804816352;
#10;x=804916352;
#10;x=805016352;
#10;x=805116352;
#10;x=805216352;
#10;x=805316352;
#10;x=805416352;
#10;x=805516352;
#10;x=805616352;
#10;x=805716352;
#10;x=805816352;
#10;x=805916352;
#10;x=806016352;
#10;x=806116352;
#10;x=806216352;
#10;x=806316352;
#10;x=806416352;
#10;x=806516352;
#10;x=806616352;
#10;x=806716352;
#10;x=806816352;
#10;x=806916352;
#10;x=807016352;
#10;x=807116352;
#10;x=807216352;
#10;x=807316352;
#10;x=807416352;
#10;x=807516352;
#10;x=807616352;
#10;x=807716352;
#10;x=807816352;
#10;x=807916352;
#10;x=808016352;
#10;x=808116352;
#10;x=808216352;
#10;x=808316352;
#10;x=808416352;
#10;x=808516352;
#10;x=808616352;
#10;x=808716352;
#10;x=808816352;
#10;x=808916352;
#10;x=809016352;
#10;x=809116352;
#10;x=809216352;
#10;x=809316352;
#10;x=809416352;
#10;x=809516352;
#10;x=809616352;
#10;x=809716352;
#10;x=809816352;
#10;x=809916352;
#10;x=810016352;
#10;x=810116352;
#10;x=810216352;
#10;x=810316352;
#10;x=810416352;
#10;x=810516352;
#10;x=810616352;
#10;x=810716352;
#10;x=810816352;
#10;x=810916352;
#10;x=811016352;
#10;x=811116352;
#10;x=811216352;
#10;x=811316352;
#10;x=811416352;
#10;x=811516352;
#10;x=811616352;
#10;x=811716352;
#10;x=811816352;
#10;x=811916352;
#10;x=812016352;
#10;x=812116352;
#10;x=812216352;
#10;x=812316352;
#10;x=812416352;
#10;x=812516352;
#10;x=812616352;
#10;x=812716352;
#10;x=812816352;
#10;x=812916352;
#10;x=813016352;
#10;x=813116352;
#10;x=813216352;
#10;x=813316352;
#10;x=813416352;
#10;x=813516352;
#10;x=813616352;
#10;x=813716352;
#10;x=813816352;
#10;x=813916352;
#10;x=814016352;
#10;x=814116352;
#10;x=814216352;
#10;x=814316352;
#10;x=814416352;
#10;x=814516352;
#10;x=814616352;
#10;x=814716352;
#10;x=814816352;
#10;x=814916352;
#10;x=815016352;
#10;x=815116352;
#10;x=815216352;
#10;x=815316352;
#10;x=815416352;
#10;x=815516352;
#10;x=815616352;
#10;x=815716352;
#10;x=815816352;
#10;x=815916352;
#10;x=816016352;
#10;x=816116352;
#10;x=816216352;
#10;x=816316352;
#10;x=816416352;
#10;x=816516352;
#10;x=816616352;
#10;x=816716352;
#10;x=816816352;
#10;x=816916352;
#10;x=817016352;
#10;x=817116352;
#10;x=817216352;
#10;x=817316352;
#10;x=817416352;
#10;x=817516352;
#10;x=817616352;
#10;x=817716352;
#10;x=817816352;
#10;x=817916352;
#10;x=818016352;
#10;x=818116352;
#10;x=818216352;
#10;x=818316352;
#10;x=818416352;
#10;x=818516352;
#10;x=818616352;
#10;x=818716352;
#10;x=818816352;
#10;x=818916352;
#10;x=819016352;
#10;x=819116352;
#10;x=819216352;
#10;x=819316352;
#10;x=819416352;
#10;x=819516352;
#10;x=819616352;
#10;x=819716352;
#10;x=819816352;
#10;x=819916352;
#10;x=820016352;
#10;x=820116352;
#10;x=820216352;
#10;x=820316352;
#10;x=820416352;
#10;x=820516352;
#10;x=820616352;
#10;x=820716352;
#10;x=820816352;
#10;x=820916352;
#10;x=821016352;
#10;x=821116352;
#10;x=821216352;
#10;x=821316352;
#10;x=821416352;
#10;x=821516352;
#10;x=821616352;
#10;x=821716352;
#10;x=821816352;
#10;x=821916352;
#10;x=822016352;
#10;x=822116352;
#10;x=822216352;
#10;x=822316352;
#10;x=822416352;
#10;x=822516352;
#10;x=822616352;
#10;x=822716352;
#10;x=822816352;
#10;x=822916352;
#10;x=823016352;
#10;x=823116352;
#10;x=823216352;
#10;x=823316352;
#10;x=823416352;
#10;x=823516352;
#10;x=823616352;
#10;x=823716352;
#10;x=823816352;
#10;x=823916352;
#10;x=824016352;
#10;x=824116352;
#10;x=824216352;
#10;x=824316352;
#10;x=824416352;
#10;x=824516352;
#10;x=824616352;
#10;x=824716352;
#10;x=824816352;
#10;x=824916352;
#10;x=825016352;
#10;x=825116352;
#10;x=825216352;
#10;x=825316352;
#10;x=825416352;
#10;x=825516352;
#10;x=825616352;
#10;x=825716352;
#10;x=825816352;
#10;x=825916352;
#10;x=826016352;
#10;x=826116352;
#10;x=826216352;
#10;x=826316352;
#10;x=826416352;
#10;x=826516352;
#10;x=826616352;
#10;x=826716352;
#10;x=826816352;
#10;x=826916352;
#10;x=827016352;
#10;x=827116352;
#10;x=827216352;
#10;x=827316352;
#10;x=827416352;
#10;x=827516352;
#10;x=827616352;
#10;x=827716352;
#10;x=827816352;
#10;x=827916352;
#10;x=828016352;
#10;x=828116352;
#10;x=828216352;
#10;x=828316352;
#10;x=828416352;
#10;x=828516352;
#10;x=828616352;
#10;x=828716352;
#10;x=828816352;
#10;x=828916352;
#10;x=829016352;
#10;x=829116352;
#10;x=829216352;
#10;x=829316352;
#10;x=829416352;
#10;x=829516352;
#10;x=829616352;
#10;x=829716352;
#10;x=829816352;
#10;x=829916352;
#10;x=830016352;
#10;x=830116352;
#10;x=830216352;
#10;x=830316352;
#10;x=830416352;
#10;x=830516352;
#10;x=830616352;
#10;x=830716352;
#10;x=830816352;
#10;x=830916352;
#10;x=831016352;
#10;x=831116352;
#10;x=831216352;
#10;x=831316352;
#10;x=831416352;
#10;x=831516352;
#10;x=831616352;
#10;x=831716352;
#10;x=831816352;
#10;x=831916352;
#10;x=832016352;
#10;x=832116352;
#10;x=832216352;
#10;x=832316352;
#10;x=832416352;
#10;x=832516352;
#10;x=832616352;
#10;x=832716352;
#10;x=832816352;
#10;x=832916352;
#10;x=833016352;
#10;x=833116352;
#10;x=833216352;
#10;x=833316352;
#10;x=833416352;
#10;x=833516352;
#10;x=833616352;
#10;x=833716352;
#10;x=833816352;
#10;x=833916352;
#10;x=834016352;
#10;x=834116352;
#10;x=834216352;
#10;x=834316352;
#10;x=834416352;
#10;x=834516352;
#10;x=834616352;
#10;x=834716352;
#10;x=834816352;
#10;x=834916352;
#10;x=835016352;
#10;x=835116352;
#10;x=835216352;
#10;x=835316352;
#10;x=835416352;
#10;x=835516352;
#10;x=835616352;
#10;x=835716352;
#10;x=835816352;
#10;x=835916352;
#10;x=836016352;
#10;x=836116352;
#10;x=836216352;
#10;x=836316352;
#10;x=836416352;
#10;x=836516352;
#10;x=836616352;
#10;x=836716352;
#10;x=836816352;
#10;x=836916352;
#10;x=837016352;
#10;x=837116352;
#10;x=837216352;
#10;x=837316352;
#10;x=837416352;
#10;x=837516352;
#10;x=837616352;
#10;x=837716352;
#10;x=837816352;
#10;x=837916352;
#10;x=838016352;
#10;x=838116352;
#10;x=838216352;
#10;x=838316352;
#10;x=838416352;
#10;x=838516352;
#10;x=838616352;
#10;x=838716352;
#10;x=838816352;
#10;x=838916352;
#10;x=839016352;
#10;x=839116352;
#10;x=839216352;
#10;x=839316352;
#10;x=839416352;
#10;x=839516352;
#10;x=839616352;
#10;x=839716352;
#10;x=839816352;
#10;x=839916352;
#10;x=840016352;
#10;x=840116352;
#10;x=840216352;
#10;x=840316352;
#10;x=840416352;
#10;x=840516352;
#10;x=840616352;
#10;x=840716352;
#10;x=840816352;
#10;x=840916352;
#10;x=841016352;
#10;x=841116352;
#10;x=841216352;
#10;x=841316352;
#10;x=841416352;
#10;x=841516352;
#10;x=841616352;
#10;x=841716352;
#10;x=841816352;
#10;x=841916352;
#10;x=842016352;
#10;x=842116352;
#10;x=842216352;
#10;x=842316352;
#10;x=842416352;
#10;x=842516352;
#10;x=842616352;
#10;x=842716352;
#10;x=842816352;
#10;x=842916352;
#10;x=843016352;
#10;x=843116352;
#10;x=843216352;
#10;x=843316352;
#10;x=843416352;
#10;x=843516352;
#10;x=843616352;
#10;x=843716352;
#10;x=843816352;
#10;x=843916352;
#10;x=844016352;
#10;x=844116352;
#10;x=844216352;
#10;x=844316352;
#10;x=844416352;
#10;x=844516352;
#10;x=844616352;
#10;x=844716352;
#10;x=844816352;
#10;x=844916352;
#10;x=845016352;
#10;x=845116352;
#10;x=845216352;
#10;x=845316352;
#10;x=845416352;
#10;x=845516352;
#10;x=845616352;
#10;x=845716352;
#10;x=845816352;
#10;x=845916352;
#10;x=846016352;
#10;x=846116352;
#10;x=846216352;
#10;x=846316352;
#10;x=846416352;
#10;x=846516352;
#10;x=846616352;
#10;x=846716352;
#10;x=846816352;
#10;x=846916352;
#10;x=847016352;
#10;x=847116352;
#10;x=847216352;
#10;x=847316352;
#10;x=847416352;
#10;x=847516352;
#10;x=847616352;
#10;x=847716352;
#10;x=847816352;
#10;x=847916352;
#10;x=848016352;
#10;x=848116352;
#10;x=848216352;
#10;x=848316352;
#10;x=848416352;
#10;x=848516352;
#10;x=848616352;
#10;x=848716352;
#10;x=848816352;
#10;x=848916352;
#10;x=849016352;
#10;x=849116352;
#10;x=849216352;
#10;x=849316352;
#10;x=849416352;
#10;x=849516352;
#10;x=849616352;
#10;x=849716352;
#10;x=849816352;
#10;x=849916352;
#10;x=850016352;
#10;x=850116352;
#10;x=850216352;
#10;x=850316352;
#10;x=850416352;
#10;x=850516352;
#10;x=850616352;
#10;x=850716352;
#10;x=850816352;
#10;x=850916352;
#10;x=851016352;
#10;x=851116352;
#10;x=851216352;
#10;x=851316352;
#10;x=851416352;
#10;x=851516352;
#10;x=851616352;
#10;x=851716352;
#10;x=851816352;
#10;x=851916352;
#10;x=852016352;
#10;x=852116352;
#10;x=852216352;
#10;x=852316352;
#10;x=852416352;
#10;x=852516352;
#10;x=852616352;
#10;x=852716352;
#10;x=852816352;
#10;x=852916352;
#10;x=853016352;
#10;x=853116352;
#10;x=853216352;
#10;x=853316352;
#10;x=853416352;
#10;x=853516352;
#10;x=853616352;
#10;x=853716352;
#10;x=853816352;
#10;x=853916352;
#10;x=854016352;
#10;x=854116352;
#10;x=854216352;
#10;x=854316352;
#10;x=854416352;
#10;x=854516352;
#10;x=854616352;
#10;x=854716352;
#10;x=854816352;
#10;x=854916352;
#10;x=855016352;
#10;x=855116352;
#10;x=855216352;
#10;x=855316352;
#10;x=855416352;
#10;x=855516352;
#10;x=855616352;
#10;x=855716352;
#10;x=855816352;
#10;x=855916352;
#10;x=856016352;
#10;x=856116352;
#10;x=856216352;
#10;x=856316352;
#10;x=856416352;
#10;x=856516352;
#10;x=856616352;
#10;x=856716352;
#10;x=856816352;
#10;x=856916352;
#10;x=857016352;
#10;x=857116352;
#10;x=857216352;
#10;x=857316352;
#10;x=857416352;
#10;x=857516352;
#10;x=857616352;
#10;x=857716352;
#10;x=857816352;
#10;x=857916352;
#10;x=858016352;
#10;x=858116352;
#10;x=858216352;
#10;x=858316352;
#10;x=858416352;
#10;x=858516352;
#10;x=858616352;
#10;x=858716352;
#10;x=858816352;
#10;x=858916352;
#10;x=859016352;
#10;x=859116352;
#10;x=859216352;
#10;x=859316352;
#10;x=859416352;
#10;x=859516352;
#10;x=859616352;
#10;x=859716352;
#10;x=859816352;
#10;x=859916352;
#10;x=860016352;
#10;x=860116352;
#10;x=860216352;
#10;x=860316352;
#10;x=860416352;
#10;x=860516352;
#10;x=860616352;
#10;x=860716352;
#10;x=860816352;
#10;x=860916352;
#10;x=861016352;
#10;x=861116352;
#10;x=861216352;
#10;x=861316352;
#10;x=861416352;
#10;x=861516352;
#10;x=861616352;
#10;x=861716352;
#10;x=861816352;
#10;x=861916352;
#10;x=862016352;
#10;x=862116352;
#10;x=862216352;
#10;x=862316352;
#10;x=862416352;
#10;x=862516352;
#10;x=862616352;
#10;x=862716352;
#10;x=862816352;
#10;x=862916352;
#10;x=863016352;
#10;x=863116352;
#10;x=863216352;
#10;x=863316352;
#10;x=863416352;
#10;x=863516352;
#10;x=863616352;
#10;x=863716352;
#10;x=863816352;
#10;x=863916352;
#10;x=864016352;
#10;x=864116352;
#10;x=864216352;
#10;x=864316352;
#10;x=864416352;
#10;x=864516352;
#10;x=864616352;
#10;x=864716352;
#10;x=864816352;
#10;x=864916352;
#10;x=865016352;
#10;x=865116352;
#10;x=865216352;
#10;x=865316352;
#10;x=865416352;
#10;x=865516352;
#10;x=865616352;
#10;x=865716352;
#10;x=865816352;
#10;x=865916352;
#10;x=866016352;
#10;x=866116352;
#10;x=866216352;
#10;x=866316352;
#10;x=866416352;
#10;x=866516352;
#10;x=866616352;
#10;x=866716352;
#10;x=866816352;
#10;x=866916352;
#10;x=867016352;
#10;x=867116352;
#10;x=867216352;
#10;x=867316352;
#10;x=867416352;
#10;x=867516352;
#10;x=867616352;
#10;x=867716352;
#10;x=867816352;
#10;x=867916352;
#10;x=868016352;
#10;x=868116352;
#10;x=868216352;
#10;x=868316352;
#10;x=868416352;
#10;x=868516352;
#10;x=868616352;
#10;x=868716352;
#10;x=868816352;
#10;x=868916352;
#10;x=869016352;
#10;x=869116352;
#10;x=869216352;
#10;x=869316352;
#10;x=869416352;
#10;x=869516352;
#10;x=869616352;
#10;x=869716352;
#10;x=869816352;
#10;x=869916352;
#10;x=870016352;
#10;x=870116352;
#10;x=870216352;
#10;x=870316352;
#10;x=870416352;
#10;x=870516352;
#10;x=870616352;
#10;x=870716352;
#10;x=870816352;
#10;x=870916352;
#10;x=871016352;
#10;x=871116352;
#10;x=871216352;
#10;x=871316352;
#10;x=871416352;
#10;x=871516352;
#10;x=871616352;
#10;x=871716352;
#10;x=871816352;
#10;x=871916352;
#10;x=872016352;
#10;x=872116352;
#10;x=872216352;
#10;x=872316352;
#10;x=872416352;
#10;x=872516352;
#10;x=872616352;
#10;x=872716352;
#10;x=872816352;
#10;x=872916352;
#10;x=873016352;
#10;x=873116352;
#10;x=873216352;
#10;x=873316352;
#10;x=873416352;
#10;x=873516352;
#10;x=873616352;
#10;x=873716352;
#10;x=873816352;
#10;x=873916352;
#10;x=874016352;
#10;x=874116352;
#10;x=874216352;
#10;x=874316352;
#10;x=874416352;
#10;x=874516352;
#10;x=874616352;
#10;x=874716352;
#10;x=874816352;
#10;x=874916352;
#10;x=875016352;
#10;x=875116352;
#10;x=875216352;
#10;x=875316352;
#10;x=875416352;
#10;x=875516352;
#10;x=875616352;
#10;x=875716352;
#10;x=875816352;
#10;x=875916352;
#10;x=876016352;
#10;x=876116352;
#10;x=876216352;
#10;x=876316352;
#10;x=876416352;
#10;x=876516352;
#10;x=876616352;
#10;x=876716352;
#10;x=876816352;
#10;x=876916352;
#10;x=877016352;
#10;x=877116352;
#10;x=877216352;
#10;x=877316352;
#10;x=877416352;
#10;x=877516352;
#10;x=877616352;
#10;x=877716352;
#10;x=877816352;
#10;x=877916352;
#10;x=878016352;
#10;x=878116352;
#10;x=878216352;
#10;x=878316352;
#10;x=878416352;
#10;x=878516352;
#10;x=878616352;
#10;x=878716352;
#10;x=878816352;
#10;x=878916352;
#10;x=879016352;
#10;x=879116352;
#10;x=879216352;
#10;x=879316352;
#10;x=879416352;
#10;x=879516352;
#10;x=879616352;
#10;x=879716352;
#10;x=879816352;
#10;x=879916352;
#10;x=880016352;
#10;x=880116352;
#10;x=880216352;
#10;x=880316352;
#10;x=880416352;
#10;x=880516352;
#10;x=880616352;
#10;x=880716352;
#10;x=880816352;
#10;x=880916352;
#10;x=881016352;
#10;x=881116352;
#10;x=881216352;
#10;x=881316352;
#10;x=881416352;
#10;x=881516352;
#10;x=881616352;
#10;x=881716352;
#10;x=881816352;
#10;x=881916352;
#10;x=882016352;
#10;x=882116352;
#10;x=882216352;
#10;x=882316352;
#10;x=882416352;
#10;x=882516352;
#10;x=882616352;
#10;x=882716352;
#10;x=882816352;
#10;x=882916352;
#10;x=883016352;
#10;x=883116352;
#10;x=883216352;
#10;x=883316352;
#10;x=883416352;
#10;x=883516352;
#10;x=883616352;
#10;x=883716352;
#10;x=883816352;
#10;x=883916352;
#10;x=884016352;
#10;x=884116352;
#10;x=884216352;
#10;x=884316352;
#10;x=884416352;
#10;x=884516352;
#10;x=884616352;
#10;x=884716352;
#10;x=884816352;
#10;x=884916352;
#10;x=885016352;
#10;x=885116352;
#10;x=885216352;
#10;x=885316352;
#10;x=885416352;
#10;x=885516352;
#10;x=885616352;
#10;x=885716352;
#10;x=885816352;
#10;x=885916352;
#10;x=886016352;
#10;x=886116352;
#10;x=886216352;
#10;x=886316352;
#10;x=886416352;
#10;x=886516352;
#10;x=886616352;
#10;x=886716352;
#10;x=886816352;
#10;x=886916352;
#10;x=887016352;
#10;x=887116352;
#10;x=887216352;
#10;x=887316352;
#10;x=887416352;
#10;x=887516352;
#10;x=887616352;
#10;x=887716352;
#10;x=887816352;
#10;x=887916352;
#10;x=888016352;
#10;x=888116352;
#10;x=888216352;
#10;x=888316352;
#10;x=888416352;
#10;x=888516352;
#10;x=888616352;
#10;x=888716352;
#10;x=888816352;
#10;x=888916352;
#10;x=889016352;
#10;x=889116352;
#10;x=889216352;
#10;x=889316352;
#10;x=889416352;
#10;x=889516352;
#10;x=889616352;
#10;x=889716352;
#10;x=889816352;
#10;x=889916352;
#10;x=890016352;
#10;x=890116352;
#10;x=890216352;
#10;x=890316352;
#10;x=890416352;
#10;x=890516352;
#10;x=890616352;
#10;x=890716352;
#10;x=890816352;
#10;x=890916352;
#10;x=891016352;
#10;x=891116352;
#10;x=891216352;
#10;x=891316352;
#10;x=891416352;
#10;x=891516352;
#10;x=891616352;
#10;x=891716352;
#10;x=891816352;
#10;x=891916352;
#10;x=892016352;
#10;x=892116352;
#10;x=892216352;
#10;x=892316352;
#10;x=892416352;
#10;x=892516352;
#10;x=892616352;
#10;x=892716352;
#10;x=892816352;
#10;x=892916352;
#10;x=893016352;
#10;x=893116352;
#10;x=893216352;
#10;x=893316352;
#10;x=893416352;
#10;x=893516352;
#10;x=893616352;
#10;x=893716352;
#10;x=893816352;
#10;x=893916352;
#10;x=894016352;
#10;x=894116352;
#10;x=894216352;
#10;x=894316352;
#10;x=894416352;
#10;x=894516352;
#10;x=894616352;
#10;x=894716352;
#10;x=894816352;
#10;x=894916352;
#10;x=895016352;
#10;x=895116352;
#10;x=895216352;
#10;x=895316352;
#10;x=895416352;
#10;x=895516352;
#10;x=895616352;
#10;x=895716352;
#10;x=895816352;
#10;x=895916352;
#10;x=896016352;
#10;x=896116352;
#10;x=896216352;
#10;x=896316352;
#10;x=896416352;
#10;x=896516352;
#10;x=896616352;
#10;x=896716352;
#10;x=896816352;
#10;x=896916352;
#10;x=897016352;
#10;x=897116352;
#10;x=897216352;
#10;x=897316352;
#10;x=897416352;
#10;x=897516352;
#10;x=897616352;
#10;x=897716352;
#10;x=897816352;
#10;x=897916352;
#10;x=898016352;
#10;x=898116352;
#10;x=898216352;
#10;x=898316352;
#10;x=898416352;
#10;x=898516352;
#10;x=898616352;
#10;x=898716352;
#10;x=898816352;
#10;x=898916352;
#10;x=899016352;
#10;x=899116352;
#10;x=899216352;
#10;x=899316352;
#10;x=899416352;
#10;x=899516352;
#10;x=899616352;
#10;x=899716352;
#10;x=899816352;
#10;x=899916352;
#10;x=900016352;
#10;x=900116352;
#10;x=900216352;
#10;x=900316352;
#10;x=900416352;
#10;x=900516352;
#10;x=900616352;
#10;x=900716352;
#10;x=900816352;
#10;x=900916352;
#10;x=901016352;
#10;x=901116352;
#10;x=901216352;
#10;x=901316352;
#10;x=901416352;
#10;x=901516352;
#10;x=901616352;
#10;x=901716352;
#10;x=901816352;
#10;x=901916352;
#10;x=902016352;
#10;x=902116352;
#10;x=902216352;
#10;x=902316352;
#10;x=902416352;
#10;x=902516352;
#10;x=902616352;
#10;x=902716352;
#10;x=902816352;
#10;x=902916352;
#10;x=903016352;
#10;x=903116352;
#10;x=903216352;
#10;x=903316352;
#10;x=903416352;
#10;x=903516352;
#10;x=903616352;
#10;x=903716352;
#10;x=903816352;
#10;x=903916352;
#10;x=904016352;
#10;x=904116352;
#10;x=904216352;
#10;x=904316352;
#10;x=904416352;
#10;x=904516352;
#10;x=904616352;
#10;x=904716352;
#10;x=904816352;
#10;x=904916352;
#10;x=905016352;
#10;x=905116352;
#10;x=905216352;
#10;x=905316352;
#10;x=905416352;
#10;x=905516352;
#10;x=905616352;
#10;x=905716352;
#10;x=905816352;
#10;x=905916352;
#10;x=906016352;
#10;x=906116352;
#10;x=906216352;
#10;x=906316352;
#10;x=906416352;
#10;x=906516352;
#10;x=906616352;
#10;x=906716352;
#10;x=906816352;
#10;x=906916352;
#10;x=907016352;
#10;x=907116352;
#10;x=907216352;
#10;x=907316352;
#10;x=907416352;
#10;x=907516352;
#10;x=907616352;
#10;x=907716352;
#10;x=907816352;
#10;x=907916352;
#10;x=908016352;
#10;x=908116352;
#10;x=908216352;
#10;x=908316352;
#10;x=908416352;
#10;x=908516352;
#10;x=908616352;
#10;x=908716352;
#10;x=908816352;
#10;x=908916352;
#10;x=909016352;
#10;x=909116352;
#10;x=909216352;
#10;x=909316352;
#10;x=909416352;
#10;x=909516352;
#10;x=909616352;
#10;x=909716352;
#10;x=909816352;
#10;x=909916352;
#10;x=910016352;
#10;x=910116352;
#10;x=910216352;
#10;x=910316352;
#10;x=910416352;
#10;x=910516352;
#10;x=910616352;
#10;x=910716352;
#10;x=910816352;
#10;x=910916352;
#10;x=911016352;
#10;x=911116352;
#10;x=911216352;
#10;x=911316352;
#10;x=911416352;
#10;x=911516352;
#10;x=911616352;
#10;x=911716352;
#10;x=911816352;
#10;x=911916352;
#10;x=912016352;
#10;x=912116352;
#10;x=912216352;
#10;x=912316352;
#10;x=912416352;
#10;x=912516352;
#10;x=912616352;
#10;x=912716352;
#10;x=912816352;
#10;x=912916352;
#10;x=913016352;
#10;x=913116352;
#10;x=913216352;
#10;x=913316352;
#10;x=913416352;
#10;x=913516352;
#10;x=913616352;
#10;x=913716352;
#10;x=913816352;
#10;x=913916352;
#10;x=914016352;
#10;x=914116352;
#10;x=914216352;
#10;x=914316352;
#10;x=914416352;
#10;x=914516352;
#10;x=914616352;
#10;x=914716352;
#10;x=914816352;
#10;x=914916352;
#10;x=915016352;
#10;x=915116352;
#10;x=915216352;
#10;x=915316352;
#10;x=915416352;
#10;x=915516352;
#10;x=915616352;
#10;x=915716352;
#10;x=915816352;
#10;x=915916352;
#10;x=916016352;
#10;x=916116352;
#10;x=916216352;
#10;x=916316352;
#10;x=916416352;
#10;x=916516352;
#10;x=916616352;
#10;x=916716352;
#10;x=916816352;
#10;x=916916352;
#10;x=917016352;
#10;x=917116352;
#10;x=917216352;
#10;x=917316352;
#10;x=917416352;
#10;x=917516352;
#10;x=917616352;
#10;x=917716352;
#10;x=917816352;
#10;x=917916352;
#10;x=918016352;
#10;x=918116352;
#10;x=918216352;
#10;x=918316352;
#10;x=918416352;
#10;x=918516352;
#10;x=918616352;
#10;x=918716352;
#10;x=918816352;
#10;x=918916352;
#10;x=919016352;
#10;x=919116352;
#10;x=919216352;
#10;x=919316352;
#10;x=919416352;
#10;x=919516352;
#10;x=919616352;
#10;x=919716352;
#10;x=919816352;
#10;x=919916352;
#10;x=920016352;
#10;x=920116352;
#10;x=920216352;
#10;x=920316352;
#10;x=920416352;
#10;x=920516352;
#10;x=920616352;
#10;x=920716352;
#10;x=920816352;
#10;x=920916352;
#10;x=921016352;
#10;x=921116352;
#10;x=921216352;
#10;x=921316352;
#10;x=921416352;
#10;x=921516352;
#10;x=921616352;
#10;x=921716352;
#10;x=921816352;
#10;x=921916352;
#10;x=922016352;
#10;x=922116352;
#10;x=922216352;
#10;x=922316352;
#10;x=922416352;
#10;x=922516352;
#10;x=922616352;
#10;x=922716352;
#10;x=922816352;
#10;x=922916352;
#10;x=923016352;
#10;x=923116352;
#10;x=923216352;
#10;x=923316352;
#10;x=923416352;
#10;x=923516352;
#10;x=923616352;
#10;x=923716352;
#10;x=923816352;
#10;x=923916352;
#10;x=924016352;
#10;x=924116352;
#10;x=924216352;
#10;x=924316352;
#10;x=924416352;
#10;x=924516352;
#10;x=924616352;
#10;x=924716352;
#10;x=924816352;
#10;x=924916352;
#10;x=925016352;
#10;x=925116352;
#10;x=925216352;
#10;x=925316352;
#10;x=925416352;
#10;x=925516352;
#10;x=925616352;
#10;x=925716352;
#10;x=925816352;
#10;x=925916352;
#10;x=926016352;
#10;x=926116352;
#10;x=926216352;
#10;x=926316352;
#10;x=926416352;
#10;x=926516352;
#10;x=926616352;
#10;x=926716352;
#10;x=926816352;
#10;x=926916352;
#10;x=927016352;
#10;x=927116352;
#10;x=927216352;
#10;x=927316352;
#10;x=927416352;
#10;x=927516352;
#10;x=927616352;
#10;x=927716352;
#10;x=927816352;
#10;x=927916352;
#10;x=928016352;
#10;x=928116352;
#10;x=928216352;
#10;x=928316352;
#10;x=928416352;
#10;x=928516352;
#10;x=928616352;
#10;x=928716352;
#10;x=928816352;
#10;x=928916352;
#10;x=929016352;
#10;x=929116352;
#10;x=929216352;
#10;x=929316352;
#10;x=929416352;
#10;x=929516352;
#10;x=929616352;
#10;x=929716352;
#10;x=929816352;
#10;x=929916352;
#10;x=930016352;
#10;x=930116352;
#10;x=930216352;
#10;x=930316352;
#10;x=930416352;
#10;x=930516352;
#10;x=930616352;
#10;x=930716352;
#10;x=930816352;
#10;x=930916352;
#10;x=931016352;
#10;x=931116352;
#10;x=931216352;
#10;x=931316352;
#10;x=931416352;
#10;x=931516352;
#10;x=931616352;
#10;x=931716352;
#10;x=931816352;
#10;x=931916352;
#10;x=932016352;
#10;x=932116352;
#10;x=932216352;
#10;x=932316352;
#10;x=932416352;
#10;x=932516352;
#10;x=932616352;
#10;x=932716352;
#10;x=932816352;
#10;x=932916352;
#10;x=933016352;
#10;x=933116352;
#10;x=933216352;
#10;x=933316352;
#10;x=933416352;
#10;x=933516352;
#10;x=933616352;
#10;x=933716352;
#10;x=933816352;
#10;x=933916352;
#10;x=934016352;
#10;x=934116352;
#10;x=934216352;
#10;x=934316352;
#10;x=934416352;
#10;x=934516352;
#10;x=934616352;
#10;x=934716352;
#10;x=934816352;
#10;x=934916352;
#10;x=935016352;
#10;x=935116352;
#10;x=935216352;
#10;x=935316352;
#10;x=935416352;
#10;x=935516352;
#10;x=935616352;
#10;x=935716352;
#10;x=935816352;
#10;x=935916352;
#10;x=936016352;
#10;x=936116352;
#10;x=936216352;
#10;x=936316352;
#10;x=936416352;
#10;x=936516352;
#10;x=936616352;
#10;x=936716352;
#10;x=936816352;
#10;x=936916352;
#10;x=937016352;
#10;x=937116352;
#10;x=937216352;
#10;x=937316352;
#10;x=937416352;
#10;x=937516352;
#10;x=937616352;
#10;x=937716352;
#10;x=937816352;
#10;x=937916352;
#10;x=938016352;
#10;x=938116352;
#10;x=938216352;
#10;x=938316352;
#10;x=938416352;
#10;x=938516352;
#10;x=938616352;
#10;x=938716352;
#10;x=938816352;
#10;x=938916352;
#10;x=939016352;
#10;x=939116352;
#10;x=939216352;
#10;x=939316352;
#10;x=939416352;
#10;x=939516352;
#10;x=939616352;
#10;x=939716352;
#10;x=939816352;
#10;x=939916352;
#10;x=940016352;
#10;x=940116352;
#10;x=940216352;
#10;x=940316352;
#10;x=940416352;
#10;x=940516352;
#10;x=940616352;
#10;x=940716352;
#10;x=940816352;
#10;x=940916352;
#10;x=941016352;
#10;x=941116352;
#10;x=941216352;
#10;x=941316352;
#10;x=941416352;
#10;x=941516352;
#10;x=941616352;
#10;x=941716352;
#10;x=941816352;
#10;x=941916352;
#10;x=942016352;
#10;x=942116352;
#10;x=942216352;
#10;x=942316352;
#10;x=942416352;
#10;x=942516352;
#10;x=942616352;
#10;x=942716352;
#10;x=942816352;
#10;x=942916352;
#10;x=943016352;
#10;x=943116352;
#10;x=943216352;
#10;x=943316352;
#10;x=943416352;
#10;x=943516352;
#10;x=943616352;
#10;x=943716352;
#10;x=943816352;
#10;x=943916352;
#10;x=944016352;
#10;x=944116352;
#10;x=944216352;
#10;x=944316352;
#10;x=944416352;
#10;x=944516352;
#10;x=944616352;
#10;x=944716352;
#10;x=944816352;
#10;x=944916352;
#10;x=945016352;
#10;x=945116352;
#10;x=945216352;
#10;x=945316352;
#10;x=945416352;
#10;x=945516352;
#10;x=945616352;
#10;x=945716352;
#10;x=945816352;
#10;x=945916352;
#10;x=946016352;
#10;x=946116352;
#10;x=946216352;
#10;x=946316352;
#10;x=946416352;
#10;x=946516352;
#10;x=946616352;
#10;x=946716352;
#10;x=946816352;
#10;x=946916352;
#10;x=947016352;
#10;x=947116352;
#10;x=947216352;
#10;x=947316352;
#10;x=947416352;
#10;x=947516352;
#10;x=947616352;
#10;x=947716352;
#10;x=947816352;
#10;x=947916352;
#10;x=948016352;
#10;x=948116352;
#10;x=948216352;
#10;x=948316352;
#10;x=948416352;
#10;x=948516352;
#10;x=948616352;
#10;x=948716352;
#10;x=948816352;
#10;x=948916352;
#10;x=949016352;
#10;x=949116352;
#10;x=949216352;
#10;x=949316352;
#10;x=949416352;
#10;x=949516352;
#10;x=949616352;
#10;x=949716352;
#10;x=949816352;
#10;x=949916352;
#10;x=950016352;
#10;x=950116352;
#10;x=950216352;
#10;x=950316352;
#10;x=950416352;
#10;x=950516352;
#10;x=950616352;
#10;x=950716352;
#10;x=950816352;
#10;x=950916352;
#10;x=951016352;
#10;x=951116352;
#10;x=951216352;
#10;x=951316352;
#10;x=951416352;
#10;x=951516352;
#10;x=951616352;
#10;x=951716352;
#10;x=951816352;
#10;x=951916352;
#10;x=952016352;
#10;x=952116352;
#10;x=952216352;
#10;x=952316352;
#10;x=952416352;
#10;x=952516352;
#10;x=952616352;
#10;x=952716352;
#10;x=952816352;
#10;x=952916352;
#10;x=953016352;
#10;x=953116352;
#10;x=953216352;
#10;x=953316352;
#10;x=953416352;
#10;x=953516352;
#10;x=953616352;
#10;x=953716352;
#10;x=953816352;
#10;x=953916352;
#10;x=954016352;
#10;x=954116352;
#10;x=954216352;
#10;x=954316352;
#10;x=954416352;
#10;x=954516352;
#10;x=954616352;
#10;x=954716352;
#10;x=954816352;
#10;x=954916352;
#10;x=955016352;
#10;x=955116352;
#10;x=955216352;
#10;x=955316352;
#10;x=955416352;
#10;x=955516352;
#10;x=955616352;
#10;x=955716352;
#10;x=955816352;
#10;x=955916352;
#10;x=956016352;
#10;x=956116352;
#10;x=956216352;
#10;x=956316352;
#10;x=956416352;
#10;x=956516352;
#10;x=956616352;
#10;x=956716352;
#10;x=956816352;
#10;x=956916352;
#10;x=957016352;
#10;x=957116352;
#10;x=957216352;
#10;x=957316352;
#10;x=957416352;
#10;x=957516352;
#10;x=957616352;
#10;x=957716352;
#10;x=957816352;
#10;x=957916352;
#10;x=958016352;
#10;x=958116352;
#10;x=958216352;
#10;x=958316352;
#10;x=958416352;
#10;x=958516352;
#10;x=958616352;
#10;x=958716352;
#10;x=958816352;
#10;x=958916352;
#10;x=959016352;
#10;x=959116352;
#10;x=959216352;
#10;x=959316352;
#10;x=959416352;
#10;x=959516352;
#10;x=959616352;
#10;x=959716352;
#10;x=959816352;
#10;x=959916352;
#10;x=960016352;
#10;x=960116352;
#10;x=960216352;
#10;x=960316352;
#10;x=960416352;
#10;x=960516352;
#10;x=960616352;
#10;x=960716352;
#10;x=960816352;
#10;x=960916352;
#10;x=961016352;
#10;x=961116352;
#10;x=961216352;
#10;x=961316352;
#10;x=961416352;
#10;x=961516352;
#10;x=961616352;
#10;x=961716352;
#10;x=961816352;
#10;x=961916352;
#10;x=962016352;
#10;x=962116352;
#10;x=962216352;
#10;x=962316352;
#10;x=962416352;
#10;x=962516352;
#10;x=962616352;
#10;x=962716352;
#10;x=962816352;
#10;x=962916352;
#10;x=963016352;
#10;x=963116352;
#10;x=963216352;
#10;x=963316352;
#10;x=963416352;
#10;x=963516352;
#10;x=963616352;
#10;x=963716352;
#10;x=963816352;
#10;x=963916352;
#10;x=964016352;
#10;x=964116352;
#10;x=964216352;
#10;x=964316352;
#10;x=964416352;
#10;x=964516352;
#10;x=964616352;
#10;x=964716352;
#10;x=964816352;
#10;x=964916352;
#10;x=965016352;
#10;x=965116352;
#10;x=965216352;
#10;x=965316352;
#10;x=965416352;
#10;x=965516352;
#10;x=965616352;
#10;x=965716352;
#10;x=965816352;
#10;x=965916352;
#10;x=966016352;
#10;x=966116352;
#10;x=966216352;
#10;x=966316352;
#10;x=966416352;
#10;x=966516352;
#10;x=966616352;
#10;x=966716352;
#10;x=966816352;
#10;x=966916352;
#10;x=967016352;
#10;x=967116352;
#10;x=967216352;
#10;x=967316352;
#10;x=967416352;
#10;x=967516352;
#10;x=967616352;
#10;x=967716352;
#10;x=967816352;
#10;x=967916352;
#10;x=968016352;
#10;x=968116352;
#10;x=968216352;
#10;x=968316352;
#10;x=968416352;
#10;x=968516352;
#10;x=968616352;
#10;x=968716352;
#10;x=968816352;
#10;x=968916352;
#10;x=969016352;
#10;x=969116352;
#10;x=969216352;
#10;x=969316352;
#10;x=969416352;
#10;x=969516352;
#10;x=969616352;
#10;x=969716352;
#10;x=969816352;
#10;x=969916352;
#10;x=970016352;
#10;x=970116352;
#10;x=970216352;
#10;x=970316352;
#10;x=970416352;
#10;x=970516352;
#10;x=970616352;
#10;x=970716352;
#10;x=970816352;
#10;x=970916352;
#10;x=971016352;
#10;x=971116352;
#10;x=971216352;
#10;x=971316352;
#10;x=971416352;
#10;x=971516352;
#10;x=971616352;
#10;x=971716352;
#10;x=971816352;
#10;x=971916352;
#10;x=972016352;
#10;x=972116352;
#10;x=972216352;
#10;x=972316352;
#10;x=972416352;
#10;x=972516352;
#10;x=972616352;
#10;x=972716352;
#10;x=972816352;
#10;x=972916352;
#10;x=973016352;
#10;x=973116352;
#10;x=973216352;
#10;x=973316352;
#10;x=973416352;
#10;x=973516352;
#10;x=973616352;
#10;x=973716352;
#10;x=973816352;
#10;x=973916352;
#10;x=974016352;
#10;x=974116352;
#10;x=974216352;
#10;x=974316352;
#10;x=974416352;
#10;x=974516352;
#10;x=974616352;
#10;x=974716352;
#10;x=974816352;
#10;x=974916352;
#10;x=975016352;
#10;x=975116352;
#10;x=975216352;
#10;x=975316352;
#10;x=975416352;
#10;x=975516352;
#10;x=975616352;
#10;x=975716352;
#10;x=975816352;
#10;x=975916352;
#10;x=976016352;
#10;x=976116352;
#10;x=976216352;
#10;x=976316352;
#10;x=976416352;
#10;x=976516352;
#10;x=976616352;
#10;x=976716352;
#10;x=976816352;
#10;x=976916352;
#10;x=977016352;
#10;x=977116352;
#10;x=977216352;
#10;x=977316352;
#10;x=977416352;
#10;x=977516352;
#10;x=977616352;
#10;x=977716352;
#10;x=977816352;
#10;x=977916352;
#10;x=978016352;
#10;x=978116352;
#10;x=978216352;
#10;x=978316352;
#10;x=978416352;
#10;x=978516352;
#10;x=978616352;
#10;x=978716352;
#10;x=978816352;
#10;x=978916352;
#10;x=979016352;
#10;x=979116352;
#10;x=979216352;
#10;x=979316352;
#10;x=979416352;
#10;x=979516352;
#10;x=979616352;
#10;x=979716352;
#10;x=979816352;
#10;x=979916352;
#10;x=980016352;
#10;x=980116352;
#10;x=980216352;
#10;x=980316352;
#10;x=980416352;
#10;x=980516352;
#10;x=980616352;
#10;x=980716352;
#10;x=980816352;
#10;x=980916352;
#10;x=981016352;
#10;x=981116352;
#10;x=981216352;
#10;x=981316352;
#10;x=981416352;
#10;x=981516352;
#10;x=981616352;
#10;x=981716352;
#10;x=981816352;
#10;x=981916352;
#10;x=982016352;
#10;x=982116352;
#10;x=982216352;
#10;x=982316352;
#10;x=982416352;
#10;x=982516352;
#10;x=982616352;
#10;x=982716352;
#10;x=982816352;
#10;x=982916352;
#10;x=983016352;
#10;x=983116352;
#10;x=983216352;
#10;x=983316352;
#10;x=983416352;
#10;x=983516352;
#10;x=983616352;
#10;x=983716352;
#10;x=983816352;
#10;x=983916352;
#10;x=984016352;
#10;x=984116352;
#10;x=984216352;
#10;x=984316352;
#10;x=984416352;
#10;x=984516352;
#10;x=984616352;
#10;x=984716352;
#10;x=984816352;
#10;x=984916352;
#10;x=985016352;
#10;x=985116352;
#10;x=985216352;
#10;x=985316352;
#10;x=985416352;
#10;x=985516352;
#10;x=985616352;
#10;x=985716352;
#10;x=985816352;
#10;x=985916352;
#10;x=986016352;
#10;x=986116352;
#10;x=986216352;
#10;x=986316352;
#10;x=986416352;
#10;x=986516352;
#10;x=986616352;
#10;x=986716352;
#10;x=986816352;
#10;x=986916352;
#10;x=987016352;
#10;x=987116352;
#10;x=987216352;
#10;x=987316352;
#10;x=987416352;
#10;x=987516352;
#10;x=987616352;
#10;x=987716352;
#10;x=987816352;
#10;x=987916352;
#10;x=988016352;
#10;x=988116352;
#10;x=988216352;
#10;x=988316352;
#10;x=988416352;
#10;x=988516352;
#10;x=988616352;
#10;x=988716352;
#10;x=988816352;
#10;x=988916352;
#10;x=989016352;
#10;x=989116352;
#10;x=989216352;
#10;x=989316352;
#10;x=989416352;
#10;x=989516352;
#10;x=989616352;
#10;x=989716352;
#10;x=989816352;
#10;x=989916352;
#10;x=990016352;
#10;x=990116352;
#10;x=990216352;
#10;x=990316352;
#10;x=990416352;
#10;x=990516352;
#10;x=990616352;
#10;x=990716352;
#10;x=990816352;
#10;x=990916352;
#10;x=991016352;
#10;x=991116352;
#10;x=991216352;
#10;x=991316352;
#10;x=991416352;
#10;x=991516352;
#10;x=991616352;
#10;x=991716352;
#10;x=991816352;
#10;x=991916352;
#10;x=992016352;
#10;x=992116352;
#10;x=992216352;
#10;x=992316352;
#10;x=992416352;
#10;x=992516352;
#10;x=992616352;
#10;x=992716352;
#10;x=992816352;
#10;x=992916352;
#10;x=993016352;
#10;x=993116352;
#10;x=993216352;
#10;x=993316352;
#10;x=993416352;
#10;x=993516352;
#10;x=993616352;
#10;x=993716352;
#10;x=993816352;
#10;x=993916352;
#10;x=994016352;
#10;x=994116352;
#10;x=994216352;
#10;x=994316352;
#10;x=994416352;
#10;x=994516352;
#10;x=994616352;
#10;x=994716352;
#10;x=994816352;
#10;x=994916352;
#10;x=995016352;
#10;x=995116352;
#10;x=995216352;
#10;x=995316352;
#10;x=995416352;
#10;x=995516352;
#10;x=995616352;
#10;x=995716352;
#10;x=995816352;
#10;x=995916352;
#10;x=996016352;
#10;x=996116352;
#10;x=996216352;
#10;x=996316352;
#10;x=996416352;
#10;x=996516352;
#10;x=996616352;
#10;x=996716352;
#10;x=996816352;
#10;x=996916352;
#10;x=997016352;
#10;x=997116352;
#10;x=997216352;
#10;x=997316352;
#10;x=997416352;
#10;x=997516352;
#10;x=997616352;
#10;x=997716352;
#10;x=997816352;
#10;x=997916352;
#10;x=998016352;
#10;x=998116352;
#10;x=998216352;
#10;x=998316352;
#10;x=998416352;
#10;x=998516352;
#10;x=998616352;
#10;x=998716352;
#10;x=998816352;
#10;x=998916352;
#10;x=999016352;
#10;x=999116352;
#10;x=999216352;
#10;x=999316352;
#10;x=999416352;
#10;x=999516352;
#10;x=999616352;
#10;x=999716352;
#10;x=999816352;
#10;x=999916352;
#10;x=1000016352;
#10;x=1001016352;
#10;x=1002016352;
#10;x=1003016352;
#10;x=1004016352;
#10;x=1005016352;
#10;x=1006016352;
#10;x=1007016352;
#10;x=1008016352;
#10;x=1009016352;
#10;x=1010016352;
#10;x=1011016352;
#10;x=1012016352;
#10;x=1013016352;
#10;x=1014016352;
#10;x=1015016352;
#10;x=1016016352;
#10;x=1017016352;
#10;x=1018016352;
#10;x=1019016352;
#10;x=1020016352;
#10;x=1021016352;
#10;x=1022016352;
#10;x=1023016352;
#10;x=1024016352;
#10;x=1025016352;
#10;x=1026016352;
#10;x=1027016352;
#10;x=1028016352;
#10;x=1029016352;
#10;x=1030016352;
#10;x=1031016352;
#10;x=1032016352;
#10;x=1033016352;
#10;x=1034016352;
#10;x=1035016352;
#10;x=1036016352;
#10;x=1037016352;
#10;x=1038016352;
#10;x=1039016352;
#10;x=1040016352;
#10;x=1041016352;
#10;x=1042016352;
#10;x=1043016352;
#10;x=1044016352;
#10;x=1045016352;
#10;x=1046016352;
#10;x=1047016352;
#10;x=1048016352;
#10;x=1049016352;
#10;x=1050016352;
#10;x=1051016352;
#10;x=1052016352;
#10;x=1053016352;
#10;x=1054016352;
#10;x=1055016352;
#10;x=1056016352;
#10;x=1057016352;
#10;x=1058016352;
#10;x=1059016352;
#10;x=1060016352;
#10;x=1061016352;
#10;x=1062016352;
#10;x=1063016352;
#10;x=1064016352;
#10;x=1065016352;
#10;x=1066016352;
#10;x=1067016352;
#10;x=1068016352;
#10;x=1069016352;
#10;x=1070016352;
#10;x=1071016352;
#10;x=1072016352;
#10;x=1073016352;
#10;x=1074016352;
#10;x=1075016352;
#10;x=1076016352;
#10;x=1077016352;
#10;x=1078016352;
#10;x=1079016352;
#10;x=1080016352;
#10;x=1081016352;
#10;x=1082016352;
#10;x=1083016352;
#10;x=1084016352;
#10;x=1085016352;
#10;x=1086016352;
#10;x=1087016352;
#10;x=1088016352;
#10;x=1089016352;
#10;x=1090016352;
#10;x=1091016352;
#10;x=1092016352;
#10;x=1093016352;
#10;x=1094016352;
#10;x=1095016352;
#10;x=1096016352;
#10;x=1097016352;
#10;x=1098016352;
#10;x=1099016352;
#10;x=1100016352;
#10;x=1101016352;
#10;x=1102016352;
#10;x=1103016352;
#10;x=1104016352;
#10;x=1105016352;
#10;x=1106016352;
#10;x=1107016352;
#10;x=1108016352;
#10;x=1109016352;
#10;x=1110016352;
#10;x=1111016352;
#10;x=1112016352;
#10;x=1113016352;
#10;x=1114016352;
#10;x=1115016352;
#10;x=1116016352;
#10;x=1117016352;
#10;x=1118016352;
#10;x=1119016352;
#10;x=1120016352;
#10;x=1121016352;
#10;x=1122016352;
#10;x=1123016352;
#10;x=1124016352;
#10;x=1125016352;
#10;x=1126016352;
#10;x=1127016352;
#10;x=1128016352;
#10;x=1129016352;
#10;x=1130016352;
#10;x=1131016352;
#10;x=1132016352;
#10;x=1133016352;
#10;x=1134016352;
#10;x=1135016352;
#10;x=1136016352;
#10;x=1137016352;
#10;x=1138016352;
#10;x=1139016352;
#10;x=1140016352;
#10;x=1141016352;
#10;x=1142016352;
#10;x=1143016352;
#10;x=1144016352;
#10;x=1145016352;
#10;x=1146016352;
#10;x=1147016352;
#10;x=1148016352;
#10;x=1149016352;
#10;x=1150016352;
#10;x=1151016352;
#10;x=1152016352;
#10;x=1153016352;
#10;x=1154016352;
#10;x=1155016352;
#10;x=1156016352;
#10;x=1157016352;
#10;x=1158016352;
#10;x=1159016352;
#10;x=1160016352;
#10;x=1161016352;
#10;x=1162016352;
#10;x=1163016352;
#10;x=1164016352;
#10;x=1165016352;
#10;x=1166016352;
#10;x=1167016352;
#10;x=1168016352;
#10;x=1169016352;
#10;x=1170016352;
#10;x=1171016352;
#10;x=1172016352;
#10;x=1173016352;
#10;x=1174016352;
#10;x=1175016352;
#10;x=1176016352;
#10;x=1177016352;
#10;x=1178016352;
#10;x=1179016352;
#10;x=1180016352;
#10;x=1181016352;
#10;x=1182016352;
#10;x=1183016352;
#10;x=1184016352;
#10;x=1185016352;
#10;x=1186016352;
#10;x=1187016352;
#10;x=1188016352;
#10;x=1189016352;
#10;x=1190016352;
#10;x=1191016352;
#10;x=1192016352;
#10;x=1193016352;
#10;x=1194016352;
#10;x=1195016352;
#10;x=1196016352;
#10;x=1197016352;
#10;x=1198016352;
#10;x=1199016352;
#10;x=1200016352;
#10;x=1201016352;
#10;x=1202016352;
#10;x=1203016352;
#10;x=1204016352;
#10;x=1205016352;
#10;x=1206016352;
#10;x=1207016352;
#10;x=1208016352;
#10;x=1209016352;
#10;x=1210016352;
#10;x=1211016352;
#10;x=1212016352;
#10;x=1213016352;
#10;x=1214016352;
#10;x=1215016352;
#10;x=1216016352;
#10;x=1217016352;
#10;x=1218016352;
#10;x=1219016352;
#10;x=1220016352;
#10;x=1221016352;
#10;x=1222016352;
#10;x=1223016352;
#10;x=1224016352;
#10;x=1225016352;
#10;x=1226016352;
#10;x=1227016352;
#10;x=1228016352;
#10;x=1229016352;
#10;x=1230016352;
#10;x=1231016352;
#10;x=1232016352;
#10;x=1233016352;
#10;x=1234016352;
#10;x=1235016352;
#10;x=1236016352;
#10;x=1237016352;
#10;x=1238016352;
#10;x=1239016352;
#10;x=1240016352;
#10;x=1241016352;
#10;x=1242016352;
#10;x=1243016352;
#10;x=1244016352;
#10;x=1245016352;
#10;x=1246016352;
#10;x=1247016352;
#10;x=1248016352;
#10;x=1249016352;
#10;x=1250016352;
#10;x=1251016352;
#10;x=1252016352;
#10;x=1253016352;
#10;x=1254016352;
#10;x=1255016352;
#10;x=1256016352;
#10;x=1257016352;
#10;x=1258016352;
#10;x=1259016352;
#10;x=1260016352;
#10;x=1261016352;
#10;x=1262016352;
#10;x=1263016352;
#10;x=1264016352;
#10;x=1265016352;
#10;x=1266016352;
#10;x=1267016352;
#10;x=1268016352;
#10;x=1269016352;
#10;x=1270016352;
#10;x=1271016352;
#10;x=1272016352;
#10;x=1273016352;
#10;x=1274016352;
#10;x=1275016352;
#10;x=1276016352;
#10;x=1277016352;
#10;x=1278016352;
#10;x=1279016352;
#10;x=1280016352;
#10;x=1281016352;
#10;x=1282016352;
#10;x=1283016352;
#10;x=1284016352;
#10;x=1285016352;
#10;x=1286016352;
#10;x=1287016352;
#10;x=1288016352;
#10;x=1289016352;
#10;x=1290016352;
#10;x=1291016352;
#10;x=1292016352;
#10;x=1293016352;
#10;x=1294016352;
#10;x=1295016352;
#10;x=1296016352;
#10;x=1297016352;
#10;x=1298016352;
#10;x=1299016352;
#10;x=1300016352;
#10;x=1301016352;
#10;x=1302016352;
#10;x=1303016352;
#10;x=1304016352;
#10;x=1305016352;
#10;x=1306016352;
#10;x=1307016352;
#10;x=1308016352;
#10;x=1309016352;
#10;x=1310016352;
#10;x=1311016352;
#10;x=1312016352;
#10;x=1313016352;
#10;x=1314016352;
#10;x=1315016352;
#10;x=1316016352;
#10;x=1317016352;
#10;x=1318016352;
#10;x=1319016352;
#10;x=1320016352;
#10;x=1321016352;
#10;x=1322016352;
#10;x=1323016352;
#10;x=1324016352;
#10;x=1325016352;
#10;x=1326016352;
#10;x=1327016352;
#10;x=1328016352;
#10;x=1329016352;
#10;x=1330016352;
#10;x=1331016352;
#10;x=1332016352;
#10;x=1333016352;
#10;x=1334016352;
#10;x=1335016352;
#10;x=1336016352;
#10;x=1337016352;
#10;x=1338016352;
#10;x=1339016352;
#10;x=1340016352;
#10;x=1341016352;
#10;x=1342016352;
#10;x=1343016352;
#10;x=1344016352;
#10;x=1345016352;
#10;x=1346016352;
#10;x=1347016352;
#10;x=1348016352;
#10;x=1349016352;
#10;x=1350016352;
#10;x=1351016352;
#10;x=1352016352;
#10;x=1353016352;
#10;x=1354016352;
#10;x=1355016352;
#10;x=1356016352;
#10;x=1357016352;
#10;x=1358016352;
#10;x=1359016352;
#10;x=1360016352;
#10;x=1361016352;
#10;x=1362016352;
#10;x=1363016352;
#10;x=1364016352;
#10;x=1365016352;
#10;x=1366016352;
#10;x=1367016352;
#10;x=1368016352;
#10;x=1369016352;
#10;x=1370016352;
#10;x=1371016352;
#10;x=1372016352;
#10;x=1373016352;
#10;x=1374016352;
#10;x=1375016352;
#10;x=1376016352;
#10;x=1377016352;
#10;x=1378016352;
#10;x=1379016352;
#10;x=1380016352;
#10;x=1381016352;
#10;x=1382016352;
#10;x=1383016352;
#10;x=1384016352;
#10;x=1385016352;
#10;x=1386016352;
#10;x=1387016352;
#10;x=1388016352;
#10;x=1389016352;
#10;x=1390016352;
#10;x=1391016352;
#10;x=1392016352;
#10;x=1393016352;
#10;x=1394016352;
#10;x=1395016352;
#10;x=1396016352;
#10;x=1397016352;
#10;x=1398016352;
#10;x=1399016352;
#10;x=1400016352;
#10;x=1401016352;
#10;x=1402016352;
#10;x=1403016352;
#10;x=1404016352;
#10;x=1405016352;
#10;x=1406016352;
#10;x=1407016352;
#10;x=1408016352;
#10;x=1409016352;
#10;x=1410016352;
#10;x=1411016352;
#10;x=1412016352;
#10;x=1413016352;
#10;x=1414016352;
#10;x=1415016352;
#10;x=1416016352;
#10;x=1417016352;
#10;x=1418016352;
#10;x=1419016352;
#10;x=1420016352;
#10;x=1421016352;
#10;x=1422016352;
#10;x=1423016352;
#10;x=1424016352;
#10;x=1425016352;
#10;x=1426016352;
#10;x=1427016352;
#10;x=1428016352;
#10;x=1429016352;
#10;x=1430016352;
#10;x=1431016352;
#10;x=1432016352;
#10;x=1433016352;
#10;x=1434016352;
#10;x=1435016352;
#10;x=1436016352;
#10;x=1437016352;
#10;x=1438016352;
#10;x=1439016352;
#10;x=1440016352;
#10;x=1441016352;
#10;x=1442016352;
#10;x=1443016352;
#10;x=1444016352;
#10;x=1445016352;
#10;x=1446016352;
#10;x=1447016352;
#10;x=1448016352;
#10;x=1449016352;
#10;x=1450016352;
#10;x=1451016352;
#10;x=1452016352;
#10;x=1453016352;
#10;x=1454016352;
#10;x=1455016352;
#10;x=1456016352;
#10;x=1457016352;
#10;x=1458016352;
#10;x=1459016352;
#10;x=1460016352;
#10;x=1461016352;
#10;x=1462016352;
#10;x=1463016352;
#10;x=1464016352;
#10;x=1465016352;
#10;x=1466016352;
#10;x=1467016352;
#10;x=1468016352;
#10;x=1469016352;
#10;x=1470016352;
#10;x=1471016352;
#10;x=1472016352;
#10;x=1473016352;
#10;x=1474016352;
#10;x=1475016352;
#10;x=1476016352;
#10;x=1477016352;
#10;x=1478016352;
#10;x=1479016352;
#10;x=1480016352;
#10;x=1481016352;
#10;x=1482016352;
#10;x=1483016352;
#10;x=1484016352;
#10;x=1485016352;
#10;x=1486016352;
#10;x=1487016352;
#10;x=1488016352;
#10;x=1489016352;
#10;x=1490016352;
#10;x=1491016352;
#10;x=1492016352;
#10;x=1493016352;
#10;x=1494016352;
#10;x=1495016352;
#10;x=1496016352;
#10;x=1497016352;
#10;x=1498016352;
#10;x=1499016352;
#10;x=1500016352;
#10;x=1501016352;
#10;x=1502016352;
#10;x=1503016352;
#10;x=1504016352;
#10;x=1505016352;
#10;x=1506016352;
#10;x=1507016352;
#10;x=1508016352;
#10;x=1509016352;
#10;x=1510016352;
#10;x=1511016352;
#10;x=1512016352;
#10;x=1513016352;
#10;x=1514016352;
#10;x=1515016352;
#10;x=1516016352;
#10;x=1517016352;
#10;x=1518016352;
#10;x=1519016352;
#10;x=1520016352;
#10;x=1521016352;
#10;x=1522016352;
#10;x=1523016352;
#10;x=1524016352;
#10;x=1525016352;
#10;x=1526016352;
#10;x=1527016352;
#10;x=1528016352;
#10;x=1529016352;
#10;x=1530016352;
#10;x=1531016352;
#10;x=1532016352;
#10;x=1533016352;
#10;x=1534016352;
#10;x=1535016352;
#10;x=1536016352;
#10;x=1537016352;
#10;x=1538016352;
#10;x=1539016352;
#10;x=1540016352;
#10;x=1541016352;
#10;x=1542016352;
#10;x=1543016352;
#10;x=1544016352;
#10;x=1545016352;
#10;x=1546016352;
#10;x=1547016352;
#10;x=1548016352;
#10;x=1549016352;
#10;x=1550016352;
#10;x=1551016352;
#10;x=1552016352;
#10;x=1553016352;
#10;x=1554016352;
#10;x=1555016352;
#10;x=1556016352;
#10;x=1557016352;
#10;x=1558016352;
#10;x=1559016352;
#10;x=1560016352;
#10;x=1561016352;
#10;x=1562016352;
#10;x=1563016352;
#10;x=1564016352;
#10;x=1565016352;
#10;x=1566016352;
#10;x=1567016352;
#10;x=1568016352;
#10;x=1569016352;
#10;x=1570016352;
#10;x=1571016352;
#10;x=1572016352;
#10;x=1573016352;
#10;x=1574016352;
#10;x=1575016352;
#10;x=1576016352;
#10;x=1577016352;
#10;x=1578016352;
#10;x=1579016352;
#10;x=1580016352;
#10;x=1581016352;
#10;x=1582016352;
#10;x=1583016352;
#10;x=1584016352;
#10;x=1585016352;
#10;x=1586016352;
#10;x=1587016352;
#10;x=1588016352;
#10;x=1589016352;
#10;x=1590016352;
#10;x=1591016352;
#10;x=1592016352;
#10;x=1593016352;
#10;x=1594016352;
#10;x=1595016352;
#10;x=1596016352;
#10;x=1597016352;
#10;x=1598016352;
#10;x=1599016352;
#10;x=1600016352;
#10;x=1601016352;
#10;x=1602016352;
#10;x=1603016352;
#10;x=1604016352;
#10;x=1605016352;
#10;x=1606016352;
#10;x=1607016352;
#10;x=1608016352;
#10;x=1609016352;
#10;x=1610016352;
#10;x=1611016352;
#10;x=1612016352;
#10;x=1613016352;
#10;x=1614016352;
#10;x=1615016352;
#10;x=1616016352;
#10;x=1617016352;
#10;x=1618016352;
#10;x=1619016352;
#10;x=1620016352;
#10;x=1621016352;
#10;x=1622016352;
#10;x=1623016352;
#10;x=1624016352;
#10;x=1625016352;
#10;x=1626016352;
#10;x=1627016352;
#10;x=1628016352;
#10;x=1629016352;
#10;x=1630016352;
#10;x=1631016352;
#10;x=1632016352;
#10;x=1633016352;
#10;x=1634016352;
#10;x=1635016352;
#10;x=1636016352;
#10;x=1637016352;
#10;x=1638016352;
#10;x=1639016352;
#10;x=1640016352;
#10;x=1641016352;
#10;x=1642016352;
#10;x=1643016352;
#10;x=1644016352;
#10;x=1645016352;
#10;x=1646016352;
#10;x=1647016352;
#10;x=1648016352;
#10;x=1649016352;
#10;x=1650016352;
#10;x=1651016352;
#10;x=1652016352;
#10;x=1653016352;
#10;x=1654016352;
#10;x=1655016352;
#10;x=1656016352;
#10;x=1657016352;
#10;x=1658016352;
#10;x=1659016352;
#10;x=1660016352;
#10;x=1661016352;
#10;x=1662016352;
#10;x=1663016352;
#10;x=1664016352;
#10;x=1665016352;
#10;x=1666016352;
#10;x=1667016352;
#10;x=1668016352;
#10;x=1669016352;
#10;x=1670016352;
#10;x=1671016352;
#10;x=1672016352;
#10;x=1673016352;
#10;x=1674016352;
#10;x=1675016352;
#10;x=1676016352;
#10;x=1677016352;
#10;x=1678016352;
#10;x=1679016352;
#10;x=1680016352;
#10;x=1681016352;
#10;x=1682016352;
#10;x=1683016352;
#10;x=1684016352;
#10;x=1685016352;
#10;x=1686016352;
#10;x=1687016352;
#10;x=1688016352;
#10;x=1689016352;
#10;x=1690016352;
#10;x=1691016352;
#10;x=1692016352;
#10;x=1693016352;
#10;x=1694016352;
#10;x=1695016352;
#10;x=1696016352;
#10;x=1697016352;
#10;x=1698016352;
#10;x=1699016352;
#10;x=1700016352;
#10;x=1701016352;
#10;x=1702016352;
#10;x=1703016352;
#10;x=1704016352;
#10;x=1705016352;
#10;x=1706016352;
#10;x=1707016352;
#10;x=1708016352;
#10;x=1709016352;
#10;x=1710016352;
#10;x=1711016352;
#10;x=1712016352;
#10;x=1713016352;
#10;x=1714016352;
#10;x=1715016352;
#10;x=1716016352;
#10;x=1717016352;
#10;x=1718016352;
#10;x=1719016352;
#10;x=1720016352;
#10;x=1721016352;
#10;x=1722016352;
#10;x=1723016352;
#10;x=1724016352;
#10;x=1725016352;
#10;x=1726016352;
#10;x=1727016352;
#10;x=1728016352;
#10;x=1729016352;
#10;x=1730016352;
#10;x=1731016352;
#10;x=1732016352;
#10;x=1733016352;
#10;x=1734016352;
#10;x=1735016352;
#10;x=1736016352;
#10;x=1737016352;
#10;x=1738016352;
#10;x=1739016352;
#10;x=1740016352;
#10;x=1741016352;
#10;x=1742016352;
#10;x=1743016352;
#10;x=1744016352;
#10;x=1745016352;
#10;x=1746016352;
#10;x=1747016352;
#10;x=1748016352;
#10;x=1749016352;
#10;x=1750016352;
#10;x=1751016352;
#10;x=1752016352;
#10;x=1753016352;
#10;x=1754016352;
#10;x=1755016352;
#10;x=1756016352;
#10;x=1757016352;
#10;x=1758016352;
#10;x=1759016352;
#10;x=1760016352;
#10;x=1761016352;
#10;x=1762016352;
#10;x=1763016352;
#10;x=1764016352;
#10;x=1765016352;
#10;x=1766016352;
#10;x=1767016352;
#10;x=1768016352;
#10;x=1769016352;
#10;x=1770016352;
#10;x=1771016352;
#10;x=1772016352;
#10;x=1773016352;
#10;x=1774016352;
#10;x=1775016352;
#10;x=1776016352;
#10;x=1777016352;
#10;x=1778016352;
#10;x=1779016352;
#10;x=1780016352;
#10;x=1781016352;
#10;x=1782016352;
#10;x=1783016352;
#10;x=1784016352;
#10;x=1785016352;
#10;x=1786016352;
#10;x=1787016352;
#10;x=1788016352;
#10;x=1789016352;
#10;x=1790016352;
#10;x=1791016352;
#10;x=1792016352;
#10;x=1793016352;
#10;x=1794016352;
#10;x=1795016352;
#10;x=1796016352;
#10;x=1797016352;
#10;x=1798016352;
#10;x=1799016352;
#10;x=1800016352;
#10;x=1801016352;
#10;x=1802016352;
#10;x=1803016352;
#10;x=1804016352;
#10;x=1805016352;
#10;x=1806016352;
#10;x=1807016352;
#10;x=1808016352;
#10;x=1809016352;
#10;x=1810016352;
#10;x=1811016352;
#10;x=1812016352;
#10;x=1813016352;
#10;x=1814016352;
#10;x=1815016352;
#10;x=1816016352;
#10;x=1817016352;
#10;x=1818016352;
#10;x=1819016352;
#10;x=1820016352;
#10;x=1821016352;
#10;x=1822016352;
#10;x=1823016352;
#10;x=1824016352;
#10;x=1825016352;
#10;x=1826016352;
#10;x=1827016352;
#10;x=1828016352;
#10;x=1829016352;
#10;x=1830016352;
#10;x=1831016352;
#10;x=1832016352;
#10;x=1833016352;
#10;x=1834016352;
#10;x=1835016352;
#10;x=1836016352;
#10;x=1837016352;
#10;x=1838016352;
#10;x=1839016352;
#10;x=1840016352;
#10;x=1841016352;
#10;x=1842016352;
#10;x=1843016352;
#10;x=1844016352;
#10;x=1845016352;
#10;x=1846016352;
#10;x=1847016352;
#10;x=1848016352;
#10;x=1849016352;
#10;x=1850016352;
#10;x=1851016352;
#10;x=1852016352;
#10;x=1853016352;
#10;x=1854016352;
#10;x=1855016352;
#10;x=1856016352;
#10;x=1857016352;
#10;x=1858016352;
#10;x=1859016352;
#10;x=1860016352;
#10;x=1861016352;
#10;x=1862016352;
#10;x=1863016352;
#10;x=1864016352;
#10;x=1865016352;
#10;x=1866016352;
#10;x=1867016352;
#10;x=1868016352;
#10;x=1869016352;
#10;x=1870016352;
#10;x=1871016352;
#10;x=1872016352;
#10;x=1873016352;
#10;x=1874016352;
#10;x=1875016352;
#10;x=1876016352;
#10;x=1877016352;
#10;x=1878016352;
#10;x=1879016352;
#10;x=1880016352;
#10;x=1881016352;
#10;x=1882016352;
#10;x=1883016352;
#10;x=1884016352;
#10;x=1885016352;
#10;x=1886016352;
#10;x=1887016352;
#10;x=1888016352;
#10;x=1889016352;
#10;x=1890016352;
#10;x=1891016352;
#10;x=1892016352;
#10;x=1893016352;
#10;x=1894016352;
#10;x=1895016352;
#10;x=1896016352;
#10;x=1897016352;
#10;x=1898016352;
#10;x=1899016352;
#10;x=1900016352;
#10;x=1901016352;
#10;x=1902016352;
#10;x=1903016352;
#10;x=1904016352;
#10;x=1905016352;
#10;x=1906016352;
#10;x=1907016352;
#10;x=1908016352;
#10;x=1909016352;
#10;x=1910016352;
#10;x=1911016352;
#10;x=1912016352;
#10;x=1913016352;
#10;x=1914016352;
#10;x=1915016352;
#10;x=1916016352;
#10;x=1917016352;
#10;x=1918016352;
#10;x=1919016352;
#10;x=1920016352;
#10;x=1921016352;
#10;x=1922016352;
#10;x=1923016352;
#10;x=1924016352;
#10;x=1925016352;
#10;x=1926016352;
#10;x=1927016352;
#10;x=1928016352;
#10;x=1929016352;
#10;x=1930016352;
#10;x=1931016352;
#10;x=1932016352;
#10;x=1933016352;
#10;x=1934016352;
#10;x=1935016352;
#10;x=1936016352;
#10;x=1937016352;
#10;x=1938016352;
#10;x=1939016352;
#10;x=1940016352;
#10;x=1941016352;
#10;x=1942016352;
#10;x=1943016352;
#10;x=1944016352;
#10;x=1945016352;
#10;x=1946016352;
#10;x=1947016352;
#10;x=1948016352;
#10;x=1949016352;
#10;x=1950016352;
#10;x=1951016352;
#10;x=1952016352;
#10;x=1953016352;
#10;x=1954016352;
#10;x=1955016352;
#10;x=1956016352;
#10;x=1957016352;
#10;x=1958016352;
#10;x=1959016352;
#10;x=1960016352;
#10;x=1961016352;
#10;x=1962016352;
#10;x=1963016352;
#10;x=1964016352;
#10;x=1965016352;
#10;x=1966016352;
#10;x=1967016352;
#10;x=1968016352;
#10;x=1969016352;
#10;x=1970016352;
#10;x=1971016352;
#10;x=1972016352;
#10;x=1973016352;
#10;x=1974016352;
#10;x=1975016352;
#10;x=1976016352;
#10;x=1977016352;
#10;x=1978016352;
#10;x=1979016352;
#10;x=1980016352;
#10;x=1981016352;
#10;x=1982016352;
#10;x=1983016352;
#10;x=1984016352;
#10;x=1985016352;
#10;x=1986016352;
#10;x=1987016352;
#10;x=1988016352;
#10;x=1989016352;
#10;x=1990016352;
#10;x=1991016352;
#10;x=1992016352;
#10;x=1993016352;
#10;x=1994016352;
#10;x=1995016352;
#10;x=1996016352;
#10;x=1997016352;
#10;x=1998016352;
#10;x=1999016352;
#10;x=2000016352;
#10;x=2001016352;
#10;x=2002016352;
#10;x=2003016352;
#10;x=2004016352;
#10;x=2005016352;
#10;x=2006016352;
#10;x=2007016352;
#10;x=2008016352;
#10;x=2009016352;
#10;x=2010016352;
#10;x=2011016352;
#10;x=2012016352;
#10;x=2013016352;
#10;x=2014016352;
#10;x=2015016352;
#10;x=2016016352;
#10;x=2017016352;
#10;x=2018016352;
#10;x=2019016352;
#10;x=2020016352;
#10;x=2021016352;
#10;x=2022016352;
#10;x=2023016352;
#10;x=2024016352;
#10;x=2025016352;
#10;x=2026016352;
#10;x=2027016352;
#10;x=2028016352;
#10;x=2029016352;
#10;x=2030016352;
#10;x=2031016352;
#10;x=2032016352;
#10;x=2033016352;
#10;x=2034016352;
#10;x=2035016352;
#10;x=2036016352;
#10;x=2037016352;
#10;x=2038016352;
#10;x=2039016352;
#10;x=2040016352;
#10;x=2041016352;
#10;x=2042016352;
#10;x=2043016352;
#10;x=2044016352;
#10;x=2045016352;
#10;x=2046016352;
#10;x=2047016352;
#10;x=2048016352;
#10;x=2049016352;
#10;x=2050016352;
#10;x=2051016352;
#10;x=2052016352;
#10;x=2053016352;
#10;x=2054016352;
#10;x=2055016352;
#10;x=2056016352;
#10;x=2057016352;
#10;x=2058016352;
#10;x=2059016352;
#10;x=2060016352;
#10;x=2061016352;
#10;x=2062016352;
#10;x=2063016352;
#10;x=2064016352;
#10;x=2065016352;
#10;x=2066016352;
#10;x=2067016352;
#10;x=2068016352;
#10;x=2069016352;
#10;x=2070016352;
#10;x=2071016352;
#10;x=2072016352;
#10;x=2073016352;
#10;x=2074016352;
#10;x=2075016352;
#10;x=2076016352;
#10;x=2077016352;
#10;x=2078016352;
#10;x=2079016352;
#10;x=2080016352;
#10;x=2081016352;
#10;x=2082016352;
#10;x=2083016352;
#10;x=2084016352;
#10;x=2085016352;
#10;x=2086016352;
#10;x=2087016352;
#10;x=2088016352;
#10;x=2089016352;
#10;x=2090016352;
#10;x=2091016352;
#10;x=2092016352;
#10;x=2093016352;
#10;x=2094016352;
#10;x=2095016352;
#10;x=2096016352;
#10;x=2097016352;
#10;x=2098016352;
#10;x=2099016352;
#10;x=2100016352;
#10;x=2101016352;
#10;x=2102016352;
#10;x=2103016352;
#10;x=2104016352;
#10;x=2105016352;
#10;x=2106016352;
#10;x=2107016352;
#10;x=2108016352;
#10;x=2109016352;
#10;x=2110016352;
#10;x=2111016352;
#10;x=2112016352;
#10;x=2113016352;
#10;x=2114016352;
#10;x=2115016352;
#10;x=2116016352;
#10;x=2117016352;
#10;x=2118016352;
#10;x=2119016352;
#10;x=2120016352;
#10;x=2121016352;
#10;x=2122016352;
#10;x=2123016352;
#10;x=2124016352;
#10;x=2125016352;
#10;x=2126016352;
#10;x=2127016352;
#10;x=2128016352;
#10;x=2129016352;
#10;x=2130016352;
#10;x=2131016352;
#10;x=2132016352;
#10;x=2133016352;
#10;x=2134016352;
#10;x=2135016352;
#10;x=2136016352;
#10;x=2137016352;
#10;x=2138016352;
#10;x=2139016352;
#10;x=2140016352;
#10;x=2141016352;
#10;x=2142016352;
#10;x=2143016352;
#10;x=2144016352;
#10;x=2145016352;
#10;x=2146016352;
#10;x=2147016352;

        #10;
        $finish;
    end
    
    // Monitor
    always @(posedge clk) begin
        $display("%d, %d", x, y);
    end
    
endmodule
