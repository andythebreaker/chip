`include "systolic_array.v"
module connect_main_mem_with_pe_array(
  //input mem addr 
)