`include "memory32x20.sv"

module Memory32x20_TB;
  // Parameters
  `define addr_width 20
  `define addr_height 1048576
  `define mem_width 32
  `define M1(x) (x-1)

  // Inputs
  logic clk;
  logic rst;
  logic [`M1(`addr_width):0] addr;
  logic we;
  logic [`M1(`mem_width):0] data_in;
  
  // Outputs
  logic [`M1(`mem_width):0] data_out;
  
  // Instantiate the module under test
  Memory32x20 dut (
    .clk(clk),
    .rst(rst),
    .addr(addr),
    .we(we),
    .data_in(data_in),
    .data_out(data_out)
  );
  
  // Clock generator
  always #5 clk = ~clk;

  initial begin
    $fsdbDumpfile("Memory32x20_TB.fsdb");
    $fsdbDumpvars("+all");
  end
  
  initial begin
    // Initialize inputs
    clk = 0;
    rst = 1;
    addr = 0;
    we = 0;
    data_in = 0;
    
    // Reset the module
    #10 rst = 0;
    
    // Write data to memory

#10 addr = 20'd0; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd19; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd20; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd21; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd22; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd23; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd24; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd25; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd26; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd27; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd28; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd29; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd30; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd31; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd32; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd33; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd34; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd35; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd36; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd37; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd38; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd39; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd40; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd41; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd42; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd43; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd44; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd45; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd46; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd47; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd48; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd49; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd50; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd51; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd52; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd53; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd54; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd55; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd56; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd57; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd58; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd59; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd60; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd61; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd62; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd63; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd64; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd65; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd66; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd67; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd68; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd69; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd70; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd71; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd72; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd73; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd74; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd75; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd76; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd77; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd78; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd79; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd80; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd81; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd82; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd83; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd84; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd85; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd86; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd87; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd88; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd89; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd90; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd91; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd92; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd93; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd94; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd95; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd96; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd97; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd98; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd99; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd100; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd102; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd103; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd104; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd105; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd106; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd107; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd108; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd109; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd110; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd111; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd112; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd113; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd114; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd115; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd116; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd117; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd118; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd119; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd120; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd121; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd122; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd123; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd124; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd125; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd126; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd127; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd128; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd129; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd130; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd131; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd132; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd133; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd135; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd137; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd138; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd139; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd140; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd141; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd142; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd143; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd144; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd145; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd146; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd147; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd148; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd149; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd150; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd151; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd152; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd153; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd154; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd155; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd156; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd157; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd158; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd159; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd160; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd161; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd162; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd163; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd164; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd165; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd166; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd167; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd168; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd169; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd170; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd171; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd172; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd173; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd174; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd175; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd176; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd177; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd178; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd179; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd180; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd181; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd182; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd183; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd184; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd185; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd186; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd187; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd188; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd189; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd190; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd191; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd192; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd193; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd194; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd195; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd196; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd197; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd198; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd199; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd200; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd201; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd202; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd203; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd204; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd205; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd206; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd207; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd208; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd209; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd210; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd211; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd212; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd213; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd214; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd215; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd216; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd217; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd218; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd219; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd220; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd221; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd222; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd223; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd224; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd225; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd226; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd227; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd228; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd229; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd230; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd231; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd232; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd233; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd234; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd235; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd236; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd237; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd238; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd239; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd240; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd241; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd242; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd243; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd244; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd245; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd246; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd247; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd249; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd250; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd251; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd252; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd253; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd254; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd255; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd256; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd257; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd258; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd259; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd260; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd261; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd262; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd263; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd264; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd265; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd266; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd267; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd268; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd269; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd271; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd272; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd273; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd274; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd275; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd277; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd278; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd279; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd280; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd281; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd282; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd283; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd284; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd285; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd286; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd287; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd288; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd289; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd290; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd291; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd292; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd293; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd294; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd295; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd296; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd298; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd299; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd300; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd301; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd302; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd303; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd304; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd305; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd306; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd307; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd308; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd309; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd310; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd311; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd312; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd313; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd314; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd315; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd316; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd318; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd319; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd320; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd321; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd322; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd323; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd324; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd325; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd328; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd329; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd330; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd331; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd333; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd334; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd335; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd337; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd338; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd339; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd340; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd341; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd342; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd343; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd344; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd346; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd347; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd348; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd349; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd350; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd351; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd352; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd353; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd354; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd355; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd356; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd357; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd358; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd359; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd360; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd361; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd362; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd363; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd364; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd365; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd366; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd367; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd368; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd369; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd370; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd371; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd372; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd374; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd375; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd376; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd377; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd378; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd379; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd383; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd384; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd385; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd386; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd387; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd389; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd390; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd391; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd392; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd393; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd394; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd395; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd396; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd397; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd398; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd399; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd400; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd402; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd403; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd404; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd405; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd406; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd407; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd411; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd412; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd413; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd414; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd415; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd416; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd417; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd418; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd419; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd420; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd421; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd422; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd423; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd424; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd425; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd426; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd427; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd428; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd430; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd431; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd432; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd433; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd434; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd435; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd436; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd438; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd439; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd440; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd441; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd442; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd443; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd444; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd445; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd446; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd447; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd448; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd449; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd450; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd451; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd452; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd453; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd454; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd455; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd456; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd457; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd459; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd460; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd461; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd462; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd463; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd464; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd465; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd466; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd467; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd468; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd469; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd470; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd471; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd472; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd473; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd474; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd475; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd476; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd477; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd478; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd479; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd480; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd481; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd482; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd484; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd485; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd486; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd487; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd488; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd489; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd490; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd491; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd492; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd493; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd494; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd495; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd496; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd497; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd498; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd499; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd500; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd501; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd502; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd503; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd504; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd505; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd506; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd507; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd508; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd509; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd510; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd511; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd512; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd514; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd515; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd516; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd517; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd518; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd519; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd520; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd521; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd522; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd523; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd524; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd525; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd526; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd527; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd528; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd529; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd530; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd531; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd532; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd533; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd534; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd535; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd536; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd537; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd538; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd539; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd540; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd542; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd543; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd544; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd545; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd546; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd547; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd548; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd549; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd550; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd551; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd552; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd553; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd554; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd555; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd556; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd557; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd558; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd559; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd560; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd561; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd562; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd563; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd564; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd565; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd566; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd567; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd568; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd569; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd570; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd571; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd572; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd573; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd574; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd575; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd576; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd577; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd578; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd579; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd580; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd581; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd582; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd583; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd584; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd585; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd586; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd587; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd588; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd589; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd590; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd591; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd592; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd593; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd594; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd595; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd596; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd597; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd598; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd599; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd600; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd601; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd602; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd603; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd604; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd605; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd606; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd607; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd608; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd609; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd610; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd611; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd612; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd613; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd614; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd615; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd616; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd617; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd618; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd619; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd620; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd621; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd622; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd623; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd624; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd625; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd626; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd627; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd628; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd629; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd630; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd631; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd632; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd633; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd634; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd635; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd636; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd637; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd638; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd639; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd640; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd641; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd642; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd643; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd644; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd645; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd646; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd647; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd648; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd649; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd650; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd651; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd652; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd653; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd654; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd655; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd656; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd657; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd658; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd659; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd660; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd661; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd663; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd664; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd665; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd666; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd667; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd668; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd669; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd670; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd671; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd672; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd673; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd674; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd675; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd676; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd677; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd678; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd679; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd680; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd681; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd682; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd683; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd684; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd685; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd686; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd687; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd688; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd689; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd690; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd691; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd692; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd693; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd694; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd695; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd696; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd697; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd698; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd699; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd700; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd701; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd702; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd703; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd704; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd705; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd706; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd707; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd708; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd709; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd710; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd712; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd713; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd714; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd715; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd716; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd717; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd718; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd719; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd720; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd721; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd722; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd723; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd724; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd725; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd726; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd727; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd728; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd729; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd730; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd731; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd732; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd733; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd734; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd735; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd736; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd737; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd738; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd739; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd740; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd741; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd742; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd743; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd744; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd746; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd747; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd748; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd749; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd750; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd751; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd752; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd753; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd754; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd755; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd756; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd757; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd758; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd759; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd760; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd761; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd762; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd763; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd764; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd765; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd767; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd768; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd769; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd770; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd771; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd773; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd774; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd775; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd776; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd777; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd778; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd779; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd780; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd781; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd782; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd783; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd784; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd785; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd786; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd787; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd788; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd789; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd790; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd791; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd792; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd793; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd795; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd796; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd797; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd798; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd799; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd800; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd801; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd802; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd803; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd804; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd805; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd806; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd807; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd808; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd809; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd810; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd811; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd812; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd813; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd814; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd815; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd816; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd817; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd818; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd819; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd820; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd821; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd822; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd823; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd824; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd825; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd826; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd827; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd828; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd829; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd830; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd831; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd832; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd833; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd834; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd835; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd836; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd837; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd838; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd839; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd840; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd841; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd842; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd843; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd844; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd845; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd846; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd847; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd848; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd849; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd850; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd851; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd852; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd853; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd854; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd855; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd856; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd857; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd858; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd859; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd860; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd861; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd862; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd863; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd864; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd865; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd866; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd867; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd868; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd869; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd870; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd871; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd872; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd873; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd874; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd875; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd876; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd877; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd878; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd879; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd880; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd881; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd882; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd883; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd884; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd885; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd887; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd888; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd889; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd890; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd891; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd892; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd893; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd894; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd895; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd896; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd897; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd898; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd899; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd900; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd901; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd902; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd903; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd904; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd905; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd906; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd907; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd908; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd909; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd910; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd911; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd912; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd914; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd915; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd916; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd917; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd918; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd919; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd920; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd921; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd922; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd923; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd924; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd925; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd926; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd927; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd928; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd929; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd930; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd931; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd932; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd933; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd934; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd935; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd936; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd937; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd938; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd939; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd940; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd941; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd942; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd943; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd944; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd945; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd946; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd947; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd948; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd949; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd950; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd951; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd952; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd953; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd954; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd955; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd956; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd957; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd958; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd959; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd960; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd961; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd962; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd963; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd964; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd965; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd966; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd967; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd968; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd969; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd970; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd971; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd972; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd973; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd974; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd975; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd976; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd977; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd978; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd979; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd980; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd981; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd982; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd983; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd984; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd985; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd986; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd987; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd988; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd989; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd990; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd991; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd993; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd994; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd995; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd996; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd997; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd998; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd999; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1000; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1001; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1002; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1003; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1004; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1005; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1006; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1007; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1008; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1009; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1010; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1011; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1012; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1013; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1014; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1015; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1016; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1017; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1018; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1020; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1021; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1022; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1023; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1024; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1025; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1026; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1027; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1028; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1029; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1030; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1031; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd1032; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1033; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1034; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1035; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1036; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1037; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1038; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1039; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1040; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1041; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1042; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1043; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1044; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1045; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1046; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1047; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1048; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1049; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1050; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1051; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1052; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1053; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1054; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1055; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1056; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1057; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1058; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1059; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1060; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1062; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1063; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1064; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1065; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1066; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1067; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1068; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1069; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1070; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1071; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1072; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1073; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1074; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1075; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1076; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1077; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1078; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1079; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1080; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1081; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1082; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1083; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1084; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1085; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1086; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1087; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1088; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1089; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1090; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1091; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1092; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1093; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1094; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1095; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1096; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1097; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1098; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1099; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1100; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1102; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1103; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1104; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1105; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1106; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1107; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1108; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1109; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1110; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1111; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1112; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1113; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1114; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1115; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1116; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1117; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1118; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1119; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1120; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1121; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1122; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1123; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1124; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1125; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1126; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1127; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1128; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1129; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1130; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1131; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1132; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1133; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd1134; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1135; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1136; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd1137; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1138; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1139; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1140; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1141; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1142; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1143; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1144; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1145; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1146; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1147; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1148; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1149; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1150; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1151; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1152; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1153; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1154; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1155; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1156; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1157; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1158; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1159; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1160; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1161; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1162; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd1163; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1164; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd6;
#10 addr = 20'd1165; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1166; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1167; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1168; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1169; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1170; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1171; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1172; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1173; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1174; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1175; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1176; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1177; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1178; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1179; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1180; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1181; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1182; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1183; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1184; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1185; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1186; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1187; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1189; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1190; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1191; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1192; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd1193; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1194; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1195; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1196; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1197; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1198; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1199; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1200; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1201; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1202; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1203; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1204; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1205; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1206; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1207; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1208; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1209; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1210; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1211; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1212; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1213; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1214; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1215; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1216; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd1217; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1218; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1219; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1220; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd1221; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1222; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1223; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1224; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1225; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1226; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1227; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1228; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1229; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1230; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1231; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1232; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1233; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1234; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1235; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1236; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1237; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1238; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1239; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1240; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1241; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1242; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1243; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1244; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1245; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1246; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1247; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd1248; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1249; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1250; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1251; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1252; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1253; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1254; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1255; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1256; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1257; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1258; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1259; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1260; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1261; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1262; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1263; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1264; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1265; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1266; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1267; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1268; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1269; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1271; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1272; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1273; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1274; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1275; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1276; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd1277; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1278; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1279; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1280; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1281; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1282; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1283; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1284; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1285; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1286; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1287; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1288; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1289; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1290; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1291; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1292; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1293; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1294; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1295; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1296; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1298; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1299; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1300; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1301; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1302; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1303; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1304; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1305; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1306; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1307; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1308; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1309; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1310; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1311; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1312; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1313; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1314; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1315; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1316; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1317; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1318; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1319; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1320; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1321; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1322; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1323; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd1324; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1325; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1328; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1329; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1330; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1331; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1332; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1333; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1334; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1335; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1336; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1337; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1338; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd1339; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1340; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1341; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1342; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1343; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1344; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1345; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1346; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1347; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1348; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1349; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1350; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1351; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1352; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1353; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1354; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1355; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1356; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1357; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1358; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1359; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1360; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1361; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1362; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1363; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1364; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1365; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1366; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1367; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1368; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1369; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1370; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1371; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1372; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1373; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1374; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1375; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1376; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1377; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1378; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1379; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1383; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd1384; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1385; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1386; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1387; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd1388; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1389; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd1390; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1391; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1392; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1393; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1394; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1395; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1396; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1397; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1398; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1399; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1401; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1402; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1403; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1404; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1405; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1406; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1407; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1410; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1411; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1412; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1413; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1414; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1415; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1416; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1417; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd3;
#10 addr = 20'd1418; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1419; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1420; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1421; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd1422; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1423; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1424; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1425; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1426; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1427; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1428; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1429; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1430; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1431; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1432; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1433; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1434; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd1435; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1436; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1438; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1440; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1441; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1442; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1443; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1444; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1445; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd5;
#10 addr = 20'd1446; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1447; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1448; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1449; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1450; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd1451; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1452; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1453; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd1454; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1455; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1456; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1457; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1458; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1459; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1460; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1461; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1462; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd1463; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1464; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1465; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1466; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1467; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1468; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1469; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1470; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1471; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1472; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1473; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd9;
#10 addr = 20'd1474; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1475; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1476; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1477; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1478; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd3;
#10 addr = 20'd1479; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1480; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1481; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd1482; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1483; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1484; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1485; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1486; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1487; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1488; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1489; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1490; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd1491; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1492; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1493; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1495; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1496; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1497; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1498; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1499; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1500; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1501; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd1502; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1503; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1504; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd10;
#10 addr = 20'd1505; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd1506; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd3;
#10 addr = 20'd1507; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1508; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1509; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1510; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1511; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1512; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1513; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1514; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1515; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1516; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1517; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1518; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd1519; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1520; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1521; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1523; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1524; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1525; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1526; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1527; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1528; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1529; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd1530; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1531; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1532; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd1533; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1534; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd4;
#10 addr = 20'd1535; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1536; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1537; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1538; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1539; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1540; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1541; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1542; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1543; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1544; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1545; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1546; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1547; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1548; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1549; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1550; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd1551; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd1552; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1553; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1554; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1555; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1556; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1557; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1558; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1559; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1560; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd1561; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1562; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd5;
#10 addr = 20'd1563; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1564; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1565; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1566; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1567; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1568; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1569; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1570; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1571; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1572; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1573; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1574; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1575; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1576; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1577; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1578; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd1579; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1580; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1581; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1582; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1583; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1584; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1585; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1586; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1588; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1589; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1590; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd5;
#10 addr = 20'd1591; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1592; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1593; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1594; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1595; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1596; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1597; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1598; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1599; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1600; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1601; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1602; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1603; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1604; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1605; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd1607; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1608; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1609; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1610; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1611; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1612; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1613; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd1614; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1615; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1616; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1617; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1618; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd1619; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1620; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1621; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1622; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1623; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1624; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1625; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1626; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1627; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1628; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1629; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1630; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd1631; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1632; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1633; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1636; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1637; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1638; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1639; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1640; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1641; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1642; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1643; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd1644; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd1645; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1646; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd1647; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1648; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1649; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1650; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1651; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1652; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1653; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1654; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1655; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1656; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1657; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1658; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd1659; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1660; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1661; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1663; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1664; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1665; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1666; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1667; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1668; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1669; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1670; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1671; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd1672; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd1673; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1674; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd1675; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1676; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1677; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1678; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1679; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1680; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1682; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1683; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1684; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1685; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1686; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd1687; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1688; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1689; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1690; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1691; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1692; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1693; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1694; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1695; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1696; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1697; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1698; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1699; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd1700; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1701; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1702; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd1703; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1704; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1705; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1706; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1707; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1708; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1709; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1710; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1711; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1712; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1713; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1714; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd1715; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1716; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1717; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1718; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1719; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1720; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1721; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1722; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1723; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1724; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1725; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1726; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1727; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1728; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1729; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1730; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd1731; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1732; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1733; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1734; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1735; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1736; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1737; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1738; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1739; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1740; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1741; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1742; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd1743; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1744; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd1746; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1747; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1748; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1749; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1750; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1751; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1752; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1753; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1754; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd1755; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1756; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1757; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1758; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd1759; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1760; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1761; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1762; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1763; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1764; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1765; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1767; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1768; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1769; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1770; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1771; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1773; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1774; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1775; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1776; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1777; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1778; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1779; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1780; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1781; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1782; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd1783; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1784; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1785; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1786; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1787; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1788; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd1789; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1790; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1791; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1792; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1793; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1795; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1796; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1797; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1798; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd1799; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1800; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1801; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1802; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1803; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1804; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1805; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1806; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1807; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1808; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1809; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1810; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1811; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1812; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1813; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1814; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1815; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd1816; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1817; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1818; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1819; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1820; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1822; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1823; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1824; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1825; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1826; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd1827; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1828; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1829; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1830; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1831; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1832; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1833; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1834; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1835; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1836; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1837; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1838; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1839; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1840; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1841; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd1842; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1843; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1844; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1845; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1846; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1847; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1848; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1849; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1850; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1851; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1852; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1853; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1854; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1855; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd1856; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1857; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1858; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1859; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1860; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1861; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1862; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1863; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1864; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1865; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1866; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1867; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1868; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1869; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1870; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1871; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1872; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1873; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1874; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1875; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1876; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1877; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1878; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1879; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1880; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1881; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1882; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1883; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1884; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd1885; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1886; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1887; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1888; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1889; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1890; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1891; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1892; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1893; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1894; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1895; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1896; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1897; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd1898; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd1899; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1900; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1901; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1902; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1903; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1904; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1905; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1906; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1907; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1908; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1909; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1910; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1911; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd1912; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd1913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1914; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1915; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1917; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1918; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1919; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd1920; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1921; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd1922; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1923; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1924; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1925; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1926; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1927; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1928; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1929; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1930; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1931; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1932; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1933; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1934; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1935; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1936; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1937; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1938; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1939; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1940; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1941; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1942; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1943; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1944; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1945; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd1946; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1947; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1948; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1949; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd1950; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1951; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1952; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1953; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd1954; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1955; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1956; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1957; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd1958; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1959; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1960; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1961; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1962; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1963; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1964; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1965; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1966; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1967; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd1968; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd1969; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd1970; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1971; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1972; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd1973; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd1974; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1975; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd1976; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1977; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd1978; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1979; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1980; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd1981; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1982; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1983; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd1984; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1985; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd1986; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1987; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd1988; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1989; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd1990; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd1991; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1992; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1993; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd1994; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd1995; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd1996; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1997; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd1998; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd1999; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2000; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2001; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2002; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2003; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2004; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2005; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2006; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2007; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2008; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2009; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2010; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2011; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2012; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2013; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2014; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2015; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2016; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2017; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2018; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2020; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2021; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2022; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2023; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2024; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2025; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2026; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2027; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2028; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2029; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2030; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2031; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2032; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2033; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2034; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2035; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2036; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2037; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2038; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2039; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2040; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2041; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2042; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2043; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2044; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2045; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2046; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2047; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2048; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2049; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2050; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2051; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2052; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2053; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2054; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2055; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2056; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2057; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2058; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2059; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2060; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2061; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2062; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2063; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2064; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd2065; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2066; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2067; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2068; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2069; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2070; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2071; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2072; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2073; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2074; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2075; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2076; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2077; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2078; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2079; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2080; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2081; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2082; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2083; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2084; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2085; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd2086; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2087; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2088; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd2089; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2090; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2091; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2092; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd2093; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2094; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2095; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2096; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2097; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2098; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2099; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2100; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2102; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2103; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2104; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2105; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2106; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2107; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2108; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2109; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2110; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2111; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd2112; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2113; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2114; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2115; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2116; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2117; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2118; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2119; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2120; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd2121; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd2122; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2123; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2124; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2125; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2126; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2127; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2128; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2129; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2130; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2131; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2132; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2133; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2134; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2135; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2137; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2138; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2139; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2140; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2141; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2142; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2143; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd2144; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd2145; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2146; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2147; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2148; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2149; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd2150; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2151; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2152; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2153; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2154; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2155; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2156; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2158; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2159; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2160; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2161; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2162; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2163; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2164; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2165; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2166; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2167; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2168; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2169; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd2170; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2171; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd2172; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2173; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2174; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2175; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2176; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd2177; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2178; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2179; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2180; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2181; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2182; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2183; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2184; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2186; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2187; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2188; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2189; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2190; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2191; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2192; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2193; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2194; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2195; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2196; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2197; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2198; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2199; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd2200; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd2201; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2202; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2203; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2204; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2205; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2206; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2207; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2208; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2209; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2210; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2211; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2212; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2213; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2214; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2215; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2216; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2217; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2218; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2219; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2220; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2221; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2222; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2223; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2224; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2225; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2226; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd2227; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd2228; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2229; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2230; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2231; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2232; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2233; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd7;
#10 addr = 20'd2234; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2235; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2236; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2237; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2238; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2239; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2240; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2241; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2242; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2243; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2244; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2245; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2246; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd2247; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2249; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2250; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2251; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2252; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2253; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2254; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2255; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd2256; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2257; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2258; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2259; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2260; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2261; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd2262; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2263; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2264; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2265; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2266; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2267; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2268; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2269; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2270; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2271; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2272; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2273; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2274; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2275; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2276; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2277; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2278; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2279; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2280; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2281; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2282; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd2283; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2284; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2285; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2286; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2287; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2288; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2289; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd2290; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2291; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd2292; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2293; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2294; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2295; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2296; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2298; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2299; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2300; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2301; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2302; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2303; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2304; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2305; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2306; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2307; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2308; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2309; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2310; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd2;
#10 addr = 20'd2311; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd2312; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2313; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2314; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2315; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2316; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2317; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2318; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2319; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2320; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2321; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2322; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2323; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2324; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2325; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2326; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2327; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2328; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2329; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2330; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2331; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2332; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2333; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2334; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2335; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2337; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2338; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd2339; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2340; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2341; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2342; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd2343; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2344; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2345; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2346; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2347; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2348; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2349; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2350; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2351; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2352; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2353; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2354; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2355; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2356; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2357; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2358; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd2359; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2360; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2361; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2362; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2363; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2364; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2365; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2366; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd2367; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2368; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2369; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2370; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd2371; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2372; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2373; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2374; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2375; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2376; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2377; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2378; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2379; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2381; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2383; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2384; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2385; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2386; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd2387; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2389; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2390; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2391; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2392; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2393; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd2394; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd2395; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2396; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2397; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2398; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2399; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2400; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2401; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2402; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2403; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2404; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2405; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2406; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2407; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2409; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2411; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2412; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2413; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2414; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2415; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2416; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2417; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2418; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2419; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2420; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd2421; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd2422; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd2423; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2424; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2425; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2426; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2427; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2428; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2429; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2430; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2431; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2432; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2433; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2434; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2435; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2436; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2437; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2438; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2440; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2441; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2442; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd2443; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2444; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2445; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2446; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2447; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2448; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2449; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2450; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd2451; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2452; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2453; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2454; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd2455; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2456; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd2457; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2458; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2459; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2460; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2461; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2462; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2463; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2464; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2465; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2466; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2468; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2469; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2470; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd2471; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2472; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2473; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2474; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2475; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2476; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2477; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd2478; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2479; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2480; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2481; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2482; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2484; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2485; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2486; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2487; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2488; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2489; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2490; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2491; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2492; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2493; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2494; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2495; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2496; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2497; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2498; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2499; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2500; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2501; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2502; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2503; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2504; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd2505; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd2506; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd2507; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2508; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2509; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2510; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2511; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2512; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2513; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2514; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2515; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2516; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2517; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2518; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2519; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2520; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2521; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2522; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2524; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2525; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2526; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2527; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2528; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2529; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2530; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2531; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2532; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2533; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2534; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd2535; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2536; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2537; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2538; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2539; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2540; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2541; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2542; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2543; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2544; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2545; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2546; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2547; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2548; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2549; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2550; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2551; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2552; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2553; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2554; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2555; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2556; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2557; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2558; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2559; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2560; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2561; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd2562; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2563; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2564; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2565; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2566; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2567; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2568; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2569; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2570; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2571; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2572; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2573; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2574; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2575; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2576; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2577; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2578; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2579; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2580; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2581; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2582; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2583; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2584; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2585; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2586; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2588; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2589; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2590; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2591; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2592; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2593; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2594; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2595; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2596; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2597; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2598; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2599; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2600; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2601; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2602; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2603; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2604; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2605; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2606; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2607; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2608; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2609; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2610; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2611; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2612; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2613; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2614; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2615; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2616; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2617; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2618; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2619; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2620; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2621; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2622; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2623; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2624; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2625; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2626; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2627; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2629; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2630; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2631; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2632; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2633; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2634; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2635; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2636; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2637; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2638; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2639; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2640; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2641; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2642; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2643; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2644; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2645; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2646; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2647; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2648; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2649; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2650; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2651; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2652; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2653; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2654; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd2655; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2656; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2657; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2658; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2659; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2660; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2661; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2662; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2663; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2664; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2665; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2666; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2667; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2668; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2669; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2670; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2671; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2672; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2673; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd2674; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2675; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2676; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2677; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2678; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2679; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2680; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2681; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2682; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd2683; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2684; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2685; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2686; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2687; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2688; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2689; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2690; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2691; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2692; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2693; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2694; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2695; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2696; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2697; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2698; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2699; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2700; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd2701; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd2702; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2703; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2704; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2705; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2706; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2707; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2708; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2709; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2710; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2711; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2712; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2713; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2714; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2715; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2716; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2717; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2718; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2719; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2720; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2721; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2722; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2723; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2724; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2725; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd2726; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2727; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2728; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd2729; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd2730; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2731; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2732; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2733; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2734; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2735; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2736; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2737; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2738; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2739; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2740; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2741; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2742; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2743; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2744; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2746; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2747; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2748; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2749; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2750; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2751; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2752; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2753; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2754; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2755; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2756; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2757; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2758; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2759; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2760; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2761; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2762; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2763; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2764; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2765; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2766; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd2767; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2768; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2769; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2770; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2771; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2773; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2774; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2775; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2776; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2777; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2778; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2779; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2780; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2781; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2782; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2783; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2784; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2785; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2786; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2787; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2788; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2789; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2790; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2791; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd2792; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2793; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2794; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd2795; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2796; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2797; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2798; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2799; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2800; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2801; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2802; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2803; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2804; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2805; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2806; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2807; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2808; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2809; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2810; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2811; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2812; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2813; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2814; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd2815; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2816; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2817; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2818; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2819; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd2820; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2822; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2823; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2824; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2825; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2826; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2827; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2828; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2829; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2830; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2831; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2832; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2833; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2834; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2835; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2836; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2837; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2838; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd2839; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2840; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd2841; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2842; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2843; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2844; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2845; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2846; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd2847; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd2848; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd2849; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2850; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2851; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd2852; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2853; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2854; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2855; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2856; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2857; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2858; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2859; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2860; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2861; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2862; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2863; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2864; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd2865; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2866; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2867; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2868; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd2869; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2870; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd2871; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2872; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2873; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2874; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd2875; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd2876; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2877; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2878; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2879; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2880; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2881; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2882; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2883; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2884; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2885; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd2886; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2887; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2888; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2889; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2890; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2891; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2892; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd2893; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2894; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2895; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2896; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2897; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2898; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2899; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2900; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2901; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2902; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd2903; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2904; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2905; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd2906; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2907; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2908; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2909; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2910; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2911; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2912; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2914; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2915; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2916; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2917; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2918; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2919; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd2920; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2921; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd2922; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2923; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2924; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2925; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2926; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2927; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2928; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2929; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd2930; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2931; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd2932; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2933; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2934; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd2935; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2936; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2937; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2938; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2939; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2940; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2941; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2942; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2943; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2944; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2945; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2946; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2947; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2948; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd2949; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2950; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2951; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd2952; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2953; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2954; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd2955; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd2956; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2957; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2958; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2959; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2960; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2961; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2962; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2963; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2964; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2965; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2966; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2967; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2968; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2969; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2970; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2971; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2972; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2973; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2974; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd2975; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd2976; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd2977; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2978; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd2979; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd2980; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd2981; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2982; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2983; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd2984; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd2985; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd2986; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd2987; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd2988; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2989; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2990; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2991; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd2993; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2994; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2995; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2996; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd2997; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd2998; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd2999; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3000; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3001; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3002; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd3003; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd3004; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3005; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3006; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3007; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3008; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd3009; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3010; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3011; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3012; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3013; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3014; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3015; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3016; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3017; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3018; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3019; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3020; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3021; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3022; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3023; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3024; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3025; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3026; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3027; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3028; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3029; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3030; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd3031; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3032; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3033; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3034; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3035; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3036; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3037; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd3038; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3039; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3040; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3042; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3043; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3044; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3045; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3046; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3047; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3048; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3049; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3050; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3051; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3052; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3053; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3054; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3055; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3056; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3057; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3058; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3059; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd3060; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3062; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3063; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3064; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3065; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd3066; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3067; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3068; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3069; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3070; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3071; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3072; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3073; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3074; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3076; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3077; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3078; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3079; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3080; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3081; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3082; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3083; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3084; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3085; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3086; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3087; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd3088; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3089; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3090; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3091; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3092; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3093; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd3094; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3095; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3096; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3097; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd3098; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3099; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3100; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3101; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3102; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3103; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3104; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3105; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3106; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3107; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3108; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3109; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3110; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3111; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3112; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3113; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3114; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3115; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3116; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3117; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3118; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3119; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3120; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3121; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3122; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd3123; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3124; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3125; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3126; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3127; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3128; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3129; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3130; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3131; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3132; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3133; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3134; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3135; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3136; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3137; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3138; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3139; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3140; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3141; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3142; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3143; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3144; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3145; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3146; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3147; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3148; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd3149; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3150; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3151; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3152; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3153; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3154; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3155; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3156; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3158; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3159; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3160; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3161; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3162; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3163; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3164; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3165; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3166; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3167; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3168; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3169; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3170; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3171; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd3172; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3173; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3174; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd3175; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd8;
#10 addr = 20'd3176; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd3177; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3178; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3179; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3180; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3181; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3182; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3183; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3184; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3186; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3187; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3189; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3190; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3191; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3192; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3193; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3194; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3195; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3196; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3197; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd3198; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3199; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd3200; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3201; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3202; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd3203; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3204; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd3205; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3206; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd3207; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3208; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3209; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3210; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3211; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3212; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3213; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3214; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3215; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3216; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3217; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3218; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3219; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3220; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3221; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3222; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3223; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3224; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3225; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd3226; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd3227; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd3228; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3229; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3230; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3231; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd3232; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd3233; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3234; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd3235; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3236; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3237; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3238; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3239; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3240; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3241; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3242; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3243; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3244; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3245; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3246; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3247; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3249; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3250; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3251; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3252; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3253; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd3254; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3255; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd3256; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd3257; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3258; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3259; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3260; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd3261; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3262; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd11;
#10 addr = 20'd3263; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3264; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3265; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3266; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3267; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3268; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3269; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3270; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3271; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3272; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3273; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3274; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3275; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3277; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3278; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3279; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3280; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3281; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd3282; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3283; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3284; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3285; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3286; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3287; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd3288; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3289; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3290; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd12;
#10 addr = 20'd3291; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3292; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3293; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3294; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3295; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3296; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3297; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3298; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3299; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3300; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3301; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3302; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3303; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3304; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3305; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3306; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3307; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3308; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3309; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd3310; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3311; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3312; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd3313; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3314; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3315; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3316; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd3317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3318; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd3319; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3320; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3321; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3322; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3323; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3324; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3325; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3328; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3329; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3330; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3331; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3333; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3334; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3335; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3336; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3337; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3338; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3339; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3340; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3341; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3342; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3343; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd3344; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3345; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3346; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd3347; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3348; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3349; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3350; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3351; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd3352; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3353; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3354; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3355; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3356; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3357; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3358; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3359; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3360; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3361; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3362; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3363; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3364; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3365; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3366; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3367; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3368; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd3369; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3370; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3371; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd3372; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd3373; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3374; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3375; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3376; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3377; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3378; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3379; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3380; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3381; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3382; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3383; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3384; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3385; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3386; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3387; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3389; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3390; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3391; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3392; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3393; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3394; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd3395; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3396; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd3397; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3398; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3399; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3400; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3401; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3402; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3403; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3404; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3405; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3406; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3407; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3408; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3409; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3410; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3411; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3412; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3413; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3414; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3415; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3416; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3417; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3418; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3419; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3420; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd3421; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3422; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd3423; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3424; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3425; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3426; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3427; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd3428; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3429; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3430; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3431; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3432; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3433; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3434; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3435; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3436; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3437; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3438; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3439; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3440; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3441; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3442; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3443; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3444; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3445; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3446; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3447; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3448; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd3449; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3450; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3451; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3452; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3453; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3454; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3455; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3456; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3457; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3458; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3459; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3460; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3461; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3462; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3463; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3464; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3465; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3466; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3467; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3468; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3469; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3470; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3471; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3472; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3473; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3474; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3475; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3476; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3477; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3478; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3479; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3480; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3481; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3482; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3484; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3485; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3486; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3487; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3488; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3489; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3490; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3491; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3492; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3493; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3494; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3495; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3496; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3497; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3498; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3499; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3500; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3501; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3502; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3503; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3504; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3505; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3506; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3507; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3508; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd3509; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3510; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3511; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd3512; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3513; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3514; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd3515; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3516; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3517; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3518; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3519; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3520; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3521; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3522; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3523; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3524; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3525; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3526; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3527; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3528; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3529; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3530; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3531; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3532; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3533; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd3534; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3535; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3536; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3537; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd3538; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd3539; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd3540; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3541; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3542; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd3543; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3544; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd3545; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3546; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3547; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3548; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3549; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3550; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3551; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3552; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3553; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3554; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3555; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3556; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3557; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3558; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3559; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3560; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3561; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3562; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3563; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3564; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd3565; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3566; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd3567; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd3568; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3569; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3570; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3571; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3572; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd3573; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3574; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3575; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3576; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3577; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3579; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3580; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3581; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3582; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3583; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3584; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3585; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3586; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3588; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3589; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3590; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3591; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3592; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd3593; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3594; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3595; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd3596; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3597; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3598; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3599; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3600; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd3601; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3602; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3603; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3604; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3605; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3607; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3608; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3609; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3610; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3611; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3612; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3613; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3614; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3615; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3616; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3617; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3618; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3619; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3620; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3621; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3622; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3623; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd3624; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3625; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3626; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3627; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3628; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd3629; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3630; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3631; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3632; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3633; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3634; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3636; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3637; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3638; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3639; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3640; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3641; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3642; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3643; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3644; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3645; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3646; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd3647; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3648; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3649; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3650; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3651; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3652; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3653; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3654; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3655; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3656; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3657; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3658; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3659; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3661; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3662; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3663; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3664; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3665; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3666; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3667; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3668; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3669; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3670; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3671; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3672; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3673; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3674; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd3675; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3676; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3677; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd3678; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3679; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3680; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3681; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3682; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3684; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3685; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3686; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3687; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3688; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3689; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3690; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3691; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3692; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3693; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3694; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3695; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3696; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3697; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3698; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3699; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3700; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3701; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd3702; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd3703; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3704; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3705; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd3706; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3707; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3708; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3709; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3710; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3712; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd3713; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3714; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3715; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3716; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3717; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3718; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3719; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3720; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3721; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3722; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3723; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3724; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3725; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3726; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3727; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3728; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd3729; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3730; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd3731; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3732; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3733; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3734; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd3735; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3736; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3737; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3738; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3739; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3740; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3741; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3742; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3743; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3744; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3745; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3746; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3747; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3748; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3749; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3750; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3751; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3752; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3753; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3754; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3755; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3756; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3757; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd3758; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd3759; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3760; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3761; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3762; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd3763; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3764; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3765; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3766; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3767; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3768; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3769; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3770; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3771; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3772; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3773; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3774; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3775; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3776; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3777; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3778; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3779; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3780; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3781; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3782; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3783; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3784; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3785; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3786; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3787; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3788; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3789; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3790; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd3791; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3792; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3793; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3794; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3795; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3796; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd3797; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3798; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3799; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3800; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd3801; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3802; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3803; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3804; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3805; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3806; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3807; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd3808; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3809; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3810; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3811; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3812; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3813; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3814; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd3815; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3816; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd3817; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3818; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd3819; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3820; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3821; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3822; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3823; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3824; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd3825; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3826; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3827; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3828; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3829; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3830; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3831; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3832; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3833; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3834; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3835; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3836; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3837; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3838; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3839; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3840; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd3841; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3842; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd3843; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3844; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3845; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3846; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd3847; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3848; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3849; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3850; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3851; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3852; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3853; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3854; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3855; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3856; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3857; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3858; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3859; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3860; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3861; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3862; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3863; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3864; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3865; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3866; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3867; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3868; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd3869; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3870; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd11;
#10 addr = 20'd3871; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3872; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3873; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3874; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3875; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3876; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3877; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3878; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3879; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3880; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3881; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3882; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3883; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3884; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3885; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3886; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3887; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3888; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3889; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3890; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3891; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3892; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3893; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3894; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3895; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3896; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3897; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3898; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd3899; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3900; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3901; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3902; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd3903; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3904; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3905; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3906; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3907; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3908; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3909; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3910; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3911; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3912; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3913; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3914; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3915; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3917; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3918; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3919; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3920; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3921; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3922; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3923; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3924; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3925; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3926; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd3927; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3928; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3929; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd3930; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd3931; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3932; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3933; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3934; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3935; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3936; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3937; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3938; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3939; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3940; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3941; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3942; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3943; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3944; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3945; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3946; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd3947; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3948; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3949; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd3950; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd3951; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3952; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3953; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3954; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd3955; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3956; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd3957; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd3958; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3959; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3960; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3961; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3962; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3963; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd3964; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3965; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3966; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3967; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3968; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd3969; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3970; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3971; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3972; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3973; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3974; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3975; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd3976; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd3977; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd3978; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd3979; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd3980; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd3981; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd3982; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd3983; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd3984; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd3985; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd3986; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd3987; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd3988; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3989; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3990; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3991; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd3992; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd3993; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd3994; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd3995; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd3996; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd3997; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3998; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd3999; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4000; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4001; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4002; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4003; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4004; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4005; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4006; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4007; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4008; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4009; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4010; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4011; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4012; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4013; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4014; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4015; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4016; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4017; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4018; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4019; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4020; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4021; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4022; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4023; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4024; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd4025; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4026; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4027; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4028; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4029; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4030; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4031; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4032; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4033; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4034; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4035; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4036; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4037; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd4038; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4039; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4040; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4041; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4042; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd4043; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4044; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4045; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4046; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4047; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4048; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4049; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4050; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4051; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4052; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd4053; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4054; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4055; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4056; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4057; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4058; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4059; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4060; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4062; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4063; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4064; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd4065; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd4066; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4067; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4068; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4069; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4070; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4071; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4072; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4073; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4074; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4076; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd4077; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4078; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4079; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4080; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4081; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4082; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4083; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4084; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4085; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4086; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4087; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4088; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4089; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4090; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4091; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4092; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4093; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4094; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4095; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4096; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4097; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4098; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4099; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4100; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4102; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4103; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4104; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4105; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4106; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4107; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4108; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4109; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4110; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4111; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4112; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4113; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4114; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4115; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4116; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4117; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4118; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4119; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4120; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4121; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4122; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4123; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd4124; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd4125; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4126; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4127; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4128; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4129; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4130; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4131; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4132; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4133; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4135; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4136; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4137; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4138; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4139; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4140; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4141; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4142; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4143; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4144; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4145; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4146; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4147; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4148; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4149; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4150; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4151; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd4152; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd4153; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd4154; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4155; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4156; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4157; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4158; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4159; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4160; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd4161; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4162; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4163; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4164; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4165; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4166; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4167; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4168; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4169; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4170; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4171; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4172; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4173; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4174; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4175; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4176; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4177; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4178; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd4179; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4180; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4181; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd4182; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4183; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4184; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4185; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4186; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4187; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4189; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4190; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4191; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4192; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4193; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4194; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4195; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4196; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4197; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4198; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4199; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4200; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4201; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4202; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4203; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4204; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4205; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4206; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4207; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd4208; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4209; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd4210; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4211; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4212; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4213; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4214; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4215; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4216; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4217; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4218; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4219; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4220; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4221; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4222; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4223; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4224; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4225; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4226; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4227; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4228; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4229; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4230; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4231; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4232; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4233; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4234; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4235; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd4236; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4237; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd2;
#10 addr = 20'd4238; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4239; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4240; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4241; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4242; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4243; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4244; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4245; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4246; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4247; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4248; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4249; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4250; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4251; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4252; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4253; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4254; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4255; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4256; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4257; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4258; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4259; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4260; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4261; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4262; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4263; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4264; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd4265; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4266; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4267; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4268; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4269; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4271; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4272; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4273; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4274; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4275; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4276; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4277; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4278; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4279; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4280; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4281; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4282; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4283; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4284; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4285; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4286; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4287; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd4288; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4289; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4290; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4291; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4292; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd4293; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd4294; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4295; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4296; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4298; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd4299; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4300; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4301; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd4302; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4303; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4304; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4305; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4306; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4307; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4308; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4309; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4310; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4311; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4312; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4313; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4314; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4315; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd4316; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4318; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4319; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4320; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd4321; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4322; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4323; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4324; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4325; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4327; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4328; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4329; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4330; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4331; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4332; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4333; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4334; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4335; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4336; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4337; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4338; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4339; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4340; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4341; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4342; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4343; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd4344; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4345; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4346; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4347; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4348; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd4349; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4350; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4351; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4352; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4353; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4354; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4355; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4356; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd4357; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4358; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4359; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4360; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4361; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4362; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4363; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4364; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4365; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4366; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4367; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4368; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4369; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4370; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4371; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4372; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4373; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd4374; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4375; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4376; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4377; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4378; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4379; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4380; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4383; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4384; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd4385; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4386; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4387; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4388; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4389; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4390; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4391; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4392; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4393; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4394; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4395; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4396; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4397; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4398; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4399; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4400; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4401; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4402; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4403; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd4404; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4405; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4406; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4407; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4408; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4411; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4412; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4413; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4414; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4415; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4416; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4417; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4418; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4419; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4420; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4421; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4422; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4423; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4424; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4425; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4426; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4427; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4428; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd4429; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4430; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4431; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4432; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4433; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4434; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4435; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4436; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4437; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4438; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4440; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4441; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4442; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4443; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4444; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4445; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4446; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4447; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4448; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4449; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4450; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd4451; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4452; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4453; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4454; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4455; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4456; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd4457; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4458; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4459; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4460; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4461; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4462; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4463; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4464; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4465; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4466; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4468; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4469; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4470; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4471; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4472; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4473; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4474; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4475; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4476; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4477; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4478; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4479; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4480; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4481; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4482; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4483; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4484; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd4485; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4486; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd4487; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4488; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4489; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4490; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4491; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd4492; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4493; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4495; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4496; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4497; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4498; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4499; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4500; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4501; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4502; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4503; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4504; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4505; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4506; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4507; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4508; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4509; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4510; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4511; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4512; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd4513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4514; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd4515; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4516; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd4517; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4518; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4519; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4520; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4521; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4524; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4525; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4526; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4527; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4528; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4529; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4530; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4531; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4532; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4533; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4534; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4535; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4536; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4537; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4538; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4539; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4540; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4541; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4542; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4543; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4544; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4545; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4546; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4547; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4548; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4549; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4551; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4552; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4553; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4554; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4555; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4556; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4557; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4558; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4559; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4560; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4561; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4562; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4563; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4564; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4565; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4566; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4567; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4568; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4569; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4570; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4571; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4572; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4573; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4574; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4575; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4576; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4577; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4579; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4580; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4581; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4582; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4583; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4584; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4585; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4586; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4588; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd4589; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4590; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4591; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4592; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4593; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4594; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4595; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4596; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4597; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4598; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4599; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4600; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4601; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4602; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4603; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4604; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4605; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4607; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4608; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4609; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4610; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4611; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4612; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4613; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4614; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4615; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4616; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4617; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4618; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4619; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4620; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4621; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4622; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4623; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4624; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4625; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4626; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd4627; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4629; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4630; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4631; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4632; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4633; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4636; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4637; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4638; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4639; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4640; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4641; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4642; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4643; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4644; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4645; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4646; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4647; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4648; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4649; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4650; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4651; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4652; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4653; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4654; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd4655; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4656; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4657; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4658; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4659; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4661; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4663; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4664; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4665; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4666; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4667; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4668; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4669; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4670; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4671; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4672; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4673; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4674; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4675; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4676; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4677; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4678; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4679; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4680; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4682; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4684; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4685; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4686; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4687; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4688; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4689; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4690; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4691; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4692; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4693; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4694; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4695; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4696; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4697; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4698; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4699; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4700; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4701; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4702; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4703; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4704; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4705; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4706; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd4707; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd8;
#10 addr = 20'd4708; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4709; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4710; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd4712; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4713; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4714; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4715; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4716; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4717; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4718; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4719; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4720; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4721; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4722; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4723; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4724; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4725; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4726; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4727; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4728; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4729; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4730; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4731; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4732; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4733; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4734; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4735; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4736; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4737; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4738; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4739; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd4740; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4741; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4742; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4743; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4744; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4745; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4746; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4747; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4748; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4749; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4750; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4751; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4752; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4753; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4754; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4755; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4756; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4757; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4758; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4759; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4760; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4761; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4762; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4763; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd4764; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4765; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4766; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4767; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4768; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd4769; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4770; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4771; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4772; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4773; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4774; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4775; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4776; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd4777; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4778; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4779; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4780; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4781; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4782; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4783; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4784; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4785; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4786; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4787; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4788; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4789; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4790; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4791; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4792; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4793; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4794; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4795; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4796; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd4797; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4798; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4799; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4800; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4801; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4802; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4803; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4804; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4805; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4806; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4807; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4808; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4809; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4810; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4811; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4812; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd4813; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4814; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4815; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4816; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4817; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4818; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4819; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4820; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4822; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd4823; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4824; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4825; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4826; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4827; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4828; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4829; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4830; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4831; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4832; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd4833; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd4834; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4835; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4836; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4837; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4838; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4839; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4840; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4841; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4842; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4843; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4844; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4845; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4846; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4847; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4848; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4849; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4850; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd4851; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4852; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd4853; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4854; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4855; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4856; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4857; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4858; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4859; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4860; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4861; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd4862; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4863; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4864; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4865; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4866; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4867; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4868; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4869; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4870; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4871; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4872; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4873; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4874; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd4875; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd4876; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4877; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd4878; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4879; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4880; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd4881; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4882; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4883; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4884; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4885; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4887; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4888; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4889; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd4890; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4891; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4892; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4893; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4894; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4895; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4896; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4897; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4898; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4899; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd4900; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4901; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4902; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4903; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd4904; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4905; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd4906; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4907; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd4908; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd4909; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4910; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4911; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4912; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4913; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4914; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4915; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4917; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4918; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4919; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4920; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4921; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4922; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4923; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4924; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4925; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4926; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4927; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4928; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd4929; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4930; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4931; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd4932; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd4933; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd4934; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd4935; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4936; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd4937; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4938; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4939; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4940; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4941; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4942; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4943; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4944; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4945; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4946; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd4947; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4948; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd4949; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4950; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4951; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4952; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4953; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd4954; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4955; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4956; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4957; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4958; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4959; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4960; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd4961; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd4962; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd4963; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd4964; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd4965; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4966; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4967; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4968; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4969; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4970; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4971; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4972; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd4973; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd4974; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4975; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd4976; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4977; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4978; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4979; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4980; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd4981; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd4982; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4983; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4984; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd4985; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4986; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd4987; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd4988; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd4989; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd4990; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd4991; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd4992; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd4993; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4994; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4995; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd4996; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd4997; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4998; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd4999; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5000; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5001; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5002; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd5003; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5004; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5005; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5006; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5007; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5008; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5009; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd5010; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5011; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5012; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5013; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5014; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5015; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5016; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5017; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5018; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd5019; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5020; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd5021; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5022; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5023; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5024; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5025; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5026; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5027; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5028; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5029; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5030; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd5031; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5032; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5033; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5034; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5035; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5036; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5037; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5038; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5039; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5040; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5041; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5042; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5043; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd5044; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5045; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5046; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd5047; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd5048; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd5049; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5050; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5051; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5052; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5053; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5054; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5055; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5056; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5057; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5058; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd5059; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5060; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5061; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5062; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5063; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5064; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5065; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5066; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5067; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5068; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5069; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5070; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5071; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd5072; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5073; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5074; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd5075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd5076; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5077; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5078; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5079; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5080; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5081; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5082; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5083; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5084; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5085; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5086; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5087; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5088; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5089; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5090; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5091; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5092; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5093; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5094; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5095; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5096; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5097; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5098; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5099; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5100; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5101; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd5102; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5103; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd5104; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5105; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd5106; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5107; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5108; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5109; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5110; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5111; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5112; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5113; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5114; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5115; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5116; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5117; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5118; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5119; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5120; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5121; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5122; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5123; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5124; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5125; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5126; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5127; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5128; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd5129; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd5130; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd5131; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5132; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd5133; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd5134; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5135; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5136; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5137; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5138; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5139; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5140; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5141; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5142; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5143; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5144; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5145; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5146; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5147; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5148; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5149; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5150; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5151; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5152; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5153; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5154; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5155; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd5156; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd5158; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5159; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5160; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd5161; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd3;
#10 addr = 20'd5162; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5163; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5164; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5165; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5166; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5167; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5168; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5169; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5170; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5171; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5172; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5173; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5174; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5175; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5176; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5177; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5178; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5179; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5180; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5181; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5182; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5183; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5184; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd5186; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5187; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5188; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd5189; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd3;
#10 addr = 20'd5190; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5191; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5192; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5193; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5194; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5195; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5196; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5197; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5198; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5199; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5200; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5201; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5202; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5203; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5204; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5205; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5206; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5207; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5208; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5209; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5210; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5211; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5212; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5213; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd5214; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd5215; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5216; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5217; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd3;
#10 addr = 20'd5218; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5219; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5220; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5221; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5222; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5223; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5224; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5225; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5226; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5227; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5228; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5229; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5230; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5231; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5232; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5233; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5234; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5235; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5236; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5237; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5238; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5239; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5240; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5241; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd5242; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5243; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5244; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5245; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd5246; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5247; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5248; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5249; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5250; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5251; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5252; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5253; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5254; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5255; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd5256; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5257; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5258; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5259; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5260; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5261; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5262; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5263; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5264; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5265; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5266; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5267; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5268; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5269; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd5270; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5271; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5272; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd5273; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd5274; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5275; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5276; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5277; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5278; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5279; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5280; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5281; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5282; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5283; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5284; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5285; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5286; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5287; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5288; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5289; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5290; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5291; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5292; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5293; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5294; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5295; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5296; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5297; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5298; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5299; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5300; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5301; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5302; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5303; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5304; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5305; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5306; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5307; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5308; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5309; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5310; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5311; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5312; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5313; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5314; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5315; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5316; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5317; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5318; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5319; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5320; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5321; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5322; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5323; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5324; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5325; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5326; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5327; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd5328; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd5329; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd5330; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5331; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5332; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5333; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5334; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5335; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5336; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5337; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5338; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5339; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd5340; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5341; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5342; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5343; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5344; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5345; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5346; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5347; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5348; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5349; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5350; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5351; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5352; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5353; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5354; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5355; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd5356; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5357; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5358; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5359; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5360; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5361; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5362; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5363; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5364; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5365; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5366; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5367; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd5368; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5369; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5370; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5371; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5372; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5373; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5374; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5375; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5376; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5377; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5378; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5379; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5380; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5381; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5382; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5383; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5384; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd5385; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5386; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5387; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5389; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5390; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5391; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5392; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5393; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5394; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5395; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd3;
#10 addr = 20'd5396; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5397; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5398; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5399; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5400; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5401; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5402; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5403; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5404; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5405; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5406; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5407; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5408; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5409; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5410; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5411; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5412; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd5413; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5414; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5415; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5416; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5417; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5418; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5419; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5420; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5421; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5422; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5423; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd5424; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5425; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5426; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5427; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5428; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5430; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5431; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5432; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5433; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5434; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5435; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5436; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5438; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5439; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5440; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd5441; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5442; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5443; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5444; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5445; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5446; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5447; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5448; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5449; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5450; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5451; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd5452; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5453; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5454; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5455; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5456; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd5457; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5458; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5459; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5460; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5461; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5462; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5463; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5464; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5465; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5466; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5467; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5468; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5469; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd5470; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5471; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5472; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5473; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5474; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5475; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5476; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5477; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5478; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5479; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd5480; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5481; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5482; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5483; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5484; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5485; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5486; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5487; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5488; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5489; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5490; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5491; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5492; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5493; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5494; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5495; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd5496; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5497; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5498; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5499; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5500; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5501; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5502; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5503; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5504; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5505; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5506; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5507; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd5508; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5509; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5510; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5511; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5512; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5514; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5515; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5516; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5517; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5518; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5519; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5520; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5521; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5522; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5523; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5524; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5525; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5526; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5527; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5528; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5529; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5530; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5531; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5532; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5533; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5534; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5535; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5536; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5537; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5538; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5539; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd5540; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5542; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5543; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5544; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5545; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5546; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5547; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5548; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5549; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5550; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5551; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd5552; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5553; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5554; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5555; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5556; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd5557; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5558; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5559; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5560; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5561; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5562; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5563; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5564; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5565; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5566; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5567; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5568; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5569; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5570; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5571; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5572; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5573; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5574; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5575; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5576; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5577; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5578; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5579; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd5580; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5581; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd5582; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5583; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5584; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5585; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5586; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5587; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5588; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5589; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5590; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5591; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd5592; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5593; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5594; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5595; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5596; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5597; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5598; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5599; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5600; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5601; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5602; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5603; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5604; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5605; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5606; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5607; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd5608; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd5609; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5610; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5611; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5612; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5613; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5614; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5615; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5616; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5617; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5618; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5619; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5620; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5621; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5622; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5623; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd5624; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5625; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5626; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5627; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5628; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5629; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5630; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5631; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5632; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5633; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5635; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5636; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd5637; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5638; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5639; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5640; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5641; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5642; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5643; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5644; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5645; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5646; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5647; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5648; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5649; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5650; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5651; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd5652; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5653; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5654; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5655; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5656; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5657; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5658; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5659; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5661; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5663; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd5664; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5665; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5666; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5667; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5668; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5669; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5670; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5671; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5672; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5673; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5674; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5675; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5676; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5677; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5678; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5679; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5680; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5682; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5683; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5684; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5685; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5686; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5687; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5688; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5689; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5690; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5691; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd5692; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5693; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5694; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5695; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5696; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5697; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5698; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5699; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5700; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5701; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5702; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd5703; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd5704; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5705; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5706; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5707; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd5708; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5709; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5710; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5711; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5712; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5713; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5714; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5715; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5716; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5717; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5718; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5719; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd5720; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd5721; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5722; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5723; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5724; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5725; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5726; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5727; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5728; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5729; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5730; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd5731; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd5732; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5733; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5734; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd5735; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5736; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5737; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5738; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5739; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5740; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5741; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5742; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5743; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5744; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5746; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5747; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5748; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5749; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5750; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5751; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5752; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5753; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5754; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5755; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5756; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5757; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5758; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5759; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd5760; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5761; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5762; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5763; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd5764; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5765; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5767; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5768; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5769; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5770; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5771; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5772; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5773; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5774; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5775; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd5776; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5777; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5778; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5779; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5780; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5781; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5782; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5783; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5784; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5785; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5786; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5787; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd5788; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5789; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5790; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5791; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5792; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5793; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5795; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5796; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd5797; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5798; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5799; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5800; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5801; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5802; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5803; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5804; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5805; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5806; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5807; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5808; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5809; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5810; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5811; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5812; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5813; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5814; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5815; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd5816; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5817; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5818; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd5819; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5820; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5822; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5823; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5824; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5825; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5826; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5827; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5828; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5829; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5830; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5831; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5832; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5833; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5834; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5835; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5836; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5837; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5838; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5839; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5840; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5841; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5842; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5843; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5844; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5845; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5846; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd5847; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5848; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5849; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5850; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5851; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5852; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5853; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5854; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5855; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5856; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5857; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5858; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5859; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5860; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5861; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5862; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5863; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd5864; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5865; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5866; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5867; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5868; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5869; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd5870; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5871; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5872; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5873; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5874; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd5875; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd5876; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5877; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5878; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5879; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5880; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5881; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5882; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5883; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5884; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5885; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5887; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5888; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd5889; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5890; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5891; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5892; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5893; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5894; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5895; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5896; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5897; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5898; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5899; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd5900; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5901; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5902; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5903; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5904; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5905; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5906; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5907; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5908; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd5909; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5910; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5911; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5912; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5913; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5914; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5915; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5917; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5918; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5919; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd5920; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5921; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5922; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5923; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5924; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5925; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5926; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd5927; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd5928; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5929; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5930; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5931; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd5932; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5933; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5934; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5935; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5936; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5937; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5938; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5939; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5940; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5941; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd5942; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5943; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5944; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5945; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5946; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5947; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5948; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5949; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5950; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5951; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5952; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5953; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5954; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5955; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd5956; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5957; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5958; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5959; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5960; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5961; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5962; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5963; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5964; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5965; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5966; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5967; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5968; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd5969; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5970; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd5971; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd5972; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5973; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd5974; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5975; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5976; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd5977; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5978; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5979; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5980; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5981; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5982; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd5983; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd5984; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5985; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5986; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd5987; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5988; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5989; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5990; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd5991; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5992; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd5993; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5994; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd5995; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd5996; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd5997; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd5998; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd5999; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd6000; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd6001; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6002; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6003; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6004; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6005; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6006; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6007; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6008; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6009; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6010; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6011; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd6012; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6013; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6014; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6015; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6016; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6017; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6018; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6020; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd6021; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6022; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6023; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6024; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6025; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6026; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd6027; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd6028; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd6029; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6030; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6031; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6032; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6033; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6034; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6035; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6036; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6037; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6038; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6039; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd6040; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6041; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6042; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6043; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6044; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6045; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6046; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6047; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6048; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd6049; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6050; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6051; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6052; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6053; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6054; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd6055; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6056; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6057; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6058; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6059; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6060; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6061; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6062; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6063; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6064; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6065; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6066; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6067; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6068; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6069; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6070; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6071; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6072; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6073; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6074; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6075; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6076; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd6077; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6078; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6079; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6080; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6081; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd6082; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd6083; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6084; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6085; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6086; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6087; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6088; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6089; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6090; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6091; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6092; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6093; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6094; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6095; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6096; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6097; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6098; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6099; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6100; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6102; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6103; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6104; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd6105; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6106; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6107; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6108; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6109; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd6110; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6111; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd6112; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd6113; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6114; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6115; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6116; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6117; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6118; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6119; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6120; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6121; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6122; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6123; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6124; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6125; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6126; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6127; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6128; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6129; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6130; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6131; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6132; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd6133; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6135; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6136; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6137; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd6138; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd6139; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd6140; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd6141; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6142; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6143; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6144; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6145; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6146; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6147; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6148; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6149; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6150; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6151; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6152; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd6153; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6154; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6155; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6156; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6158; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6159; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6160; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd6161; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6162; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6163; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6164; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6165; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd6166; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd6167; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6168; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6169; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6170; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6171; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6172; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6173; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6174; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6175; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6176; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6177; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6178; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6179; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6180; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd6181; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6182; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6183; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6184; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6186; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6187; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6188; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd6189; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6190; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6191; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6192; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6193; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd6194; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6195; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6196; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6197; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6198; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6199; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6200; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6201; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6202; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6203; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6204; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6205; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6206; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6207; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6208; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd6209; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6210; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6211; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6212; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6213; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6214; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6215; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6216; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd6217; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6218; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6219; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6220; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6221; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd6222; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6223; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6224; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6225; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6226; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6227; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6228; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6229; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6230; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6231; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6232; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6233; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6234; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6235; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd6236; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd6237; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6238; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6239; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6240; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6241; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6242; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6243; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6244; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd6245; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6246; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6247; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6248; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6249; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd6250; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd6251; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6252; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd6253; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd6254; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6255; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6256; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6257; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6258; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6259; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6260; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6261; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6262; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6263; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd6264; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd6265; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6266; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6267; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6268; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6269; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6270; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6271; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6272; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6273; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6274; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6275; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6276; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6277; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6278; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6279; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6280; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6281; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6282; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6283; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6284; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6285; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6286; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6287; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6288; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6289; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6290; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6291; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6292; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6293; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6294; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd6295; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6296; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6298; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6299; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd6300; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6301; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6302; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6303; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6304; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6305; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6306; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6307; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6308; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6309; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6310; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6311; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6312; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6313; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6314; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6315; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6316; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6318; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6319; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6320; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6321; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6322; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd6323; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6324; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6325; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6326; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6327; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd6328; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6329; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6330; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6331; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd6332; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6333; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6334; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6335; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6337; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6338; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6339; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6340; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6341; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6342; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6343; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6344; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6346; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6347; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6348; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6349; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6350; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd6351; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6352; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6353; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6354; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6355; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd6356; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6357; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6358; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6359; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6360; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6361; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6362; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6363; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6364; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6365; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6366; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6367; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6368; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6369; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6370; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6371; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6372; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6374; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6375; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6376; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6377; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6378; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6379; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6382; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6383; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6384; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6385; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6386; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6387; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6388; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6389; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6390; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6391; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6392; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6393; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6394; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6395; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6396; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6397; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6398; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6399; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6400; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6402; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6403; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6404; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6405; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6406; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6407; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6410; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6411; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6412; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6413; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6414; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6415; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6416; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6417; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6418; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6419; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6420; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6421; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6422; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6423; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6424; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6425; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6426; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6427; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6428; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6430; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6431; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6432; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6433; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6434; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6435; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6436; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6438; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6440; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6441; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6442; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6443; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6444; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6445; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6446; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6447; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6448; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6449; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6450; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6451; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6452; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6453; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6454; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6455; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6456; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6457; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6459; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6460; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6461; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6462; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6463; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6464; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6465; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6466; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6468; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6469; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6470; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6471; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6472; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6473; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6474; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6475; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6476; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6477; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6478; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6479; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6480; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6481; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6482; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6483; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6484; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6485; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6486; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6487; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6488; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6489; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6490; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd6491; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6492; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6493; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6495; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6496; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6497; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6498; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6499; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6500; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6501; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6502; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6503; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6504; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6505; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6506; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6507; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6508; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6509; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6510; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6511; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6512; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6514; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6515; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6516; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6517; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6518; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd6519; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6520; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6521; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd6523; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6524; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6525; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6526; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6527; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6528; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6529; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6530; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6531; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6532; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6533; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6534; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6535; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6536; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6537; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6538; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6539; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6540; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6542; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6543; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6544; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6545; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6546; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd6547; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6548; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6549; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd6551; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6552; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6553; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6554; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6555; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6556; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6557; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6558; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6559; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6560; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6561; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6562; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6563; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6564; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6565; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6566; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6567; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6568; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6569; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6570; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6571; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6572; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6573; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6574; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd6575; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6576; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6577; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd6579; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6580; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6581; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6582; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6583; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6584; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6585; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6586; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6587; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6588; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6589; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6590; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6591; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6592; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6593; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6594; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6595; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6596; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6597; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6598; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6599; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6600; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6601; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6602; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd6603; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd6604; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6605; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd6607; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6608; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6609; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6610; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6611; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6612; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6613; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6614; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6615; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6616; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6617; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6618; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6619; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6620; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6621; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6622; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6623; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6624; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6625; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6626; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6627; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6629; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6630; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd6631; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd6632; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6633; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6635; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6636; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6637; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6638; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6639; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6640; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6641; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6642; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6643; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6644; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6645; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6646; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6647; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6648; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6649; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6650; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6651; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6652; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6653; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6654; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6655; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6656; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6657; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6658; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd6659; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd6660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6661; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6662; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6663; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd6664; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6665; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6666; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6667; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6668; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6669; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6670; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6671; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6672; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6673; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6674; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6675; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6676; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6677; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6678; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6679; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6680; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6681; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6682; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6684; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6685; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6686; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6687; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd6688; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6689; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6690; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6691; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6692; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6693; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6694; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6695; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6696; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6697; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6698; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6699; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6700; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6701; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6702; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6703; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6704; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6705; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6706; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6707; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6708; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6709; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6710; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6712; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6713; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6714; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6715; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6716; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6717; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6718; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd6719; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6720; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6721; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6722; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6723; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6724; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6725; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6726; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6727; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6728; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6729; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6730; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6731; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6732; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6733; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6734; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6735; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6736; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6737; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6738; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6739; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6740; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6741; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6742; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6743; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6744; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6745; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd6746; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6747; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6748; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6749; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6750; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6751; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6752; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6753; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6754; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6755; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6756; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6757; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6758; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6759; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6760; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6761; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6762; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6763; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6764; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6765; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6766; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6767; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6768; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6769; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6770; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6771; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6772; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6773; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd6774; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd6775; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6776; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd6777; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6778; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6779; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6780; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6781; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6782; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6783; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6784; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6785; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6786; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6787; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6788; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6789; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6790; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6791; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6792; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6793; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6794; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6795; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6796; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6797; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6798; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6799; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6800; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6801; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd6802; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd6803; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6804; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6805; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6806; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6807; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6808; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6809; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6810; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6811; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6812; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6813; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6814; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6815; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6816; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6817; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6818; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6819; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6820; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6821; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6822; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6823; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6824; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6825; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6826; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6827; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6828; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6829; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6830; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd6831; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6832; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6833; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6834; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6835; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6836; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6837; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6838; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6839; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6840; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6841; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6842; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6843; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6844; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd6845; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6846; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6847; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6848; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6849; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6850; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6851; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6852; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6853; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6854; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6855; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6856; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6857; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6858; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd6859; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6860; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6861; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6862; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6863; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6864; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6865; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6866; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6867; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6868; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6869; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6870; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6871; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6872; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd6873; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6874; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6875; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6876; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6877; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6878; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6879; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6880; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6881; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6882; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6883; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6884; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6885; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6886; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd6887; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6888; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6889; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6890; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6891; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6892; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6893; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6894; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6895; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6896; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6897; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6898; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6899; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6900; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd6901; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd6902; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6903; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6904; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6905; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6906; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6907; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6908; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6909; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6910; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd6911; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd6912; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6914; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6915; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6916; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd6917; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6918; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6919; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6920; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6921; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6922; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6923; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd6924; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6925; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6926; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6927; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd6928; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd6929; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6930; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6931; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6932; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6933; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6934; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6935; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6936; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6937; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6938; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6939; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd6940; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6941; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6942; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6943; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6944; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6945; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6946; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6947; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd6948; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6949; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6950; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6951; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6952; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6953; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6954; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6955; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6956; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd6957; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6958; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6959; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6960; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6961; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6962; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6963; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6964; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6965; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6966; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6967; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd6968; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd6969; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6970; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6971; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6972; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd6973; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd6974; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6975; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd6976; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6977; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd6978; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6979; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6980; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6981; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6982; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6983; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd6984; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd6985; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd6986; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd6987; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd6988; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd6989; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd6990; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6991; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6993; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd6994; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd6995; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd6996; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd1;
#10 addr = 20'd6997; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6998; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd6999; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7000; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7001; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7002; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7003; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7004; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7005; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7006; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7007; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7008; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7009; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7010; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7011; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7012; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7013; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7014; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd7015; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7016; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7017; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7018; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7019; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7020; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7021; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7022; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7023; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd7024; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd9;data_in[31:28] = 4'd0;
#10 addr = 20'd7025; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7026; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7027; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7028; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7029; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7030; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7031; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7032; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7033; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7034; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7035; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7036; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7037; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7038; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7039; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd7040; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7042; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7043; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7044; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7045; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7046; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7047; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7048; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7049; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7050; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7051; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd7052; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd5;data_in[31:28] = 4'd0;
#10 addr = 20'd7053; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7054; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7055; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7056; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7057; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7058; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7059; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7060; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7062; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7063; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7064; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7065; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7066; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7067; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7068; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7069; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7070; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7071; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7072; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7073; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7074; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7076; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7077; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7078; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7079; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7080; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7081; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7082; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7083; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7084; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7085; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7086; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7087; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7088; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7089; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7090; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7091; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7092; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd7093; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7094; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7095; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7096; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7097; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7098; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7099; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7100; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7101; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7102; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7103; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7104; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7105; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7106; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7107; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7108; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7109; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7110; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7111; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7112; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd7113; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7114; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7115; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7116; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7117; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7118; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7119; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7120; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7121; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7122; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7123; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7124; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7125; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7126; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7127; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7128; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7129; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7130; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7131; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7132; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7133; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7134; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7135; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7136; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7137; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7138; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7139; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7140; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd7141; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7142; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7143; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7144; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7145; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7146; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7147; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7148; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7149; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7150; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7151; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7152; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7153; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7154; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7155; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7156; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7158; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7159; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7160; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7161; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7162; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7163; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7164; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7165; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7166; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7167; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7168; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7169; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7170; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7171; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7172; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7173; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7174; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7175; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7176; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7177; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7178; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7179; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7180; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7181; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7182; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7183; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd7184; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7186; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7187; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7188; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7189; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7190; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7191; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7192; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7193; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7194; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7195; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd6;
#10 addr = 20'd7196; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7197; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7198; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7199; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7200; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7201; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7202; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7203; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7204; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7205; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7206; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7207; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7208; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7209; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7210; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7211; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7212; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7213; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7214; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7215; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7216; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7217; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7218; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7219; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7220; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7221; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7222; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7223; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd7224; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7225; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7226; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7227; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7228; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7229; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7230; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7231; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7232; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7233; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7234; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7235; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7236; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7237; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7238; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7239; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7240; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7241; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7242; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7243; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7244; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7245; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7246; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7247; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7248; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7249; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7250; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7251; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd7252; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7253; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7254; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7255; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7256; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7257; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7258; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7259; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7260; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7261; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7262; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7263; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7264; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7265; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7266; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7267; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7268; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7269; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7270; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7271; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd7272; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7273; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7274; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7275; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd7276; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7277; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7278; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd7279; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7280; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7281; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7282; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7283; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7284; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7285; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7286; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7287; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7288; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7289; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7290; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7291; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7292; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7293; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd7294; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd7295; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7296; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd8;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd7297; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7298; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7299; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7300; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7301; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7302; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7303; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd1;
#10 addr = 20'd7304; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7305; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7306; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7307; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7308; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7309; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7310; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7311; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7312; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7313; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7314; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7315; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7316; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7318; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7319; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7320; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7321; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7322; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7323; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7324; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7325; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7326; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7328; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7329; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7330; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7331; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd7332; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7333; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7334; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7335; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7336; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7337; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7338; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7339; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7340; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7341; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7342; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7343; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7344; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7346; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7347; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7348; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7349; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7350; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7351; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7352; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7353; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7354; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7355; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7356; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7357; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7358; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7359; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7360; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7361; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7362; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7363; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7364; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7365; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7366; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7367; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7368; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7369; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7370; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7371; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7372; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7374; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7375; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7376; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7377; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7378; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7379; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7380; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd7381; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7382; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7383; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7384; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7385; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7386; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7387; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd7388; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7389; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7390; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7391; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7392; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7393; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7394; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7395; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7396; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7397; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7398; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7399; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7402; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7403; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7404; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7405; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7406; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7407; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd7408; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd2;
#10 addr = 20'd7409; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd7410; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7411; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7412; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7413; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7414; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7415; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd7416; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7417; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7418; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7419; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7420; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7421; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7422; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7423; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7424; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7425; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7426; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7427; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7428; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7430; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7431; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7432; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7433; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7434; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7435; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7436; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd6;
#10 addr = 20'd7437; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7438; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7439; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7440; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7441; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7442; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7443; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7444; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7445; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7446; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7447; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7448; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7449; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7450; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7451; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7452; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7453; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7454; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7455; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7456; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7457; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7459; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7460; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7461; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7462; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7463; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7464; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd7465; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7466; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7467; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7468; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd7469; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7470; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7471; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7472; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7473; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7474; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd7475; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7476; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7477; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7478; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7479; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7480; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7481; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7482; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7484; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7485; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7486; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7487; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7488; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd7489; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7490; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7491; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7492; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd7493; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7494; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7495; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7496; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd7497; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7498; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7499; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7500; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7501; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7502; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7503; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7504; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7505; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7506; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7507; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7508; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7509; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7510; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7511; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7512; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7514; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7515; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7516; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7517; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7518; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7519; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7520; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7521; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7522; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7523; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7524; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd7525; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7526; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7527; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7528; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7529; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7530; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7531; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7532; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7533; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7534; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7535; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7536; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7537; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7538; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7539; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7540; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7542; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7543; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7544; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7545; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7546; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7547; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7548; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7549; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7550; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7551; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7552; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7553; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7554; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7555; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7556; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7557; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7558; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7559; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7560; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7561; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7562; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7563; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7564; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7565; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7566; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7567; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7568; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7569; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7570; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7571; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7572; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7573; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7574; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7575; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7576; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7577; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7578; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7579; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7580; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7581; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7582; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7583; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7584; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7585; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7586; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7588; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7589; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7590; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7591; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7592; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7593; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7594; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7595; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7596; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7597; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7598; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7599; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7600; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7601; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7602; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7603; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7604; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd7605; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7606; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7607; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7608; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7609; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7610; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd7611; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7612; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7613; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7614; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd7615; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7616; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7617; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7618; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7619; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7620; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7621; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7622; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7623; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7624; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7625; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7626; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7627; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd7628; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7629; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7630; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7631; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7632; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd7633; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd7634; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7636; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7637; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd7638; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd1;
#10 addr = 20'd7639; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd7640; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7641; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7642; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7643; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7644; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7645; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7646; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7647; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7648; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7649; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7650; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7651; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7652; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7653; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7654; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7655; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd7656; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7657; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7658; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7659; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7660; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7661; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd7662; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7663; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7664; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7665; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7666; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd7667; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7668; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7669; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7670; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7671; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7672; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7673; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7674; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7675; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7676; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7677; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7678; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd7679; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7680; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7681; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7682; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7683; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7684; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7685; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7686; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7687; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7688; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7689; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd10;data_in[31:28] = 4'd2;
#10 addr = 20'd7690; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7691; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7692; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7693; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd4;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7694; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd7695; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7696; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7697; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd7698; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7699; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7700; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7701; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7702; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7703; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7704; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd7705; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7706; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd7707; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7708; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7709; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7710; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7711; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7712; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7713; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7714; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7715; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7716; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7717; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd5;
#10 addr = 20'd7718; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7719; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7720; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd7721; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7722; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd7723; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7724; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7725; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd7726; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd7727; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7728; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7729; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7730; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7731; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7732; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7733; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7734; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd7735; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7736; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7737; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7738; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7739; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7740; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7741; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7742; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7743; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7744; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7745; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd9;
#10 addr = 20'd7746; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7747; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7748; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd7749; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7750; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd7751; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7752; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7753; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd7754; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7755; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7756; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7757; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7758; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7759; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7760; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7761; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7762; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd12;
#10 addr = 20'd7763; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7764; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7765; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7767; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7768; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7769; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7770; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7771; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7772; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7773; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd7774; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7775; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7776; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd7777; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7778; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd11;data_in[31:28] = 4'd1;
#10 addr = 20'd7779; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7780; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7781; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7782; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7783; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7784; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7785; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7786; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7787; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7788; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7789; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7790; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd13;
#10 addr = 20'd7791; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7792; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7793; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7795; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7796; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7797; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7798; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7799; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7800; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7801; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd7802; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7803; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd7804; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd5;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd7805; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7806; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd2;
#10 addr = 20'd7807; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7808; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7809; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7810; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7811; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7812; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7813; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7814; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7815; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd7816; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7817; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7818; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd7819; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7820; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd7821; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7822; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd7823; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd7824; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7825; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7826; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7827; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7828; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7829; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd7830; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7831; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd7832; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7833; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7834; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd3;
#10 addr = 20'd7835; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7836; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7837; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7838; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7839; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7840; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd7841; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7842; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7843; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7844; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7845; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7846; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7847; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7848; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7849; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd7850; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7851; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7852; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd7853; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7854; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7855; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7856; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7857; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7858; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7859; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7860; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd7861; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7862; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd3;
#10 addr = 20'd7863; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7864; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7865; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd7866; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7867; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7868; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7869; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7870; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7871; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7872; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7873; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7874; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd7875; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7876; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7877; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd7878; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd7879; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd7880; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7881; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7882; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7883; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7884; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7885; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7886; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7887; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd7888; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd7889; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7890; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd2;
#10 addr = 20'd7891; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7892; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7893; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7894; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7895; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7896; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7897; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7898; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7899; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7900; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7901; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7902; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd7903; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7904; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd7905; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7906; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7907; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7908; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7909; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7910; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7911; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7912; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7913; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7914; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7915; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7916; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd7917; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7918; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd2;
#10 addr = 20'd7919; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7920; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7921; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7922; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7923; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7924; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7925; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7926; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7927; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7928; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7929; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7930; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd8;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd7931; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7932; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7933; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7934; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd7935; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7936; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd7937; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7938; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7939; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7940; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7941; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7942; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7943; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd7944; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7945; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7946; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd10;data_in[31:28] = 4'd1;
#10 addr = 20'd7947; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7948; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7949; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7950; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7951; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7952; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7953; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7954; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7955; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7956; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7957; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7958; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd9;data_in[27:24] = 4'd13;data_in[31:28] = 4'd9;
#10 addr = 20'd7959; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7960; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7961; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd7962; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7963; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd7964; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7965; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7966; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7967; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd7968; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd7969; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7970; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7971; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd7972; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7973; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd7974; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd8;data_in[31:28] = 4'd0;
#10 addr = 20'd7975; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd7976; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd7977; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7978; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7979; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd7980; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7981; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7982; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd7983; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd7984; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7985; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd7986; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd8;
#10 addr = 20'd7987; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd7988; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7989; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd7990; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd7991; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7992; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7993; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd7994; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7995; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd7996; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7997; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd7998; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd7999; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8000; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8001; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8002; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd8003; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8004; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8005; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8006; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8007; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8008; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8009; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8010; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8011; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8012; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8013; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8014; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd8015; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8016; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8017; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd8018; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd8019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8020; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8021; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8022; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8023; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8024; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8025; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8026; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd8027; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8028; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8029; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8030; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd5;data_in[31:28] = 4'd0;
#10 addr = 20'd8031; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8032; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8033; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8034; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8035; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8036; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8037; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8038; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8039; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8040; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8041; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8042; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd8043; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8044; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8045; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8046; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8047; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8048; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8049; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8050; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8051; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8052; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8053; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8054; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd8055; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8056; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8057; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8058; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd8059; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8060; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8061; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8062; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8063; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8064; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8065; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8066; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8067; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8068; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8069; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8070; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd8071; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8072; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8073; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8074; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8076; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8077; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8078; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8079; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8080; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8081; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8082; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8083; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8084; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8085; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8086; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd8087; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8088; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd8089; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8090; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8091; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8092; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8093; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8094; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8095; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8096; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8097; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8098; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8099; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8100; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8101; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8102; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8103; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8104; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8105; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8106; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8107; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8108; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8109; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8110; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8111; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8112; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8113; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8114; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd8115; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8116; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd8117; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8118; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8119; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8120; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8121; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8122; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8123; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8124; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8125; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8126; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8127; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8128; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8129; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8130; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8131; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8132; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8133; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8134; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8135; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8136; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8137; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8138; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8139; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8140; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8141; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8142; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd5;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd8143; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8144; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd8145; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8146; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8147; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8148; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8149; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8150; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8151; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8152; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8153; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8154; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8155; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8156; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8158; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8159; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8160; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8161; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8162; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8163; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8164; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8165; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8166; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8167; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8168; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8169; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd8170; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8171; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8172; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8173; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8174; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8175; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8176; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8177; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8178; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8179; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8180; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8181; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8182; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8183; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8184; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8186; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8187; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8189; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8190; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8191; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8192; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8193; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8194; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8195; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8196; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8197; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8198; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd7;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8199; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8200; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8201; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8202; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8203; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8204; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8205; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8206; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8207; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8208; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8209; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8210; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8211; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8212; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8213; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8214; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8215; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8216; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8217; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8218; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8219; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8220; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8221; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8222; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8223; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8224; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8225; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd8226; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8227; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8228; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8229; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8230; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8231; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8232; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8233; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8234; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8235; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8236; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8237; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8238; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8239; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd8240; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd8241; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd8242; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8243; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8244; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8245; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8246; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8247; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8248; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8249; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8250; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8251; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8252; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8253; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8254; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8255; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8256; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8257; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8258; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8259; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8260; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8261; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8262; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8263; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8264; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8265; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8266; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8267; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8268; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8269; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8271; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8272; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8273; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8274; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8275; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8276; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8277; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8278; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8279; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8280; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8281; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8282; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd7;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8283; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8284; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8285; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8286; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8287; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8288; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8289; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8290; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8291; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8292; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8293; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8294; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8295; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8296; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8297; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd8298; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8299; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8300; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8301; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd8302; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8303; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8304; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8305; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8306; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8307; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8308; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd8309; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8310; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8311; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8312; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8313; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8314; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8315; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8316; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8317; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8318; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8319; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8320; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8321; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8322; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8323; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8324; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8325; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8326; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8328; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8329; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8330; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8331; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8332; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8333; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8334; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8335; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8336; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd8337; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8338; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8339; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8340; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8341; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8342; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8343; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8344; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8345; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8346; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8347; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8348; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8349; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8350; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8351; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8352; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8353; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8354; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8355; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8356; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8357; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8358; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8359; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8360; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd8361; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8362; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8363; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8364; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd8365; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd8366; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd14;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8367; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8368; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8369; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8370; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8371; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8372; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8373; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8374; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8375; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8376; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8377; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8378; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8379; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8381; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8383; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd8384; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8385; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8386; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8387; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd8388; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8389; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8390; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8391; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8392; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd8393; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd8394; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8395; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8396; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8397; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8398; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8399; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8401; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8402; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8403; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8404; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8405; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8406; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8407; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8411; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8412; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8413; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8414; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd8415; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd7;
#10 addr = 20'd8416; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd8417; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8418; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8419; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8420; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8421; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd8422; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd7;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8423; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8424; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8425; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8426; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8427; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8428; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8429; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8430; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8431; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8432; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8433; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8434; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8435; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8436; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8438; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd8440; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8441; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8442; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8443; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd4;
#10 addr = 20'd8444; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8445; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8446; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8447; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8448; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd8449; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd8450; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8451; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd8452; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8453; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8454; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8455; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8456; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8457; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8458; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8459; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8460; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8461; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8462; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8463; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8464; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8465; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8466; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8467; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8468; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8469; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8470; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8471; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd3;
#10 addr = 20'd8472; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8473; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8474; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8475; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8476; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8477; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd8478; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8479; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd8480; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8481; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8482; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8483; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8484; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8485; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8486; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8487; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8488; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8489; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8490; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8491; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8492; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8493; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8495; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8496; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8497; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd8498; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd8499; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd8500; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8501; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8502; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8503; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8504; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8505; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd9;
#10 addr = 20'd8506; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8507; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd8508; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8509; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8510; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8511; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8512; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8513; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8514; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8515; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8516; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8517; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8518; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8519; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8520; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8521; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd8522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8524; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8525; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8526; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd8527; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd8528; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8529; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8530; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8531; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd8532; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8533; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd1;
#10 addr = 20'd8534; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8535; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd8536; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8537; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8538; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8539; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8540; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8541; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8542; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8543; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8544; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8545; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8546; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd7;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8547; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8548; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8549; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8551; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8552; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8553; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8554; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd8555; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8556; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8557; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8558; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8559; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8560; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8561; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8562; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8563; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd8564; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8565; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8566; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8567; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8568; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8569; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8570; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8571; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8572; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8573; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8574; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8575; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8576; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8577; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8579; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8580; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8581; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8582; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd8583; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd8584; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8585; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8586; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8587; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8588; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8589; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd5;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8590; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8591; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8592; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8593; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8594; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8595; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8596; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8597; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8598; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8599; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8600; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8601; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8602; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd8603; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8604; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8605; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8607; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8608; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8609; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd8610; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd8611; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8612; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8613; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8614; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd8615; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8616; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8617; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8618; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8619; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8620; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8621; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8622; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8623; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8624; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8625; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8626; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8627; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8628; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8629; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8630; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd8;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd8631; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd8632; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8633; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8635; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd8636; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd8637; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8638; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd8639; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8640; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8641; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8642; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd8643; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8644; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8645; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8646; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8647; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8648; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8649; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8650; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8651; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8652; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8653; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8654; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8655; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8656; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8657; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8658; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd8659; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8660; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8661; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8663; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8664; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd8665; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd8666; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd8667; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8668; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8669; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8670; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd8671; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8672; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd8673; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd6;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8674; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8675; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8676; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8677; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8678; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8679; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8680; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8682; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8684; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8685; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8686; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8687; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8688; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8689; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8690; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8691; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8692; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd8693; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd8694; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd8695; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8696; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8697; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8698; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8699; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd8700; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd8701; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8702; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8703; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8704; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8705; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8706; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8707; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8708; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8709; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8710; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8712; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8713; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8714; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd8;data_in[31:28] = 4'd13;
#10 addr = 20'd8715; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd8716; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8717; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8718; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8719; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8720; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8721; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8722; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd8723; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8724; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8725; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8726; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd8727; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8728; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd8729; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8730; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8731; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8732; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8733; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8734; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8735; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8736; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8737; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8738; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8739; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8740; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8741; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8742; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd11;
#10 addr = 20'd8743; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd8744; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8746; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8747; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd8748; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8749; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd8750; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd0;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8751; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd8752; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8753; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8754; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8755; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd8756; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd8757; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8758; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8759; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd8760; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8761; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8762; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8763; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8764; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8765; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8766; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8767; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8768; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8769; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8770; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd8771; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd8772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8773; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8774; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8775; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8776; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd8777; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd0;
#10 addr = 20'd8778; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd8779; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8780; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8781; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8782; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8783; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8784; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8785; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8786; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8787; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8788; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8789; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8790; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8791; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8792; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8793; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8794; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8795; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8796; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8797; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8798; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8799; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd8800; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8801; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8802; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8803; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd3;
#10 addr = 20'd8804; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8805; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd8806; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd8807; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8808; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8809; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8810; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8811; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8812; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8813; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8814; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8815; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd8816; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8817; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8818; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8819; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8820; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8822; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8823; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8824; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8825; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8826; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8827; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd8828; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8829; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8830; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd8831; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8832; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8833; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd8834; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8835; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8836; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8837; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8838; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd8839; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd8840; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8841; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8842; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8843; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd8844; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8845; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8846; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8847; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8848; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8849; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8850; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8851; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8852; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8853; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8854; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8855; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd8856; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8857; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd8858; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd8859; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8860; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8861; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8862; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8863; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8864; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8865; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8866; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8867; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8868; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd8869; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8870; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8871; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8872; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8873; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8874; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8875; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8876; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8877; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8878; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8879; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8880; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8881; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8882; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8883; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd8884; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8885; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8887; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8888; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8889; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8890; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8891; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8892; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8893; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8894; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8895; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8896; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8897; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8898; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8899; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8900; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8901; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd8902; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8903; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8904; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8905; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8906; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8907; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8908; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8909; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8910; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8911; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd8912; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8914; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8915; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8916; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8917; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd8918; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8919; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd8920; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8921; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8922; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8923; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8924; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd8925; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8926; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8927; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8928; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8929; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8930; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8931; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8932; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8933; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8934; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8935; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8936; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8937; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8938; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8939; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8940; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd8941; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8942; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8943; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8944; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8945; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd8946; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8947; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8948; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8949; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8950; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8951; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8952; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8953; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8954; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd8955; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8956; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8957; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8958; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8959; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8960; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8961; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8962; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8963; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8964; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8965; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8966; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd8967; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd8968; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd8969; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd8970; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8971; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd8972; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8973; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd8974; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8975; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd8976; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd8977; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd8978; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd8979; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8980; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8981; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd8982; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd8983; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8984; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8985; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8986; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8987; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd8988; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8989; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd8990; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd8991; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd8992; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8993; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8994; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd8995; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd8996; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd8997; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd8998; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd8999; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9000; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9001; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd9002; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9003; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9004; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9005; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd9006; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9007; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9008; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9009; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9010; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9011; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9012; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9013; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9014; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9015; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9016; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9017; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9018; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9019; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9020; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9021; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9022; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9023; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9024; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9025; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9026; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9027; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9028; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9029; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9030; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd9031; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd9032; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9033; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9034; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9035; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9036; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9037; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9038; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd9039; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9040; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9041; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9042; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9043; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9044; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9045; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9046; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9047; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9048; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9049; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9050; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9051; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd14;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9052; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9053; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9054; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9055; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9056; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9057; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9058; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd9059; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9060; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9061; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9062; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9063; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd9064; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9065; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9066; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd9067; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9068; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9069; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9070; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9071; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9072; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9073; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9074; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9075; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9076; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9077; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9078; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9079; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9080; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9081; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9082; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9083; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9084; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9085; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9086; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9087; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9088; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9089; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9090; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9091; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd9092; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9093; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9094; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9095; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9096; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9097; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9098; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9099; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9100; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9101; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9102; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9103; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9104; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9105; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9106; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9107; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9108; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9109; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9110; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9111; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9112; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd4;
#10 addr = 20'd9113; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9114; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd9115; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9116; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9117; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9118; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd9119; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd9120; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9121; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9122; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9123; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd9124; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9125; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9126; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9127; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9128; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9129; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9130; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9131; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9132; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9133; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9135; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9137; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9138; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9139; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9140; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd8;
#10 addr = 20'd9141; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9142; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd9143; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9144; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9145; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9146; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd9147; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd9148; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9149; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9150; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9151; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9152; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9153; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9154; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9155; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9156; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9157; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9158; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9159; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9160; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9161; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9162; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9163; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9164; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9165; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9166; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9167; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9168; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9169; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9170; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd9171; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9172; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9173; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9174; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9175; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd8;
#10 addr = 20'd9176; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9177; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9178; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9179; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9180; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9181; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9182; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9183; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9184; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9185; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9186; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9187; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9188; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9189; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9190; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9191; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9192; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9193; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9194; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9195; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9196; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9197; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9198; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd9199; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9200; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9201; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9202; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd9203; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd9204; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9205; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9206; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9207; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9208; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9209; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9210; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9211; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9212; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9213; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9214; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9215; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9216; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9217; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9218; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9219; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9220; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9221; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9222; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9223; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9224; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd7;
#10 addr = 20'd9225; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9226; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9227; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9228; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9229; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9230; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd9231; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd9232; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9233; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9234; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9235; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9236; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9237; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9238; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9239; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9240; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9241; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9242; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9243; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9244; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9245; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9246; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9247; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9248; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd9249; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9250; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9251; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd3;
#10 addr = 20'd9252; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd9253; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9254; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9255; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9256; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9257; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9258; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd9259; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd9260; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9261; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9262; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9263; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9264; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9265; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9266; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9267; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9268; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9269; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9270; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9271; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9272; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9273; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9274; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd9275; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9276; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd9277; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9278; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9279; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd9280; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9281; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9282; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9283; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9284; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9285; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9286; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9287; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9288; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9289; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9290; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9291; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9292; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9293; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9294; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9295; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9296; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9297; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9298; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9299; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9300; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9301; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9302; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd9303; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd7;data_in[31:28] = 4'd11;
#10 addr = 20'd9304; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9305; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9306; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9307; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9308; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9309; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9310; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9311; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd9312; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9313; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9314; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd9315; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9316; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9317; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9318; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9319; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9320; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9321; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9322; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9323; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9324; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9325; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9326; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9327; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9328; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9329; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9330; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9331; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9333; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9334; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9335; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9336; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9337; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9338; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9339; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd9340; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9341; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9342; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9343; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9344; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9345; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9346; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9347; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9348; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9349; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9350; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9351; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9352; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9353; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9354; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9355; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9356; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9357; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9358; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9359; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9360; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9361; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9362; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9363; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9364; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9365; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd9366; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd9367; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9368; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9369; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9370; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9371; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9372; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9373; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9374; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9375; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9376; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9377; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9378; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9379; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9380; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9381; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9382; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9383; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9384; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9385; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9386; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9387; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9388; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9389; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd9390; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9391; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9392; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9393; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd9394; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd9395; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9396; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9397; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9398; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9399; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9400; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9401; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9402; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd9403; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9404; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9405; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9406; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9407; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9408; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9409; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9410; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9411; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9412; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9413; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9414; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9415; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9416; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd9417; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd3;
#10 addr = 20'd9418; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9419; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd3;
#10 addr = 20'd9420; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd9421; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9422; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9423; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9424; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9425; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd9426; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9427; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9428; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9429; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9430; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9431; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9432; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9433; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9434; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9435; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9436; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9437; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9438; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9439; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9440; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9441; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd9442; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9443; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9444; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9445; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9446; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd9447; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd8;
#10 addr = 20'd9448; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd9449; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9450; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9451; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9452; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9453; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9454; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9455; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9456; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9457; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9458; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9459; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9460; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9461; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9462; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9463; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9464; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9465; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9466; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9467; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9468; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9469; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd9470; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9471; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd9472; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9473; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9474; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9475; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9476; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd9477; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9478; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd9479; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9480; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd9481; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9482; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9483; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9484; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9485; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9486; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9487; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9488; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9489; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9490; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9491; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9492; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9493; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9494; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9495; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9496; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9497; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd6;data_in[31:28] = 4'd12;
#10 addr = 20'd9498; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd9499; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd6;
#10 addr = 20'd9500; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9501; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9502; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9503; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd9504; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd9505; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9506; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd10;
#10 addr = 20'd9507; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9508; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd9509; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd9;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9510; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9511; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9512; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9513; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9514; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9515; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9516; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9517; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9518; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9519; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9520; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9521; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9522; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9523; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9524; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9525; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd9526; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9527; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9528; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9529; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9530; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9531; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9532; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd9533; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9534; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd10;
#10 addr = 20'd9535; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9536; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9537; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9538; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9539; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9540; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9541; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9542; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9543; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9544; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9545; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9546; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9547; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9548; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9549; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9550; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9551; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9552; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9553; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd9;
#10 addr = 20'd9554; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9555; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9556; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9557; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9558; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9559; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd9560; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9561; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9562; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd12;
#10 addr = 20'd9563; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9564; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd9565; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9566; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9567; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9568; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9569; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9570; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9571; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9572; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9573; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9574; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9575; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9576; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9577; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9578; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9579; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9580; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9581; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd7;
#10 addr = 20'd9582; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9583; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9584; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9585; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9586; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9587; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd9588; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd9589; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9590; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd9591; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9592; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd9593; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd9594; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9595; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9596; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9597; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9598; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9599; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9600; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9601; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9602; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9603; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9604; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9605; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9606; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9607; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9608; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9609; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd9610; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd15;data_in[19:16] = 4'd10;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9611; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9612; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9613; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9614; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9615; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9616; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9617; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9618; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9619; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9620; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd9621; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9622; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9623; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9624; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9625; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9626; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9627; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9629; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9630; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9631; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9632; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9633; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9634; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9635; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9636; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd9637; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9638; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9639; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9640; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9641; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9642; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9643; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd9644; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd9645; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9646; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9647; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9648; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd9649; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9650; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9651; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd9652; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9653; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd9654; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9655; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9656; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9657; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9658; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9659; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9661; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9662; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9663; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9664; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd9665; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9666; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd9667; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9668; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9669; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9670; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9671; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9672; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9673; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9674; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9675; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9676; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd9677; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9678; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9679; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd9680; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9681; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd9682; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9684; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9685; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9686; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9687; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9688; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9689; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9690; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9691; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9692; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9693; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9694; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd9695; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9696; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9697; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9698; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9699; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd9700; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9701; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9702; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd9703; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9704; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd9705; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9706; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9707; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd9708; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9709; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd9710; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9711; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9712; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9713; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9714; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9715; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9716; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9717; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9718; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9719; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9720; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9721; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9722; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9723; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9724; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd9725; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9726; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9727; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9728; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9729; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9730; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9731; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9732; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd9733; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9734; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9735; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9736; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9737; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd9738; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9739; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9740; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9741; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9742; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9743; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9744; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9745; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9746; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9747; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9748; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9749; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9750; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9751; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9752; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9753; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9754; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd9755; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9756; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9757; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9758; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9759; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9760; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd9761; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9762; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd9763; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9764; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9765; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd9766; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9767; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9768; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9769; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9770; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9771; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9772; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9773; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9774; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9775; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd9776; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9777; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd9778; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd9779; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9780; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd2;
#10 addr = 20'd9781; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9782; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9783; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd9784; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9785; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9786; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9787; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9788; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd9789; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9790; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9791; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9792; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9793; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9795; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9796; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9797; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9798; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9799; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9800; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9801; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd9802; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9803; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9804; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd9805; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd9806; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9807; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9808; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9809; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9810; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd5;
#10 addr = 20'd9811; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd9812; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9813; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9814; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd9815; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9816; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd9817; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9818; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9819; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9820; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9821; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9822; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9823; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9824; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9825; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9826; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9827; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9828; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9829; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9830; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9831; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9832; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9833; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9834; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9835; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9836; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9837; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9838; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd8;
#10 addr = 20'd9839; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd5;
#10 addr = 20'd9840; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9841; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9842; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9843; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd9844; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd9845; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9846; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd9847; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9848; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd9849; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9850; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9851; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9852; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9853; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9854; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9855; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9856; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9857; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9858; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd9859; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9860; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9861; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9862; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9863; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9864; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd1;
#10 addr = 20'd9865; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9866; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd9867; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd9868; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9869; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9870; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9871; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9872; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd9873; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9874; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9875; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9876; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9877; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9878; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9879; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9880; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9881; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd9882; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9883; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9884; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9885; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9886; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd9887; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9888; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9889; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9890; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9891; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9892; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9893; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9894; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9895; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9896; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9897; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9898; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9899; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9900; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd9901; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9902; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9903; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9904; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9905; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9906; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9907; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9908; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9909; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd9910; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9911; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9912; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9913; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd9914; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9915; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9916; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9917; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd9918; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd9919; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9920; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd9921; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9922; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd9923; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9924; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9925; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd9926; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9927; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9928; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd9929; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9930; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9931; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd9932; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9933; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9934; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9935; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9936; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9937; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd9938; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9939; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9940; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9941; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd9942; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9943; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9944; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9945; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9946; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd9947; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9948; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9949; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9950; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9951; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd6;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9952; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd9953; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9954; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9955; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9956; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd9957; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9958; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd9959; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9960; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9961; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd9962; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9963; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9964; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9965; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9966; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9967; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9968; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9969; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9970; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9971; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd9972; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd9973; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd9974; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd9975; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd9976; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd9977; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd1;
#10 addr = 20'd9978; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd9979; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd9980; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd9981; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9982; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9983; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd9984; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd9985; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd9986; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd9987; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd9988; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd9989; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9990; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd9991; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9993; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9994; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd9995; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd9996; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd9997; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd9998; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd9999; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10000; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10001; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10002; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10003; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10004; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10005; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd10006; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd10007; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10008; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10009; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10010; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10011; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10012; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10013; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10014; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10015; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10016; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10017; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10018; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10019; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10020; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10021; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10022; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd10023; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10024; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10025; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10026; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10027; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10028; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10029; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd10030; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10031; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10032; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10033; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10034; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd10035; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10036; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10037; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10038; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd10039; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10040; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10042; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10043; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10044; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10045; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10046; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10047; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10048; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10049; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10050; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10051; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10052; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10053; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10054; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10055; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10056; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd10057; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10058; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10059; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10060; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10062; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd10063; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10064; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10065; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10066; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10067; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10068; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10069; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10070; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10071; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10072; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10073; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10074; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10075; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10076; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10077; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10078; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10079; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10080; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10081; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10082; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10083; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10084; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10085; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10086; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd10087; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10088; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd10089; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10090; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd10091; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10092; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10093; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10094; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10095; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10096; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10097; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10098; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10099; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10100; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10101; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10102; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10103; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10104; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10105; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10106; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10107; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10108; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10109; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10110; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10111; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10112; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10113; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd10114; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd10115; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10116; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd10117; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10118; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd10119; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10120; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10121; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10122; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10123; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10124; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10125; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10126; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10127; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10128; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10129; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10130; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10131; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10132; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10133; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10134; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10135; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10136; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10137; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10138; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10139; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10140; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd10141; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10142; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd10143; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10144; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd10145; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10146; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd10147; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10148; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10149; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10150; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10151; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10152; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10153; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10154; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10155; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10156; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10157; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10158; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10159; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10160; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10161; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10162; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10163; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10164; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10165; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10166; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10167; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd10168; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10169; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10170; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd10171; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10172; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10173; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd10174; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd10175; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10176; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10177; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10178; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10179; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10180; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd10181; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10182; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10183; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10184; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10185; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10186; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10187; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10189; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10190; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10191; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10192; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10193; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10194; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10195; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10196; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10197; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10198; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd8;
#10 addr = 20'd10199; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd1;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10200; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd10201; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd10202; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd2;
#10 addr = 20'd10203; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10204; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10205; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10206; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10207; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10208; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10209; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10210; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10211; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10212; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd10213; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10214; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10215; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10216; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10217; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10218; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10219; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10220; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10221; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10222; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10223; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10224; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10225; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd10226; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd10227; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10228; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd8;
#10 addr = 20'd10229; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd5;
#10 addr = 20'd10230; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10231; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10232; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10233; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10234; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10235; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10236; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10237; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10238; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10239; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10240; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd10241; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10242; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10243; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10244; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10245; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10246; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10247; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10248; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10249; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10250; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10251; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10252; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10253; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd6;
#10 addr = 20'd10254; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10255; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10256; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd10257; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd7;
#10 addr = 20'd10258; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10259; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10260; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10261; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10262; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10263; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10264; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10265; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10266; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10267; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10268; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd10269; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10270; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10271; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10272; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10273; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10274; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10275; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10276; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10277; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10278; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10279; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10280; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10281; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd10282; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10283; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10284; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10285; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10286; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd5;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10287; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10288; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10289; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10290; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10291; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10292; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10293; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10294; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10295; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10296; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd10297; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10298; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10299; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10300; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10301; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd10302; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10303; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10304; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10305; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10306; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10307; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10308; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10309; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd2;
#10 addr = 20'd10310; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10311; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10312; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10313; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10314; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10315; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10316; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10318; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10319; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10320; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd10321; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10322; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10323; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10324; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd10325; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10326; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10327; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10328; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10329; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10330; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10331; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10332; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10333; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10334; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10335; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10336; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd10337; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd10338; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10339; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10340; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10341; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10342; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10343; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10344; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10346; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10347; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10348; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10349; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10350; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10351; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10352; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd10353; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10354; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10355; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10356; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd10357; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10358; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10359; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10360; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10361; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10362; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10363; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10364; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd10365; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10366; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10367; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10368; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd5;
#10 addr = 20'd10369; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10370; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd12;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10371; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10372; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10374; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10375; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10376; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10377; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10378; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10379; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10380; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10382; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10383; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10384; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd10385; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10386; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10387; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10388; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10389; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10390; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10391; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10392; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10393; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10394; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10395; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd10396; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd10397; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10398; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10399; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10402; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10403; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10404; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd10405; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10406; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10407; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10408; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10409; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10410; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10411; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10412; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd10413; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10414; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10415; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10416; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10417; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10418; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10419; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10420; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10421; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10422; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd10423; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd7;
#10 addr = 20'd10424; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd10425; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd8;
#10 addr = 20'd10426; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10427; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd10428; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10430; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10431; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10432; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10433; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10434; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10435; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10436; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10437; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10438; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10439; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10440; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd10441; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10442; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10443; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10444; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10445; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10446; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10447; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10448; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10449; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10450; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd10451; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10452; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd10453; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd10454; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10455; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10456; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10457; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10459; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10460; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd10461; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10462; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10463; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10464; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10465; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10466; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10467; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10468; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd10469; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10470; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10471; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10472; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10473; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10474; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10475; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10476; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10477; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10478; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10479; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd2;
#10 addr = 20'd10480; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10481; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd10482; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10483; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10484; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10485; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10486; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10487; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10488; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10489; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10490; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10491; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10492; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10493; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10494; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10495; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10496; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd10497; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10498; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10499; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10500; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10501; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10502; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10503; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10504; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10505; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10506; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10507; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10508; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd10509; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd10510; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10511; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10512; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10514; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10515; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10516; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10517; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10518; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10519; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10520; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10521; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10522; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10523; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10524; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd10525; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10526; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10527; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd10528; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10529; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10530; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10531; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd10532; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd10533; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10534; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10535; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10536; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd10537; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10538; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10539; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd10540; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10542; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10543; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10544; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd10545; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd2;
#10 addr = 20'd10546; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10547; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10548; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10549; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10550; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10551; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10552; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd10553; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10554; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10555; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10556; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10557; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10558; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10559; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd10560; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10561; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10562; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd10563; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10564; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd10565; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10566; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10567; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10568; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10569; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10570; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10571; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10572; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10573; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd10574; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10575; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10576; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10577; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10578; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10579; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10580; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10581; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10582; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10583; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10584; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10585; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10586; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10587; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10588; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd10589; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10590; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd10591; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10592; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd9;
#10 addr = 20'd10593; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10594; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10595; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10596; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10597; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10598; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd10599; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10600; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10601; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10602; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10603; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10604; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10605; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10606; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10607; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10608; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10609; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10610; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10611; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10612; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10613; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10614; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10615; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd2;
#10 addr = 20'd10616; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10617; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10618; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10619; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd10620; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd4;
#10 addr = 20'd10621; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10622; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10623; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10624; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10625; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10626; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10627; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd10629; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10630; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10631; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10632; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10633; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10634; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10636; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10637; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10638; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10639; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10640; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10641; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10642; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10643; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10644; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10645; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10646; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10647; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10648; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd12;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10649; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd4;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10650; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10651; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10652; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10653; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10654; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10655; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10656; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd10657; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10658; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10659; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10660; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10661; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10662; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10663; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10664; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10665; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10666; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10667; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10668; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10669; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10670; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10671; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10672; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10673; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10674; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd10675; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd10676; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd10677; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10678; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10679; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10680; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10682; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10683; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10684; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10685; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10686; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10687; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10688; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10689; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10690; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10691; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10692; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10693; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10694; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10695; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10696; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10697; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10698; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10699; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10700; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd4;
#10 addr = 20'd10701; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10702; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd10703; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10704; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd12;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd10705; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10706; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10707; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10708; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10709; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10710; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10711; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10712; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10713; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10714; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10715; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10716; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10717; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10718; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10719; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10720; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10721; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10722; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10723; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10724; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10725; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10726; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10727; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10728; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd5;
#10 addr = 20'd10729; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10730; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd10731; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10732; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd10733; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10734; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10735; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd10736; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10737; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10738; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd10739; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10740; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10741; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10742; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10743; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10744; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10745; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10746; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10747; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10748; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10749; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10750; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10751; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10752; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10753; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10754; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd10755; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd10756; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd10757; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10758; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10759; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd10760; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd10761; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10762; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10763; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10764; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10765; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10767; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10768; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10769; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10770; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10771; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10772; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10773; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10774; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10775; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10776; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10777; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10778; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10779; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10780; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10781; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10782; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10783; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd10784; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd10785; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10786; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd10787; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd10788; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd3;
#10 addr = 20'd10789; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10790; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10791; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10792; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10793; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10795; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10796; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10797; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10798; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10799; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10800; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10801; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10802; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10803; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10804; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10805; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10806; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10807; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10808; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10809; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10810; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd10811; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10812; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10813; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10814; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10815; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10816; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd10817; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10818; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10819; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10820; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10821; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10822; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10823; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10824; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10825; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10826; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10827; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10828; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10829; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10830; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10831; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10832; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd10833; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd10834; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10835; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10836; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10837; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10838; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10839; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10840; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd10841; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10842; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10843; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd10844; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd10845; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10846; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10847; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10848; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10849; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10850; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10851; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd10852; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10853; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10854; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10855; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10856; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10857; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10858; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10859; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10860; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd10861; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10862; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10863; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10864; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10865; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10866; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10867; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10868; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10869; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10870; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10871; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10872; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10873; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10874; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10875; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10876; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10877; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10878; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10879; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd10880; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10881; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10882; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10883; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10884; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10885; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10886; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10887; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10888; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd10889; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10890; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10891; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10892; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10893; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10894; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10895; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10896; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10897; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10898; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd10899; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd10900; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10901; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10902; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10903; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10904; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd10905; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10906; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10907; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10908; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10909; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10910; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10911; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10912; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10913; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10914; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10915; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10917; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10918; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10919; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd10920; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10921; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10922; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10923; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10924; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd10925; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10926; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd5;
#10 addr = 20'd10927; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10928; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10929; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10930; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10931; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10932; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10933; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd10934; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10935; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd10936; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10937; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10938; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10939; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10940; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10941; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10942; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10943; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10944; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10945; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10946; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10947; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd10948; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10949; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd10950; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10951; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10952; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd10953; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10954; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10955; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10956; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10957; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10958; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd10959; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10960; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10961; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10962; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd10963; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10964; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd10965; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10966; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10967; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd10968; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10969; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10970; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10971; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10972; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd10973; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd10974; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd10975; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd10976; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10977; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd10978; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd10979; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd10980; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10981; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10982; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd10983; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd10984; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10985; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd10986; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10987; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10988; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10989; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd10990; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd10991; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd10993; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd10994; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd10995; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd10996; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10997; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd10998; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd10999; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11000; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11001; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11002; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd11003; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11004; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11005; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11006; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11007; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd11008; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11009; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11010; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11011; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd11012; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11013; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11014; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11015; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11016; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11017; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11018; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11020; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd11021; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11022; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11023; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11024; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd11025; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11026; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11027; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11028; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11029; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11030; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd11031; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11032; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd11033; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11034; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11035; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd13;data_in[31:28] = 4'd6;
#10 addr = 20'd11036; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11037; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11038; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11039; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd11040; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd11041; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11042; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11043; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11044; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11045; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11046; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11047; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11048; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd11049; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11050; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11051; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11052; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd11053; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11054; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11055; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11056; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11057; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11058; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd11059; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11060; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11061; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11062; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11063; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd12;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd11064; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11065; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11066; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11067; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd11068; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd11069; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11070; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11071; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11072; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11073; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11074; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11076; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11077; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11078; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11079; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11080; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11081; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11082; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11083; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11084; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11085; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11086; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd11087; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11088; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11089; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11090; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11091; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11092; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11093; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11094; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd2;
#10 addr = 20'd11095; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11096; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11097; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11098; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11099; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11100; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11101; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11102; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11103; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11104; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11105; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11106; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11107; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11108; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11109; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11110; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11111; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11112; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11113; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11114; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11115; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11116; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11117; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11118; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11119; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11120; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11121; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11122; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11123; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11124; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd11125; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11126; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11127; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11128; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11129; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11130; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11131; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11132; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11133; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd11134; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11135; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11136; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11137; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11138; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11139; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11140; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11141; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11142; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11143; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11144; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11145; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11146; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11147; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd11148; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd11149; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11150; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11151; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11152; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd11153; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11154; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11155; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11156; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11157; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11158; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11159; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11160; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11161; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11162; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11163; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11164; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11165; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11166; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11167; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11168; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11169; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11170; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11171; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11172; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11173; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11174; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11175; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd11176; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11177; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd11178; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd11179; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11180; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd3;
#10 addr = 20'd11181; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11182; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11183; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11184; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11185; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11186; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11187; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11188; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11189; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd11190; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11191; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11192; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11193; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11194; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11195; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11196; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11197; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd11198; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11199; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11200; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11201; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11202; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11203; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd11204; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11205; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd11206; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11207; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11208; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd11209; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11210; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11211; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11212; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11213; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11214; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11215; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11216; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11217; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd11218; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd11219; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11220; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11221; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11222; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11223; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11224; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11225; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd11226; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11227; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11228; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11229; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11230; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11231; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11232; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd11233; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11234; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd11235; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11236; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd11237; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11238; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11239; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11240; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11241; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11242; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11243; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11244; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11245; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11246; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11247; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11248; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd11249; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11250; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11251; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11252; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11253; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd11254; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11255; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11256; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11257; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11258; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11259; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11260; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd11261; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11262; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd11263; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd11264; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11265; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11266; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11267; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11268; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11269; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11270; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11271; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11272; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11273; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd11274; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd3;
#10 addr = 20'd11275; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11276; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11277; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11278; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11279; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11280; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11281; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd11282; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11283; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11284; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11285; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11286; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11287; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11288; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11289; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11290; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11291; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11292; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd0;
#10 addr = 20'd11293; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd10;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11294; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11295; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11296; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11297; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11298; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11299; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11300; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11301; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11302; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd11303; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11304; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11305; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11306; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11307; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11308; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11309; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd11310; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11311; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11312; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd11313; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11314; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11315; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd11316; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11317; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11318; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11319; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11320; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd11321; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11322; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11323; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11324; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11325; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11327; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11328; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11329; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11330; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11331; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11332; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11333; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11334; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11335; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11337; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd2;
#10 addr = 20'd11338; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11339; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11340; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11341; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11342; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11343; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd2;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd11344; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11345; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11346; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd11347; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd11348; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11349; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd9;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11350; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11351; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11352; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd11353; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11354; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11355; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11356; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11357; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11358; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11359; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11360; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11361; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11362; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11363; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11364; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11365; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd11366; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11367; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11368; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11369; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11370; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11371; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11372; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11373; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd11374; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd11375; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd11376; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11377; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd9;data_in[19:16] = 4'd1;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd0;
#10 addr = 20'd11378; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11379; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11380; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd11381; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11382; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11383; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11384; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11385; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11386; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11387; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd6;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11388; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11389; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11390; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11391; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11392; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11393; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11394; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11395; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11396; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11397; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11398; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11399; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11400; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11401; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd11402; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd11403; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11404; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd11405; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd0;
#10 addr = 20'd11406; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11407; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11408; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11409; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11411; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11412; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11413; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11414; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11415; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11416; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11417; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11418; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11419; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11420; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11421; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11422; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11423; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11424; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd11425; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11426; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11427; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd11428; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11429; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd1;
#10 addr = 20'd11430; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11431; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11432; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd11433; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd0;
#10 addr = 20'd11434; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11435; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11436; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11437; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11438; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11440; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11441; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11442; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11443; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd8;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11444; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11445; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11446; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11447; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11448; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11449; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11450; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11451; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11452; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd11453; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11454; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11455; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11456; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11457; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd1;
#10 addr = 20'd11458; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11459; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11460; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11461; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd0;
#10 addr = 20'd11462; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11463; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11464; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11465; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11466; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11468; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11469; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11470; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11471; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11472; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11473; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11474; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11475; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11476; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11477; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11478; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11479; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11480; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11481; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11482; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11483; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11484; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11485; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd0;
#10 addr = 20'd11486; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd11487; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11488; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11489; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd7;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd0;
#10 addr = 20'd11490; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11491; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11492; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11493; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11495; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11496; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11497; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11498; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11499; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd8;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11500; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11501; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11502; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11503; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd11504; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11505; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11506; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11507; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11508; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11509; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11510; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11511; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd11512; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11513; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd0;
#10 addr = 20'd11514; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11515; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11516; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11517; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd6;data_in[23:20] = 4'd12;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd11518; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11519; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11520; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11521; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11524; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11525; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11526; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11527; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd11528; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11529; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11530; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11531; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11532; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11533; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11534; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11535; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11536; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11537; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11538; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11539; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11540; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11541; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd11542; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11543; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11544; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd11545; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd6;data_in[23:20] = 4'd11;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd11546; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11547; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11548; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11549; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11551; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11552; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11553; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11554; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11555; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd6;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd11556; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11557; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11558; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd11559; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd11560; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11561; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11562; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11563; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11564; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11565; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11566; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11567; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11568; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11569; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11570; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11571; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11572; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd11573; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11574; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11575; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11576; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11577; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11579; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11580; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11581; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11582; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11583; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11584; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd11585; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11586; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11587; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11588; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11589; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11590; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11591; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11592; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11593; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11594; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11595; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd11596; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11597; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11598; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11599; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd11600; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11601; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd11602; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11603; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11604; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11605; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11607; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11608; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11609; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11610; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11611; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd11612; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd11613; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11614; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11615; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11616; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11617; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11618; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11619; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11620; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11621; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11622; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11623; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11624; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11625; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11626; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11627; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd11628; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11629; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11630; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11631; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11632; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11633; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11635; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11636; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11637; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11638; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11639; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd7;data_in[31:28] = 4'd0;
#10 addr = 20'd11640; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11641; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11642; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11643; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd11644; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11645; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11646; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11647; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11648; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11649; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11650; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11651; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11652; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11653; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11654; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11655; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11656; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd11657; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11658; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11659; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11660; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11661; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11662; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11663; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11664; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11665; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11666; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11667; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd0;
#10 addr = 20'd11668; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd11669; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11670; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11671; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11672; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd11673; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11674; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11675; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11676; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11677; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11678; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11679; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11680; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11681; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11682; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11683; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11684; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd11685; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11686; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11687; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11688; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11689; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11690; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11691; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11692; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11693; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11694; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11695; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd2;
#10 addr = 20'd11696; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11697; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11698; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11699; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11700; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd11701; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11702; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11703; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11704; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11705; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11706; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11707; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11708; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11709; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11710; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11711; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd11712; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11713; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11714; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11715; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11716; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11717; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11718; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11719; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11720; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11721; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd11722; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11723; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd5;
#10 addr = 20'd11724; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11725; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11726; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11727; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd11728; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd11729; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11730; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11731; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11732; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11733; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11734; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11735; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11736; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11737; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11738; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11739; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd5;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11740; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11741; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11742; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11743; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11744; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11745; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11746; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11747; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11748; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11749; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11750; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11751; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd8;
#10 addr = 20'd11752; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11753; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11754; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11755; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11756; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd11757; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11758; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11759; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11760; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11761; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd2;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11762; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11763; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11764; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11765; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11766; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11767; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd11768; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd11769; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11770; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11771; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11773; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11774; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11775; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11776; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11777; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11778; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11779; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd11780; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11781; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11782; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11783; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11784; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd11785; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11786; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11787; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11788; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11789; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11790; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11791; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11792; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11793; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11794; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11795; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11796; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11797; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11798; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11799; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11800; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11801; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11802; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11803; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11804; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11805; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11806; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11807; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11808; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11809; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11810; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11811; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd11812; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd11813; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11814; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11815; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11816; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11817; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11818; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11819; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11820; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11821; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11822; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11823; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd0;
#10 addr = 20'd11824; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd11825; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11826; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11827; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11828; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd11829; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11830; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11831; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd11832; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11833; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11834; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11835; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11836; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11837; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11838; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11839; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11840; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd11841; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11842; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11843; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11844; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11845; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11846; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11847; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd11848; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11849; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11850; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11851; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd11852; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11853; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11854; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11855; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11856; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd11857; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11858; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11859; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11860; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd11861; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11862; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11863; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd11864; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11865; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11866; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11867; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11868; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd11869; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11870; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11871; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11872; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd11873; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11874; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11875; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11876; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11877; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11878; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11879; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd11880; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd11881; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11882; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11883; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11884; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11885; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11886; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11887; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11888; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11889; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd11890; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11891; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11892; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11893; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11894; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11895; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11896; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd11897; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11898; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11899; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11900; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd11901; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11902; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11903; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11904; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11905; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11906; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11907; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd11908; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd0;
#10 addr = 20'd11909; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11910; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11911; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11912; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11914; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11915; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11916; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11917; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11918; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11919; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11920; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11921; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11922; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11923; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd11924; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd11925; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11926; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11927; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11928; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd11929; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11930; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11931; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11932; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11933; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11934; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11935; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd11936; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd11937; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11938; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd0;
#10 addr = 20'd11939; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11940; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd11941; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11942; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11943; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11944; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11945; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11946; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11947; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11948; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd11949; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11950; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11951; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd11952; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11953; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd11954; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11955; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11956; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11957; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11958; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11959; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11960; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11961; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11962; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11963; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd11964; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11965; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11966; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd11967; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd11968; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd11969; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11970; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11971; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11972; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd11973; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd11974; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd11975; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd11976; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11977; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11978; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd11979; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd11980; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11981; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd11982; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd11983; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd11984; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11985; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd6;
#10 addr = 20'd11986; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd11987; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd11988; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11989; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd11990; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11991; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd11992; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd11993; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd11994; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd11995; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11996; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd11997; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11998; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd11999; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12000; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12001; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12002; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12003; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12004; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12005; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12006; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12007; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd12008; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12009; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12010; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12011; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12012; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12013; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12014; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12015; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12016; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12017; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12018; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12019; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12020; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12021; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12022; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd12023; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12024; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12025; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12026; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12027; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12028; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12029; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12030; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12031; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12032; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd8;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12033; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12034; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12035; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd12036; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12037; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12038; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12039; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12040; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12042; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12043; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12044; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd12045; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12046; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12047; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd12048; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12049; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12050; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12051; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12052; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12053; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12054; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12055; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12056; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12057; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12058; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12059; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12060; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12061; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12062; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12063; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12064; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12065; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12066; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12067; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12068; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12069; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12070; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12071; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12072; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12073; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12074; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12075; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd12076; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12077; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12078; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12079; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12080; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12081; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12082; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12083; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12084; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12085; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12086; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12087; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12088; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12089; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12090; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd12091; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd12092; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12093; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12094; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12095; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12096; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12097; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12098; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12099; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12100; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12101; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12102; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12103; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12104; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12105; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12106; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12107; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd12108; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12109; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12110; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12111; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12112; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12113; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12114; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12115; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12116; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd8;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12117; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12118; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd0;data_in[31:28] = 4'd5;
#10 addr = 20'd12119; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12120; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12121; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12122; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12123; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12124; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12125; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12126; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12127; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12128; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12129; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12130; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12131; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12132; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12133; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12134; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12135; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd0;
#10 addr = 20'd12136; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12137; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12138; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12139; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12140; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12141; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd12142; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12143; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12144; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd9;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12145; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12146; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd5;
#10 addr = 20'd12147; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12148; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12149; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12150; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12151; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12152; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12153; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12154; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12155; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12156; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12157; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12158; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12159; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12160; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12161; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12162; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12163; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12164; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12165; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12166; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12167; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12168; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12169; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12170; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12171; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12172; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12173; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12174; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd12175; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd12176; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12177; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12178; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12179; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12180; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12181; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12182; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12183; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12184; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12185; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12186; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12187; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12188; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12189; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12190; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12191; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd1;data_in[27:24] = 4'd0;data_in[31:28] = 4'd2;
#10 addr = 20'd12192; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12193; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12194; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12195; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12196; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12197; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12198; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12199; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12200; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12201; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12202; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12203; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd12204; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12205; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12206; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12207; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12208; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd12209; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12210; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12211; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd12212; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12213; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd12214; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12215; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12216; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12217; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd0;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12218; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12219; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12220; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12221; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12222; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12223; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12224; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12225; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12226; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12227; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12228; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12229; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12230; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd12231; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd12232; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12233; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd12234; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12235; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12236; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd12237; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12238; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12239; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12240; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12241; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12242; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd12243; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd4;data_in[31:28] = 4'd2;
#10 addr = 20'd12244; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12245; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12246; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12247; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12249; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12250; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12251; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12252; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12253; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12254; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12255; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12256; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12257; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12258; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12259; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd12260; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12261; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12262; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12263; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12264; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd12265; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12266; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12267; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12268; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12269; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12270; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd1;
#10 addr = 20'd12271; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd4;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12272; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd1;
#10 addr = 20'd12273; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12274; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12275; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12277; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12278; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12279; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12280; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12281; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12282; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12283; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12284; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12285; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12286; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12287; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12288; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12289; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12290; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12291; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12292; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd12293; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12294; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12295; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12296; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12297; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12298; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd0;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd12299; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd12300; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd12301; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12302; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12303; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12304; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12305; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12306; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12307; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12308; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12309; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12310; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12311; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12312; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd7;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12313; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12314; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12315; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12316; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12317; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12318; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12319; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12320; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd12321; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12322; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12323; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12324; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12325; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd4;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12326; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd12327; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12328; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12329; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12330; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12331; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12333; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12334; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12335; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12337; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12338; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12339; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12340; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12341; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12342; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12343; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12344; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12346; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12347; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12348; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd12349; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12350; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12351; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12352; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12353; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd12354; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd12355; we = 1; data_in[3:0] = 4'd0;data_in[7:4] = 4'd0;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12356; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd3;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12357; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12358; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12359; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12360; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12361; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12362; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12363; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12364; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12365; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12366; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12367; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12368; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12369; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12370; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12371; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12372; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12373; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12374; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12375; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12376; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd12377; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12378; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12379; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12380; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12381; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd4;
#10 addr = 20'd12382; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd12383; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd0;data_in[11:8] = 4'd2;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd0;data_in[31:28] = 4'd1;
#10 addr = 20'd12384; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd12385; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12386; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12387; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12389; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12390; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd12391; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12392; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12393; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12394; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12395; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12396; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd5;data_in[31:28] = 4'd2;
#10 addr = 20'd12397; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12398; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12399; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12401; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12402; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12403; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12404; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd12405; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12406; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12407; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12408; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12409; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd5;
#10 addr = 20'd12410; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd7;
#10 addr = 20'd12411; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12412; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd0;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd2;
#10 addr = 20'd12413; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12414; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12415; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12416; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12417; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12418; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12419; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12420; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12421; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12422; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12423; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12424; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd7;data_in[31:28] = 4'd2;
#10 addr = 20'd12425; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12426; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12427; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12428; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12429; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12430; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12431; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12432; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd12433; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12434; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12435; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12436; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12437; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd0;data_in[27:24] = 4'd1;data_in[31:28] = 4'd6;
#10 addr = 20'd12438; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd12439; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd1;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12440; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12441; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd2;data_in[11:8] = 4'd0;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12442; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12443; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12444; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12445; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12446; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12447; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12448; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12449; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd12450; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12451; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12452; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd2;
#10 addr = 20'd12453; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12454; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12455; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12456; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd3;
#10 addr = 20'd12457; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd2;
#10 addr = 20'd12459; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12460; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd12461; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12462; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12463; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12464; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12465; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd2;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd6;
#10 addr = 20'd12466; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12467; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd0;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12468; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd2;data_in[15:12] = 4'd3;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12469; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd0;data_in[19:16] = 4'd0;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd2;
#10 addr = 20'd12470; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12471; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12472; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12473; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12474; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12475; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12476; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12477; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd12478; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12479; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12480; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd3;
#10 addr = 20'd12481; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12482; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12484; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12485; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12486; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd1;
#10 addr = 20'd12487; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12488; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd10;
#10 addr = 20'd12489; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12490; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12491; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12492; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12493; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd12494; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12495; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd2;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd2;data_in[31:28] = 4'd0;
#10 addr = 20'd12496; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd2;data_in[31:28] = 4'd4;
#10 addr = 20'd12497; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd2;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd2;data_in[31:28] = 4'd3;
#10 addr = 20'd12498; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12499; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12500; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12501; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12502; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12503; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12504; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12505; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12506; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12507; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12508; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd5;
#10 addr = 20'd12509; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12510; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12511; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd12512; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12513; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12514; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12515; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12516; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd1;data_in[15:12] = 4'd1;data_in[19:16] = 4'd1;data_in[23:20] = 4'd1;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd12517; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12518; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12519; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd0;
#10 addr = 20'd12520; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd2;data_in[31:28] = 4'd2;
#10 addr = 20'd12521; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd2;data_in[11:8] = 4'd3;data_in[15:12] = 4'd2;data_in[19:16] = 4'd2;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12522; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd2;data_in[11:8] = 4'd1;data_in[15:12] = 4'd2;data_in[19:16] = 4'd6;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd3;
#10 addr = 20'd12523; we = 1; data_in[3:0] = 4'd2;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd1;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12524; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd1;data_in[27:24] = 4'd1;data_in[31:28] = 4'd5;
#10 addr = 20'd12525; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd1;data_in[23:20] = 4'd2;data_in[27:24] = 4'd3;data_in[31:28] = 4'd3;
#10 addr = 20'd12526; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12527; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12528; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12529; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12530; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12531; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12532; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd12533; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd12534; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd12535; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12536; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd7;
#10 addr = 20'd12537; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd12538; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12539; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12540; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd3;data_in[27:24] = 4'd3;data_in[31:28] = 4'd4;
#10 addr = 20'd12541; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12542; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd3;data_in[19:16] = 4'd2;data_in[23:20] = 4'd2;data_in[27:24] = 4'd1;data_in[31:28] = 4'd1;
#10 addr = 20'd12543; we = 1; data_in[3:0] = 4'd1;data_in[7:4] = 4'd1;data_in[11:8] = 4'd2;data_in[15:12] = 4'd2;data_in[19:16] = 4'd3;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd12544; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12545; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12546; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12547; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12548; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12549; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12550; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12551; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12552; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12553; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12554; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12555; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12556; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12557; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12558; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12559; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12560; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd12561; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12562; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12563; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12564; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12565; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12566; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12567; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12568; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12569; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12570; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12571; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd12572; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12573; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12574; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12575; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12576; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12577; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12578; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12579; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12580; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12581; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12582; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12583; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12584; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12585; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12586; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12587; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12588; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12589; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12590; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12591; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd12592; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12593; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12594; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12595; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12596; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12597; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12598; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12599; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd12600; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12601; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12602; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12603; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12604; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd12605; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12606; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12607; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12608; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12609; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12610; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12611; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12612; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12613; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12614; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12615; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12616; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd12617; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12618; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12619; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12620; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12621; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12622; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12623; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12624; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12625; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12626; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12627; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd12628; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12629; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12630; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12631; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12632; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12633; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12634; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12635; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12636; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12637; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12638; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12639; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12640; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12641; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12642; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12643; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12644; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12645; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12646; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12647; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12648; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12649; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12650; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12651; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12652; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12653; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12654; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12655; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd12656; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12657; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12658; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12659; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12660; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12661; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12662; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12663; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12664; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12665; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12666; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12667; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12668; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12669; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12670; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12671; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12672; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12673; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12674; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12675; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12676; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12677; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12678; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12679; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12680; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12681; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12682; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12683; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12684; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12685; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12686; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12687; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12688; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12689; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12690; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12691; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12692; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12693; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12694; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12695; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12696; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12697; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12698; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12699; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12700; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd12701; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12702; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd12703; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12704; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12705; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12706; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12707; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12708; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12709; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12710; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12711; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12712; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12713; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12714; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12715; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12716; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12717; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12718; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12719; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12720; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12721; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12722; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12723; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12724; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12725; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12726; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12727; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12728; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12729; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12730; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12731; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12732; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12733; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12734; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12735; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12736; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd12737; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12738; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12739; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12740; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12741; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12742; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12743; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12744; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12745; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12746; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12747; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12748; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12749; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12750; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12751; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12752; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12753; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12754; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12755; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12756; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12757; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12758; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12759; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12760; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12761; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12762; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12763; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12764; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd12765; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12766; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12767; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12768; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12769; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12770; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12771; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12772; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12773; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12774; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12775; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12776; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12777; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12778; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12779; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12780; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12781; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12782; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12783; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12784; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12785; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12786; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12787; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12788; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12789; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12790; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12791; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12792; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12793; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12794; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd12795; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12796; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12797; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12798; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12799; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12800; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12801; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12802; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12803; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12804; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12805; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12806; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12807; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12808; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12809; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12810; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12811; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12812; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12813; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12814; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12815; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12816; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12817; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12818; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12819; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12820; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12821; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12822; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd12823; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd12824; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12825; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12826; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12827; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12828; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12829; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12830; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12831; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12832; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12833; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12834; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12835; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12836; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12837; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12838; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12839; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12840; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12841; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12842; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12843; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12844; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12845; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12846; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12847; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd12848; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12849; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12850; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd12851; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12852; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12853; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12854; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12855; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12856; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12857; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12858; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12859; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12860; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12861; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12862; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12863; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12864; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12865; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12866; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12867; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12868; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12869; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12870; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12871; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12872; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12873; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12874; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12875; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd12876; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12877; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12878; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12879; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12880; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12881; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12882; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12883; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12884; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12885; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12886; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12887; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12888; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12889; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12890; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12891; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12892; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12893; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12894; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12895; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12896; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12897; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12898; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12899; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12900; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12901; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12902; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd12903; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd12904; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12905; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12906; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12907; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12908; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12909; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12910; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12911; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12912; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12913; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12914; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12915; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12916; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12917; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12918; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12919; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12920; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12921; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12922; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12923; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12924; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12925; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12926; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12927; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12928; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12929; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12930; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd12931; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd12932; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12933; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12934; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12935; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12936; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12937; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12938; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12939; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12940; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12941; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12942; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12943; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12944; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12945; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12946; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12947; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12948; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12949; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12950; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12951; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12952; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12953; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12954; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12955; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12956; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12957; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12958; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd12959; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd12960; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd12961; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12962; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd12963; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12964; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12965; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12966; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12967; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12968; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd12969; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12970; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12971; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12972; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12973; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12974; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd12975; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12976; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12977; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12978; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12979; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12980; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12981; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12982; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12983; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd12984; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12985; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd12986; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd12987; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd12988; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12989; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12990; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12991; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd12992; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12993; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12994; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd12995; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd12996; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd12997; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd12998; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd12999; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13000; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13001; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13002; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13003; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13004; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13005; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13006; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13007; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13008; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13009; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13010; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13011; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13012; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13013; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13014; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13015; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13016; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13017; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd13018; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13019; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13020; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13021; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13022; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13023; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13024; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13025; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13026; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13027; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13028; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13029; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13030; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13031; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13032; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13033; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13034; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13035; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13036; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13037; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13038; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13039; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13040; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13041; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13042; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13043; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13044; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13045; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd13046; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13047; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13048; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13049; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13050; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13051; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13052; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13053; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13054; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13055; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13056; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13057; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13058; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13059; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13060; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13061; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13062; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13063; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13064; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13065; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13066; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13067; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13068; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13069; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13070; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13071; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13072; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13073; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd13074; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13075; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13076; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13077; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13078; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13079; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13080; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13081; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13082; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13083; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13084; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13085; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13086; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13087; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13088; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13089; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13090; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13091; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13092; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13093; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13094; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13095; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13096; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13097; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13098; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13099; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13100; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13101; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13102; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13103; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13104; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13105; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13106; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13107; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13108; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13109; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13110; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13111; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13112; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13113; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13114; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13115; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13116; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13117; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13118; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13119; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13120; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13121; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13122; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13123; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13124; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13125; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13126; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13127; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13128; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13129; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13130; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13131; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13132; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13133; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13134; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13135; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13136; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13137; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13138; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13139; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13140; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13141; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13142; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13143; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13144; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13145; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13146; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13147; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13148; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13149; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13150; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13151; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13152; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13153; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13154; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13155; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13156; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13157; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13158; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13159; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13160; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13161; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13162; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13163; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13164; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13165; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13166; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13167; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13168; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13169; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13170; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13171; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13172; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13173; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13174; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13175; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13176; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13177; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13178; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13179; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13180; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13181; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13182; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13183; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13184; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13185; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13186; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13187; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13188; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13189; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13190; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13191; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13192; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13193; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13194; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13195; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13196; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13197; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13198; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13199; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13200; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13201; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13202; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13203; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13204; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13205; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13206; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13207; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13208; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13209; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13210; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13211; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13212; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13213; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13214; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13215; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13216; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13217; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13218; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13219; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13220; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13221; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13222; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13223; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13224; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13225; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13226; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13227; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13228; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13229; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13230; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13231; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13232; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13233; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13234; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13235; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13236; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13237; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13238; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13239; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13240; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd13241; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13242; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13243; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13244; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13245; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13246; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13247; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13248; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13249; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13250; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13251; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13252; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13253; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13254; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13255; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13256; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13257; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13258; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13259; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13260; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13261; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13262; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13263; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13264; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13265; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13266; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13267; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13268; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd8;
#10 addr = 20'd13269; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13271; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13272; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13273; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13274; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13275; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13276; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13277; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13278; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13279; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13280; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd13281; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13282; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13283; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13284; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13285; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13286; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13287; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13288; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13289; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13290; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13291; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13292; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13293; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13294; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13295; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd13296; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd6;
#10 addr = 20'd13297; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13298; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13299; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13300; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13301; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13302; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13303; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13304; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13305; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13306; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13307; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13308; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13309; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13310; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13311; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13312; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13313; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13314; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13315; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13316; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13317; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13318; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13319; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13320; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13321; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13322; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13323; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd13324; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd13325; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13326; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13327; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13328; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13329; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13330; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13331; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13332; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13333; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13334; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13335; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13336; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13337; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13338; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13339; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13340; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13341; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13342; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13343; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13344; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13345; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13346; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13347; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13348; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13349; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13350; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13351; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13352; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd13353; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13354; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13355; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13356; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13357; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13358; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13359; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13360; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13361; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13362; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13363; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13364; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd13365; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13366; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13367; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13368; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13369; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13370; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13371; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13372; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13373; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13374; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13375; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13376; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13377; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13378; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13379; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13380; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd13381; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13383; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd13384; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13385; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13386; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13387; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13388; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13389; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13390; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13391; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13392; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13393; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13394; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13395; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13396; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13397; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13398; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13399; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13400; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13401; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13402; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13403; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13404; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13405; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13406; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13407; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13408; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd13409; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13410; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13411; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd13412; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13413; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13414; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13415; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13416; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13417; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13418; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13419; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13420; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13421; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13422; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13423; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13424; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13425; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13426; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13427; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd13428; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13429; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd13430; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13431; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13432; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13433; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13434; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13435; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13436; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13437; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13438; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd13440; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd13441; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13442; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13443; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13444; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13445; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13446; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13447; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13448; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13449; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13450; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13451; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13452; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13453; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13454; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13455; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd13456; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13457; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13458; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13459; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13460; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13461; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13462; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13463; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13464; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13465; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13466; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd13468; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd13469; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13470; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13471; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13472; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13473; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13474; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13475; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13476; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13477; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13478; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13479; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13480; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13481; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13482; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13483; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13484; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13485; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13486; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13487; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13488; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13489; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13490; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13491; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd13492; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13493; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13494; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13495; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd13496; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13497; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13498; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13499; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13500; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13501; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13502; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13503; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13504; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13505; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13506; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13507; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13508; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13509; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13510; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13511; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd13512; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13513; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13514; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13515; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13516; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13517; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13518; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13519; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13520; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13521; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd13524; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13525; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13526; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13527; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13528; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13529; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13530; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13531; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13532; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13533; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13534; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13535; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13536; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13537; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13538; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13539; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13540; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13541; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13542; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13543; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13544; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13545; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13546; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13547; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd13548; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13549; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13551; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13552; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13553; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13554; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13555; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13556; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13557; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13558; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13559; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13560; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13561; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13562; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13563; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13564; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13565; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13566; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13567; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13568; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13569; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13570; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13571; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13572; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13573; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13574; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13575; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd8;
#10 addr = 20'd13576; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13577; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd13579; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13580; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13581; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13582; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13583; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13584; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13585; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13586; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13587; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13588; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13589; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13590; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13591; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13592; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13593; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13594; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13595; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd13596; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13597; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13598; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13599; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13600; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13601; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13602; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13603; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd13604; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13605; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13606; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd13607; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13608; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13609; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13610; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13611; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13612; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13613; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13614; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13615; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13616; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13617; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13618; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13619; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13620; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13621; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13622; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13623; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13624; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13625; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13626; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13627; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13628; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13629; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13630; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13631; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd13632; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13633; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13634; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd13635; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13636; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13637; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13638; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13639; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13640; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13641; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13642; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13643; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13644; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13645; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13646; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13647; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13648; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13649; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13650; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13651; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13652; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd13653; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13654; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13655; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13656; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13657; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13658; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13659; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13660; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13661; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13662; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd13663; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13664; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13665; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13666; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13667; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13668; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13669; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13670; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13671; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13672; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13673; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13674; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13675; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13676; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13677; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13678; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13679; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13680; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd13681; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13682; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13683; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13684; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13685; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13686; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13687; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13688; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13689; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13690; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd13691; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13692; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13693; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13694; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13695; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13696; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13697; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13698; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13699; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13700; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13701; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13702; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13703; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13704; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13705; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13706; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13707; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13708; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd9;
#10 addr = 20'd13709; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13710; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13711; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13712; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd13713; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13714; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13715; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd13716; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13717; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13718; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd13719; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13720; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13721; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13722; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13723; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13724; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13725; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13726; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13727; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13728; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13729; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13730; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13731; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13732; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13733; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13734; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13735; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13736; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd13737; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13738; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13739; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13740; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd13741; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13742; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13743; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd13744; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13745; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13746; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13747; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13748; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13749; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13750; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13751; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13752; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13753; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13754; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13755; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13756; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13757; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13758; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13759; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13760; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd13761; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13762; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13763; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13764; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13765; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13766; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13767; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13768; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd13769; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13770; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13771; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13772; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13773; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13774; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13775; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13776; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13777; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13778; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13779; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13780; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13781; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13782; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13783; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13784; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13785; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13786; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13787; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13788; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13789; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13790; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13791; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13792; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13793; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13794; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13795; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13796; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd13797; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13798; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13799; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13800; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13801; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13802; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13803; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13804; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13805; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13806; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13807; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13808; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13809; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13810; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13811; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13812; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13813; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13814; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13815; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13816; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13817; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13818; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13819; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13820; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd13821; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13822; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13823; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13824; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd13825; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13826; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13827; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13828; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13829; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13830; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13831; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13832; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13833; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13834; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13835; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13836; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13837; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13838; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13839; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13840; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13841; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13842; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13843; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13844; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13845; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13846; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13847; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13848; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13849; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd13850; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13851; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13852; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13853; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13854; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13855; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13856; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13857; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13858; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13859; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13860; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd13861; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13862; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13863; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13864; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13865; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13866; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13867; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13868; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13869; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13870; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13871; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13872; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13873; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13874; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13875; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13876; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13877; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd13878; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13879; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13880; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13881; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13882; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd13883; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13884; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13885; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd13886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13887; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13888; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13889; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13890; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13891; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13892; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13893; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13894; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13895; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd15;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13896; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13897; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13898; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13899; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd13900; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13901; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13902; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13903; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13904; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13905; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd13906; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13907; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13908; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13909; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13910; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd7;
#10 addr = 20'd13911; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13912; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13913; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd13914; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13915; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13916; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13917; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13918; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13919; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13920; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13921; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13922; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13923; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13924; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13925; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13926; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13927; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13928; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13929; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13930; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13931; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13932; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13933; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd13934; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13935; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13936; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13937; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13938; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd13939; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13940; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13941; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd13942; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13943; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13944; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13945; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13946; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13947; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13948; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13949; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13950; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd13951; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13952; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd13953; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13954; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13955; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13956; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13957; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13958; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13959; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13960; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13961; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd6;
#10 addr = 20'd13962; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13963; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13964; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd13965; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13966; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd13967; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13968; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13969; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd13970; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd13971; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13972; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd13973; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13974; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13975; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd13976; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd13977; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13978; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd13979; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13980; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd13981; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd13982; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd13983; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13984; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd13985; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13986; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13987; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13988; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13989; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd8;
#10 addr = 20'd13990; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd13991; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd13992; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd13993; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd13;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd13994; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd13995; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd13996; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd13997; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd13998; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd13999; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14000; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14001; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14002; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14003; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14004; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14005; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14006; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd15;
#10 addr = 20'd14007; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14008; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14009; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14010; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14011; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14012; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14013; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14014; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14015; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14016; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14017; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd11;
#10 addr = 20'd14018; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14019; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14020; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd14021; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd14022; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd14023; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14024; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14025; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd14026; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14027; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14028; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14029; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14030; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14031; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14032; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14033; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14034; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd15;
#10 addr = 20'd14035; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14036; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14037; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14038; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14039; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14040; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14041; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14042; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14043; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14044; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14045; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14046; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14047; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14048; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd14049; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14050; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd4;
#10 addr = 20'd14051; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14052; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14053; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14054; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14055; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14056; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14057; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14058; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14059; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14060; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14061; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14062; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd14063; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14064; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14065; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14066; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14067; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14068; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14069; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14070; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14071; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14072; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14073; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd14074; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14075; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14076; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd3;data_in[23:20] = 4'd7;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd14077; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14078; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd5;
#10 addr = 20'd14079; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14080; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14081; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14082; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14083; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14084; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14085; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14086; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14087; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14088; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14089; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14090; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd14091; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14092; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14093; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14094; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14095; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14096; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14097; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14098; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14099; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14100; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14101; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14102; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14103; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14104; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd14105; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14106; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd7;
#10 addr = 20'd14107; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14108; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14109; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14110; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14111; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14112; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14113; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14114; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14115; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14116; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14117; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14118; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14119; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14120; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14121; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14122; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14123; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14124; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14125; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14126; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14127; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14128; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14129; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14130; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14131; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14132; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14133; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14134; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd6;
#10 addr = 20'd14135; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14137; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14138; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14139; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14140; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14141; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14142; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14143; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14144; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14145; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14146; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14147; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14148; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14149; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14150; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14151; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14152; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14153; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14154; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14155; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14156; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14157; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14158; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14159; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14160; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14161; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14162; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd6;
#10 addr = 20'd14163; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14164; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14165; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14166; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14167; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14168; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14169; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14170; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14171; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14172; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14173; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14174; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14175; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14176; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14177; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14178; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14179; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14180; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14181; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14182; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14183; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14184; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14185; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14186; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14187; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd14188; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14189; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14190; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd5;
#10 addr = 20'd14191; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14192; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14193; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14194; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14195; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14196; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14197; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14198; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14199; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14200; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14201; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14202; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14203; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14204; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14205; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14206; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14207; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14208; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14209; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14210; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14211; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14212; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14213; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14214; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14215; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14216; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14217; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14218; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd5;
#10 addr = 20'd14219; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14220; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14221; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14222; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14223; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14224; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14225; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14226; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14227; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14228; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14229; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14230; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14231; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14232; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14233; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14234; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14235; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14236; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14237; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14238; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14239; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14240; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14241; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14242; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14243; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14244; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14245; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14246; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd11;data_in[31:28] = 4'd4;
#10 addr = 20'd14247; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14249; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14250; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14251; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14252; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14253; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14254; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14255; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14256; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14257; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14258; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14259; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14260; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14261; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14262; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14263; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14264; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14265; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14266; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14267; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14268; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14269; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14270; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14271; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14272; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14273; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14274; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd14275; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14277; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14278; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14279; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14280; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14281; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14282; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14283; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14284; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14285; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14286; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14287; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14288; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14289; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14290; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14291; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14292; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14293; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14294; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14295; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14296; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14297; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14298; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14299; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14300; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14301; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14302; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd14303; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14304; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd14305; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14306; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14307; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14308; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14309; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14310; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14311; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14312; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14313; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14314; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14315; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14316; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14317; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14318; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14319; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14320; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14321; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14322; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14323; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14324; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14325; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14326; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd14327; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14328; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14329; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14330; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd14331; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd14333; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14334; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14335; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14336; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14337; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14338; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14339; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14340; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14341; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14342; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14343; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14344; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14345; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14346; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14347; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14348; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14349; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14350; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14351; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14352; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14353; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14354; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14355; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14356; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14357; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14358; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd14359; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14360; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd14361; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14362; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14363; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14364; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14365; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14366; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14367; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14368; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14369; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14370; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14371; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14372; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14373; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14374; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14375; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14376; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14377; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14378; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14379; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14380; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14381; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14382; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14383; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14384; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14385; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14386; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd11;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd14387; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd14389; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14390; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14391; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14392; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14393; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14394; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14395; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14396; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14397; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14398; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14399; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14400; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14401; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14402; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14403; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14404; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14405; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14406; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14407; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14408; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14409; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14410; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14411; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14412; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14413; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14414; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd9;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd14415; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14416; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14417; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14418; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14419; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14420; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14421; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14422; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14423; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14424; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14425; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14426; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14427; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14428; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14429; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14430; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14431; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14432; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14433; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14434; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14435; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14436; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14437; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14438; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14439; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14440; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14441; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd14442; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd14443; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14444; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14445; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14446; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14447; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14448; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14449; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14450; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14451; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14452; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14453; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14454; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14455; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14456; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd14457; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14458; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14459; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14460; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14461; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14462; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14463; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14464; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14465; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd14466; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14467; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14468; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14469; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14470; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14471; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14472; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14473; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14474; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14475; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14476; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14477; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14478; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14479; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14480; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14481; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14482; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14483; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14484; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14485; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14486; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14487; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14488; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14489; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14490; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14491; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14492; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14493; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14494; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14495; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14496; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14497; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd14498; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14499; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14500; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14501; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14502; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14503; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14504; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14505; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14506; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14507; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14508; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14509; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14510; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14511; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd14512; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd14513; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd14514; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14515; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14516; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14517; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14518; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14519; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14520; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14521; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14522; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14523; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14524; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14525; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14526; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14527; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14528; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14529; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14530; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14531; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14532; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14533; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14534; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14535; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14536; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14537; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14538; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14539; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd14540; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14541; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14542; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14543; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14544; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14545; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14546; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14547; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14548; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14549; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14550; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14551; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14552; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14553; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14554; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14555; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14556; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14557; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14558; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14559; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14560; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14561; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14562; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14563; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14564; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14565; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14566; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14567; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14568; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14569; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14570; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14571; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14572; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14573; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14574; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14575; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14576; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14577; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14578; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14579; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14580; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14581; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14582; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14583; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14584; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14585; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14586; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14587; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14588; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14589; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14590; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14591; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14592; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14593; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14594; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14595; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14596; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14597; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14598; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14599; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14600; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14601; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14602; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14603; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14604; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14605; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14606; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14607; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14608; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14609; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14610; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14611; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14612; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14613; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14614; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14615; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14616; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14617; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14618; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14619; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14620; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14621; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14622; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14623; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14624; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14625; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14626; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14627; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14628; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14629; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14630; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14631; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14632; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14633; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14634; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14635; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14636; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd12;
#10 addr = 20'd14637; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd14638; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd9;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14639; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14640; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14641; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14642; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14643; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14644; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14645; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14646; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14647; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14648; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14649; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14650; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14651; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14652; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14653; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14654; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14655; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd14656; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14657; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14658; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14659; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14660; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14661; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14662; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14663; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14664; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14665; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14666; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14667; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14668; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14669; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14670; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14671; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14672; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14673; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14674; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14675; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14676; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14677; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14678; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14679; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14680; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14681; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14682; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14683; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd14684; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd14685; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14686; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14687; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd14688; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14689; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14690; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14691; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14692; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14693; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd14694; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14695; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14696; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14697; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14698; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14699; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14700; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14701; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14702; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14703; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14704; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14705; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14706; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14707; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14708; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14709; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14710; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14711; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14712; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd14713; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14714; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd14715; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd14716; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14717; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14718; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14719; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14720; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14721; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14722; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14723; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd14724; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14725; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14726; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14727; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14728; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14729; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14730; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14731; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14732; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14733; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14734; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14735; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14736; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14737; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd14738; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14739; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14740; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd14741; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd14742; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd14743; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd14744; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14745; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14746; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14747; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14748; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd14749; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14750; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14751; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd14752; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14753; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14754; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14755; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14756; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14757; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14758; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14759; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14760; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd14761; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14762; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14763; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd14764; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14765; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14766; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14767; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14768; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd14769; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd14770; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd14771; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd12;
#10 addr = 20'd14772; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14773; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14774; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14775; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14776; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14777; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd12;
#10 addr = 20'd14778; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14779; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd14780; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14781; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14782; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14783; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14784; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14785; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14786; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14787; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14788; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14789; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14790; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14791; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14792; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14793; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14794; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14795; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd14796; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd14797; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14798; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14799; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14800; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14801; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14802; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14803; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd14804; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14805; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd14806; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14807; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd14808; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14809; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14810; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14811; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14812; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14813; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14814; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14815; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14816; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14817; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14818; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14819; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd14820; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14821; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14822; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14823; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14824; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14825; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14826; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd14827; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd3;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd14828; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14829; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14830; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14831; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14832; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14833; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd14834; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14835; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd14836; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14837; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14838; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14839; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14840; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14841; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14842; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14843; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14844; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14845; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14846; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14847; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14848; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14849; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14850; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14851; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14852; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14853; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd14854; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd14855; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14856; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14857; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14858; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14859; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd14860; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14861; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd14862; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14863; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd14864; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14865; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14866; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14867; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14868; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14869; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14870; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14871; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14872; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14873; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14874; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14875; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14876; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14877; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14878; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14879; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd14880; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14881; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd14882; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd3;
#10 addr = 20'd14883; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14884; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14885; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14886; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14887; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd14888; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14889; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14890; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14891; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14892; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14893; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14894; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14895; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14896; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14897; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14898; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14899; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14900; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14901; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14902; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14903; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14904; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14905; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14906; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14907; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd14908; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd14909; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd14910; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd14911; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14912; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14913; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14914; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd14915; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14916; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14917; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd14918; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd14919; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14920; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14921; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14922; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14923; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14924; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14925; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14926; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14927; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd14928; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14929; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14930; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14931; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14932; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14933; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14934; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14935; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd14936; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd14937; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd14938; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd14939; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd14940; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14941; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14942; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd14943; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14944; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14945; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14946; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14947; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd14948; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14949; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14950; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14951; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14952; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14953; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14954; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14955; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14956; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14957; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14958; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14959; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14960; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14961; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14962; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd14963; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd14964; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd14965; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14966; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd3;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd3;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd14967; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14968; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14969; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14970; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd14971; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd14972; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd14973; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14974; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14975; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14976; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14977; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14978; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14979; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14980; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14981; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd14982; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd14983; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd14984; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd14985; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd14986; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd14987; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd14988; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd14989; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd14990; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd14991; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd14992; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd14993; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd14994; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd3;data_in[19:16] = 4'd5;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd14995; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14996; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14997; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd14998; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd14999; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15000; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd10;
#10 addr = 20'd15001; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15002; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15003; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15004; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15005; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15006; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15007; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15008; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15009; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15010; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15011; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15012; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15013; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15014; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd15;
#10 addr = 20'd15015; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd15016; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15017; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15018; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15019; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15020; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15021; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15022; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15023; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15024; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15025; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15026; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd15027; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15028; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15029; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15030; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15031; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15032; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15033; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15034; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15035; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15036; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15037; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15038; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15039; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15040; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15042; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd15043; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd12;
#10 addr = 20'd15044; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15045; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15046; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15047; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15048; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15049; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd15050; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd15051; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15052; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15053; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15054; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd15055; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15056; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd12;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15057; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15058; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15059; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15060; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15061; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15062; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15063; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15064; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15065; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15066; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15067; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15068; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15069; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15070; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15071; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15072; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15073; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15074; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15075; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15076; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15077; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15078; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15079; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15080; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15081; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15082; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15083; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15084; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15085; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15086; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15087; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15088; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15089; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15090; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15091; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15092; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15093; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15094; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15095; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15096; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15097; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15098; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd15099; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15100; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15101; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15102; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd15103; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15104; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15105; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15106; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15107; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15108; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15109; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15110; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15111; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15112; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15113; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15114; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15115; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15116; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15117; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15118; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15119; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15120; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15121; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15122; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15123; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15124; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15125; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15126; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15127; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15128; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15129; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15130; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15131; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15132; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15133; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd15135; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15136; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15137; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15138; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15139; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15140; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15141; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15142; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15143; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15144; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15145; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15146; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15147; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15148; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15149; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15150; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15151; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15152; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15153; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15154; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15155; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15156; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15157; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15158; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15159; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15160; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15161; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15162; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15163; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15164; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15165; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15166; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd15167; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15168; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15169; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15170; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15171; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15172; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15173; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15174; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15175; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15176; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15177; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15178; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15179; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15180; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15181; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15182; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15183; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15184; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15185; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15186; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15187; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15188; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15189; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15190; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd15191; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15192; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15193; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15194; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd15195; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15196; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15197; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15198; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15199; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15200; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15201; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15202; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15203; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15204; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15205; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15206; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15207; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15208; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15209; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15210; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15211; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15212; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd15213; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15214; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15215; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15216; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15217; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15218; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15219; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15220; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15221; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15222; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd15223; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15224; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15225; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15226; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15227; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15228; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15229; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15230; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15231; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15232; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15233; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15234; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15235; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15236; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15237; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15238; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15239; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15240; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15241; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd15242; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15243; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15244; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd15245; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd15246; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15247; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15248; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15249; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15250; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd15251; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15252; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15253; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15254; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15255; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15256; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15257; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15258; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15259; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15260; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15261; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15262; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15263; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15264; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15265; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15266; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15267; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15268; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15269; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd15270; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15271; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15272; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd15273; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd15274; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15275; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15276; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15277; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15278; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd15279; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15280; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15281; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15282; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd15283; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15284; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15285; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15286; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15287; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15288; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15289; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15290; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15291; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15292; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15293; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15294; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15295; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15296; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15297; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15298; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15299; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15300; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd15301; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15302; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15303; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15304; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15305; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15306; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd15307; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15308; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15309; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15310; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd15311; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15312; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15313; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15314; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15315; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15316; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15317; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15318; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15319; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15320; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15321; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15322; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15323; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15324; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15325; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15326; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15327; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd15328; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd15329; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15330; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15331; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15332; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15333; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15334; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd15335; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15336; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15337; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15338; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd11;
#10 addr = 20'd15339; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15340; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15341; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15342; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15343; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15344; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15345; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15346; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15347; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15348; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15349; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15350; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15351; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15352; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15353; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15354; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15355; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd15356; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd15357; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15358; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15359; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15360; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15361; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15362; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15363; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd15364; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15365; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15366; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd15367; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15368; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15369; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15370; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15371; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15372; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15373; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15374; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15375; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15376; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15377; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15378; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15379; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15380; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15381; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd15382; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15383; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15384; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd15385; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15386; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15387; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15388; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15389; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15390; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15391; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd15392; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15393; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15394; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15395; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15396; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15397; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15398; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15399; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15400; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15401; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15402; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15403; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15404; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15405; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15406; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15407; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15408; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd15409; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15410; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15411; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15412; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd13;
#10 addr = 20'd15413; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15414; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15415; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15416; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15417; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15418; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15419; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd13;
#10 addr = 20'd15420; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15421; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15422; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15423; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15424; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15425; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15426; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15427; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15428; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15429; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15430; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15431; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15432; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15433; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15434; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15435; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15436; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd15437; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15438; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15439; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15440; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15441; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15442; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15443; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15444; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15445; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15446; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd15447; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd12;
#10 addr = 20'd15448; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15449; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15450; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15451; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15452; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15453; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15454; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15455; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15456; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15457; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15458; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15459; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15460; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15461; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15462; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15463; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15464; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd15465; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15466; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd15467; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15468; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15469; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15470; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15471; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15472; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15473; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15474; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15475; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd15476; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15477; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15478; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15479; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15480; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15481; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15482; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15483; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15484; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15485; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15486; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15487; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15488; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15489; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15490; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15491; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15492; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15493; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15494; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15495; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15496; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd15497; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15498; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15499; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15500; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15501; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15502; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd15503; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd15504; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15505; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15506; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15507; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15508; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15509; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15510; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15511; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15512; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15513; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15514; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15515; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15516; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15517; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15518; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15519; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15520; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15521; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15522; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15523; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd15524; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15525; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15526; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15527; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15528; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15529; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15530; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15531; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15532; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15533; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15534; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15535; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15536; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15537; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15538; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15539; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15540; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15541; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15542; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15543; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15544; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15545; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15546; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd15547; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15548; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd15549; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15550; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15551; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15552; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15553; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15554; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15555; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15556; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15557; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15558; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15559; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15560; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15561; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15562; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15563; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15564; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15565; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15566; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15567; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15568; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15569; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15570; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15571; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15572; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15573; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15574; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd15;
#10 addr = 20'd15575; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd15;
#10 addr = 20'd15576; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd15577; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15578; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15579; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15580; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15581; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15582; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15583; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd15584; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15585; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15586; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd15587; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15588; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15589; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15590; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15591; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15592; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15593; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15594; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15595; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15596; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15597; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15598; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15599; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15600; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15601; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15602; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15603; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15604; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15605; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15606; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15607; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15608; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15609; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15610; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15611; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd15612; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15613; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15614; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15615; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15616; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15617; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15618; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15619; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15620; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15621; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15622; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15623; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15624; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15625; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15626; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15627; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15628; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15629; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15630; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15631; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15632; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15633; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15634; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15635; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd15636; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15637; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd15638; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15639; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15640; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15641; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15642; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15643; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15644; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15645; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15646; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15647; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15648; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15649; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15650; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15651; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15652; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15653; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15654; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15655; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15656; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15657; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15658; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15659; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15660; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15661; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd15662; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15663; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd15664; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15665; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15666; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd15667; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15668; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15669; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd15670; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15671; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15672; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15673; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15674; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15675; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15676; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15677; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15678; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15679; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15680; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15681; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15682; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15683; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15684; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15685; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15686; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15687; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15688; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15689; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15690; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd15691; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd15692; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15693; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15694; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd15695; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15696; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15697; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15698; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15699; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15700; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15701; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15702; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15703; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15704; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15705; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15706; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15707; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15708; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15709; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15710; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15711; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15712; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15713; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd15714; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15715; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd15716; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15717; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15718; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd15719; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd12;
#10 addr = 20'd15720; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15721; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15722; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15723; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15724; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15725; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd15726; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15727; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15728; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15729; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15730; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15731; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15732; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15733; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15734; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15735; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15736; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15737; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15738; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15739; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15740; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15741; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd15742; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15743; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd15744; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15745; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15746; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15747; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd15748; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15749; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15750; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15751; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15752; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15753; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15754; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15755; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15756; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15757; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15758; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15759; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15760; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15761; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15762; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15763; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15764; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15765; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15766; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15767; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd15768; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd15769; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd15;
#10 addr = 20'd15770; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd10;
#10 addr = 20'd15771; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd15772; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15773; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15774; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd15775; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd15776; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15777; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15778; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd15779; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15780; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15781; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15782; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15783; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15784; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15785; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15786; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15787; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15788; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15789; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15790; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15791; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15792; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15793; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15794; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15795; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15796; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15797; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd15798; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15799; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15800; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15801; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15802; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd15803; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15804; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15805; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd15806; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd12;
#10 addr = 20'd15807; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd15808; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15809; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15810; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15811; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15812; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15813; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15814; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15815; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15816; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15817; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15818; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15819; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15820; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15821; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15822; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15823; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15824; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15825; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd13;
#10 addr = 20'd15826; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd15827; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15828; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15829; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15830; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15831; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd15832; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15833; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd15834; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd13;
#10 addr = 20'd15835; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15836; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15837; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15838; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15839; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd15840; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd14;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15841; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15842; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15843; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15844; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15845; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15846; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15847; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15848; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15849; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15850; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15851; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15852; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15853; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd15854; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd12;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15855; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15856; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd15857; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15858; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15859; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd15860; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd15861; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15862; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd15863; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15864; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15865; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd15866; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15867; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd15868; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15869; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15870; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15871; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15872; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15873; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15874; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15875; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15876; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15877; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15878; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd15879; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15880; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15881; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd15882; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15883; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd15884; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd15885; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd15886; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15887; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd15888; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15889; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15890; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15891; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd15892; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15893; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15894; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15895; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15896; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15897; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd15898; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15899; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15900; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15901; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15902; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15903; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15904; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15905; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15906; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15907; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15908; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15909; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15910; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd15;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15911; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd15912; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd15913; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15914; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15915; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd15916; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15917; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd15918; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15919; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15920; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15921; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15922; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd15923; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15924; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd15925; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd15926; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15927; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15928; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15929; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15930; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15931; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15932; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd15933; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15934; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15935; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15936; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15937; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15938; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd15939; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15940; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd15941; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15942; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15943; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15944; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15945; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15946; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15947; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15948; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15949; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15950; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15951; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15952; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15953; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd15954; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15955; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15956; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15957; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15958; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15959; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15960; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15961; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15962; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15963; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15964; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15965; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd15966; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd15967; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15968; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15969; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd15970; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd15971; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd6;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15972; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15973; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15974; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15975; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd15976; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd15977; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd15978; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd15979; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd15980; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd15981; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd15982; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15983; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15984; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd15985; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd15986; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd15987; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd15988; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd15989; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd15990; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd15991; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd15992; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd15993; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd15994; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd15995; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd15996; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd15997; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd15998; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd15999; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16000; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16001; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16002; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16003; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16004; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16005; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16006; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16007; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16008; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16009; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd16010; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16011; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16012; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16013; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16014; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16015; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16016; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16017; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16018; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16019; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16020; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16021; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16022; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16023; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16024; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16025; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16026; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd16027; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16028; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16029; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16030; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16031; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16032; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16033; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16034; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd16035; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16036; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16037; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd16038; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16039; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16040; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16041; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16042; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16043; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16044; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16045; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16046; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16047; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16048; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16049; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16050; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16051; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16052; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16053; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16054; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16055; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16056; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16057; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16058; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16059; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16060; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16061; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16062; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd16063; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16064; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16065; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16066; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16067; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16068; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16069; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16070; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16071; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16072; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16073; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16074; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16075; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16076; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16077; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd16078; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16079; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16080; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16081; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16082; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd16083; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16084; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16085; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16086; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16087; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16088; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16089; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16090; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16091; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16092; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16093; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd16094; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16095; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16096; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16097; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16098; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16099; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16100; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16101; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16102; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16103; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16104; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16105; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16106; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16107; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16108; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16109; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16110; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd12;
#10 addr = 20'd16111; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd8;
#10 addr = 20'd16112; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16113; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16114; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16115; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16116; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16117; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16118; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16119; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd16120; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16121; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd16122; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16123; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16124; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16125; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16126; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16127; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16128; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16129; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16130; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16131; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16132; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd16133; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16134; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16135; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd16137; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16138; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd16139; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd16140; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16141; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16142; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16143; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16144; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd16145; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16146; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16147; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16148; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16149; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16150; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16151; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16152; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16153; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd16154; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16155; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16156; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16157; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16158; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16159; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16160; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16161; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16162; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16163; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16164; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16165; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16166; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16167; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd16168; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16169; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16170; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16171; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16172; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16173; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16174; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16175; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16176; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16177; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16178; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16179; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16180; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16181; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16182; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16183; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16184; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16185; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16186; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16187; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16188; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16189; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16190; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd16191; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16192; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd16193; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16194; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16195; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd16196; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16197; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16198; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16199; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16200; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16201; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16202; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16203; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16204; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16205; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16206; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16207; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16208; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16209; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16210; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16211; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16212; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16213; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16214; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16215; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16216; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd16217; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd16218; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16219; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16220; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16221; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd16222; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16223; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16224; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16225; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16226; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16227; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16228; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16229; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16230; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd16231; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16232; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16233; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16234; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16235; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16236; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16237; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16238; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16239; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16240; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16241; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16242; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16243; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16244; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd16245; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd16246; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16247; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16249; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd14;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd16250; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16251; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16252; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16253; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16254; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16255; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16256; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16257; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16258; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd16259; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd16260; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16261; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16262; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16263; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16264; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16265; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16266; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16267; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16268; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16269; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16270; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16271; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16272; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16273; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16274; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd16275; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16277; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd16278; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd16279; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd7;data_in[19:16] = 4'd3;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16280; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16281; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16282; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16283; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16284; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16285; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16286; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd16287; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd16288; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16289; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16290; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16291; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16292; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16293; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16294; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16295; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16296; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16297; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16298; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16299; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16300; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd16301; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16302; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16303; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16304; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16305; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16306; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd14;
#10 addr = 20'd16307; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16308; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16309; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16310; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16311; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16312; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16313; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16314; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd16315; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd16316; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16317; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16318; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16319; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16320; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16321; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16322; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16323; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16324; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16325; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16326; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16327; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16328; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd16329; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16330; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16331; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16332; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16333; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd15;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16334; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd3;data_in[11:8] = 4'd4;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16335; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16336; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16337; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16338; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16339; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16340; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16341; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16342; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd16343; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd16344; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16346; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16347; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16348; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16349; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16350; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16351; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16352; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16353; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16354; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16355; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16356; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd16357; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16358; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16359; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16360; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd16361; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16362; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16363; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16364; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16365; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16366; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16367; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16368; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16369; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16370; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd16371; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16372; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16374; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16375; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16376; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16377; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16378; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16379; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16380; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16381; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16382; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16383; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16384; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd16385; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16386; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd16387; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16388; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd16389; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16390; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd16391; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16392; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16393; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16394; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16395; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16396; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16397; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16398; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd16399; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16400; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16402; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16403; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16404; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16405; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16406; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16407; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16408; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16409; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16410; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16411; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16412; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd16413; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16414; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd16415; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16416; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd16417; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd16418; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16419; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16420; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16421; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16422; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16423; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16424; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16425; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16426; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16427; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16428; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16429; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16430; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16431; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16432; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16433; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16434; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16435; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16436; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16437; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16438; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16439; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd16440; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd16441; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16442; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16443; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16444; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16445; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd16446; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16447; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16448; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16449; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16450; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16451; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16452; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd16453; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16454; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16455; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16456; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16457; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16458; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16459; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16460; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16461; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16462; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16463; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16464; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16465; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16466; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16467; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd16468; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd16469; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16470; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd16471; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16472; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16473; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd16474; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd8;
#10 addr = 20'd16475; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16476; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16477; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16478; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16479; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16480; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16481; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16482; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd16483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16484; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16485; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16486; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16487; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16488; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16489; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16490; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16491; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16492; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16493; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16494; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16495; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16496; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16497; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16498; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16499; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16500; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd16501; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd3;data_in[31:28] = 4'd9;
#10 addr = 20'd16502; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16503; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16504; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16505; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16506; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16507; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16508; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16509; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16510; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd16511; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16512; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd16513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16514; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16515; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16516; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16517; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16518; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16519; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16520; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16521; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16522; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16523; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16524; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16525; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd8;
#10 addr = 20'd16526; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16527; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16528; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd16529; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd11;
#10 addr = 20'd16530; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd16531; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16532; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16533; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16534; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16535; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16536; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16537; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd16538; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16539; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16540; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd9;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd16541; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16542; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16543; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16544; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd16545; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16546; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16547; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16548; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16549; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16550; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16551; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16552; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16553; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16554; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16555; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16556; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16557; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16558; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16559; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16560; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16561; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16562; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16563; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16564; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16565; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16566; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16567; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16568; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd16569; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16570; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16571; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16572; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd16573; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16574; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16575; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16576; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16577; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16578; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16579; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16580; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd16581; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd16582; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16583; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16584; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd8;data_in[15:12] = 4'd3;data_in[19:16] = 4'd3;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16585; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16586; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16587; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16588; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16589; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16590; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16591; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16592; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16593; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16594; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16595; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16596; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd16597; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16598; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16599; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16600; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd16601; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16602; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16603; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16604; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16605; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16606; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16607; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16608; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd5;
#10 addr = 20'd16609; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd16610; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16611; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16612; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd16613; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16614; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16615; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16616; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16617; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16618; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16619; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16620; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16621; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16622; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16623; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16624; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd16625; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16626; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16627; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16628; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd16629; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16630; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16631; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16632; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16633; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16634; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16635; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16636; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd16637; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16638; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16639; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16640; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd3;data_in[27:24] = 4'd4;data_in[31:28] = 4'd9;
#10 addr = 20'd16641; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16642; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd14;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16643; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16644; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16645; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16646; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16647; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16648; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16649; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16650; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16651; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16652; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd16653; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16654; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16655; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16656; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16657; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16658; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16659; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16660; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16661; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16662; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16663; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16664; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16665; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16666; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16667; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd16668; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd12;
#10 addr = 20'd16669; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16670; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd9;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16671; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16672; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16673; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16674; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16675; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16676; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16677; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16678; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16679; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16680; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd16681; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16682; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16683; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16684; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd16685; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16686; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16687; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16688; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16689; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16690; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16691; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16692; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16693; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16694; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16695; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd11;
#10 addr = 20'd16696; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd16697; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd16698; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16699; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16700; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16701; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16702; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16703; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16704; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16705; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16706; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16707; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16708; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd16709; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16710; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16711; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16712; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd16713; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16714; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16715; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16716; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16717; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16718; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16719; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16720; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16721; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16722; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd16723; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16724; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd16725; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16726; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16727; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16728; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16729; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16730; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16731; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16732; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16733; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16734; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16735; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16736; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16737; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16738; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16739; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16740; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd16741; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16742; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16743; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16744; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16745; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16746; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16747; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16748; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16749; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16750; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16751; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd16752; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16753; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd13;data_in[31:28] = 4'd7;
#10 addr = 20'd16754; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16755; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16756; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16757; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16758; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16759; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16760; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16761; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16762; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16763; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16764; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16765; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16766; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16767; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16768; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16769; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16770; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16771; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16772; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16773; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16774; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16775; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16776; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16777; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16778; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16779; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd16780; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16781; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd16782; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16783; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16784; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16785; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16786; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16787; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16788; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16789; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16790; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16791; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16792; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd16793; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16794; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16795; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16796; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16797; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16798; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16799; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16800; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16801; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16802; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16803; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16804; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16805; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16806; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16807; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16808; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16809; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd16810; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16811; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16812; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16813; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16814; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16815; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16816; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16817; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd7;
#10 addr = 20'd16818; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16819; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16820; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd16821; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16822; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16823; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16824; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16825; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16826; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16827; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16828; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16829; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16830; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16831; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd16832; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16833; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16834; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16835; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16836; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16837; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd16838; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16839; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16840; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16841; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16842; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16843; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16844; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd16845; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd16846; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16847; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16848; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd16849; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16850; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16851; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16852; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16853; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16854; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16855; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16856; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16857; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16858; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16859; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd16860; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16861; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16862; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16863; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16864; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd16865; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16866; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16867; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16868; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16869; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16870; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd16871; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16872; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16873; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd16874; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16875; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16876; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16877; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16878; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16879; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16880; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16881; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16882; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16883; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16884; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16885; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16886; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16887; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd9;
#10 addr = 20'd16888; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16889; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16890; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16891; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16892; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd10;
#10 addr = 20'd16893; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16894; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd16895; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16896; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16897; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16898; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16899; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16900; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16901; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16902; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16903; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16904; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16905; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16906; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16907; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16908; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16909; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16910; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16911; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16912; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16913; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16914; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16915; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16916; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16917; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd16918; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16919; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd16920; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd16921; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd16922; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16923; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16924; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16925; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16926; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16927; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16928; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16929; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16930; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16931; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16932; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16933; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16934; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16935; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16936; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16937; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16938; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16939; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16940; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16941; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16942; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16943; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16944; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16945; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16946; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16947; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd16948; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd16949; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16950; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16951; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16952; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16953; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16954; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16955; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16956; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd16957; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16958; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16959; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16960; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16961; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16962; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16963; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd16964; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16965; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16966; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16967; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16968; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd16969; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16970; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16971; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd16972; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd16973; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd16974; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16975; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd16976; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd16977; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd10;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd16978; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16979; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd16980; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16981; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16982; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16983; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd16984; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16985; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd16986; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd16987; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd16988; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd16989; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16990; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd16991; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd16992; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd16993; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16994; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd16995; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd16996; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd16997; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd16998; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd16999; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17000; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17001; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17002; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17003; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd17004; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd17005; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17006; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17007; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17008; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17009; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17010; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17011; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17012; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17013; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17014; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17015; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17016; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17017; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17018; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17019; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17020; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17021; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17022; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17023; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17024; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17025; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17026; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17027; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17028; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd17029; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17030; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17031; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17032; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd17033; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17034; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17035; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17036; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17037; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17038; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17039; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd17040; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd17041; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17042; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17043; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17044; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17045; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17046; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17047; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17048; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17049; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17050; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17051; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17052; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17053; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17054; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17055; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17056; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17057; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17058; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17059; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17060; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd7;
#10 addr = 20'd17061; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17062; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17063; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17064; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17065; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17066; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17067; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd17068; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17069; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17070; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17071; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17072; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17073; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17074; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17075; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17076; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17077; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17078; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17079; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17080; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17081; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17082; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17083; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17084; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17085; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17086; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17087; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd8;
#10 addr = 20'd17088; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17089; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17090; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17091; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17092; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17093; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17094; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17095; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17096; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17097; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17098; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17099; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17100; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17101; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17102; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17103; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17104; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17105; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17106; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17107; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17108; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17109; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17110; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17111; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17112; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17113; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17114; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17115; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17116; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17117; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17118; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17119; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17120; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17121; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17122; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17123; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17124; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17125; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17126; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17127; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17128; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17129; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17130; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17131; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17132; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17133; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17134; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17135; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17136; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17137; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17138; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17139; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17140; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17141; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17142; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17143; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd17144; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17145; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17146; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17147; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17148; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17149; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17150; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17151; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17152; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17153; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17154; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17155; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17156; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17157; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17158; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17159; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17160; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17161; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17162; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17163; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17164; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17165; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17166; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17167; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17168; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17169; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17170; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd17171; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17172; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17173; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17174; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17175; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17176; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17177; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17178; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17179; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17180; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17181; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17182; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17183; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17184; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17185; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17186; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17187; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17188; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17189; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17190; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17191; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17192; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17193; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17194; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17195; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17196; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17197; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17198; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17199; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd17200; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17201; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17202; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17203; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17204; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17205; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17206; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17207; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17208; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd17209; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17210; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17211; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17212; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17213; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17214; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17215; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17216; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17217; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17218; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17219; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd17220; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17221; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17222; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17223; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17224; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17225; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17226; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17227; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd17228; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17229; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17230; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17231; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17232; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17233; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17234; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17235; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17236; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17237; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17238; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17239; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17240; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17241; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17242; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17243; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17244; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17245; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17246; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17247; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17248; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17249; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17250; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17251; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd17252; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17253; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17254; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17255; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd17256; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd4;
#10 addr = 20'd17257; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17258; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17259; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17260; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17261; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17262; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17263; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17264; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17265; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17266; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17267; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17268; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd17269; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17270; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17271; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17272; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17273; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17274; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17275; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17276; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17277; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17278; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17279; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd17280; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17281; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17282; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd17283; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd17284; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd17285; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17286; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17287; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17288; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17289; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17290; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17291; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17292; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd17293; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17294; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17295; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17296; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd17297; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17298; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17299; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17300; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd12;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17301; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17302; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd17303; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17304; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17305; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17306; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17307; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd14;data_in[31:28] = 4'd10;
#10 addr = 20'd17308; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17309; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17310; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17311; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17312; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd17313; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17314; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17315; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17316; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17317; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17318; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17319; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17320; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd17321; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17322; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17323; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17324; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17325; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17326; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17327; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17328; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17329; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17330; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd17331; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17332; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17333; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17334; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17335; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd14;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17336; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17337; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17338; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17339; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17340; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd10;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17341; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd3;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17342; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17343; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17344; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17345; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17346; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17347; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17348; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17349; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd9;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17350; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17351; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17352; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17353; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17354; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17355; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17356; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17357; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17358; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd17359; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17360; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17361; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17362; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17363; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17364; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17365; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17366; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17367; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17368; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17369; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17370; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17371; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17372; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17373; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17374; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17375; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17376; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17377; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd17378; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17379; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17380; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd11;
#10 addr = 20'd17381; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17382; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17383; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17384; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17385; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17386; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17387; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17388; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17389; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17390; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17391; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17392; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17393; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17394; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17395; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17396; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17397; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17398; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17399; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17400; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17401; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17402; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17403; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17404; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17405; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd17406; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17407; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17408; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17409; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17410; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17411; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17412; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17413; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17414; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17415; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17416; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17417; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17418; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17419; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd17420; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd17421; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17422; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17423; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17424; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd9;
#10 addr = 20'd17425; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17426; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17427; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17428; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17429; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17430; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17431; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17432; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17433; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17434; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17435; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17436; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17437; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17438; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17439; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17440; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17441; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17442; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17443; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17444; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17445; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17446; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17447; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd17448; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17449; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd17450; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17451; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17452; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd8;
#10 addr = 20'd17453; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17454; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17455; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17456; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17457; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17458; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17459; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17460; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17461; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17462; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd8;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17463; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17464; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17465; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17466; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17467; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17468; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17469; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17470; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17471; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17472; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17473; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17474; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17475; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd17476; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17477; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd3;data_in[15:12] = 4'd3;data_in[19:16] = 4'd4;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17478; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17479; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17480; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17481; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17482; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17483; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17484; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17485; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17486; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17487; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17488; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17489; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17490; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd17491; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17492; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17493; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17494; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17495; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17496; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17497; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17498; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17499; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17500; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17501; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17502; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17503; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17504; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd17505; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17506; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17507; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17508; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd17509; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17510; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17511; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17512; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17513; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17514; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17515; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17516; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17517; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17518; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17519; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17520; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17521; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17522; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17523; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17524; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17525; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd17526; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17527; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17528; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17529; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17530; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17531; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17532; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd17533; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17534; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd17535; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17536; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd17537; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17538; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17539; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17540; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17541; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17542; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17543; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17544; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17545; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17546; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd6;
#10 addr = 20'd17547; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17548; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17549; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17550; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17551; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17552; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17553; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd11;
#10 addr = 20'd17554; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17555; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17556; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17557; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17558; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17559; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17560; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17561; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17562; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd17563; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17564; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd3;
#10 addr = 20'd17565; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd12;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17566; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17567; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17568; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17569; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17570; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17571; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17572; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17573; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17574; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd12;
#10 addr = 20'd17575; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17576; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17577; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17578; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17579; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17580; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17581; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd10;
#10 addr = 20'd17582; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17583; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17584; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17585; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17586; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17587; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd7;
#10 addr = 20'd17588; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17589; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17590; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17591; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17592; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd17593; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17594; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17595; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17596; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17597; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17598; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17599; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17600; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17601; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17602; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17603; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17604; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd10;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17605; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17606; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17607; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17608; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17609; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd8;
#10 addr = 20'd17610; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17611; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17612; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17613; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd9;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17614; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17615; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd17616; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17617; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17618; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd17619; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd17620; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17621; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd11;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17622; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17623; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17624; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17625; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17626; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17627; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17628; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17629; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17630; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17631; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd11;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd17632; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17633; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17634; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17635; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17636; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17637; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd17638; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17639; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17640; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17641; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd17642; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17643; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17644; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17645; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17646; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd17647; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17648; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17649; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd12;data_in[19:16] = 4'd5;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd17650; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17651; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17652; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd17653; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17654; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17655; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17656; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17657; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17658; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17659; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17660; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17661; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17662; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17663; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17664; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17665; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd17666; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17667; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17668; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17669; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd17670; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17671; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17672; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17673; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17674; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd17675; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17676; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd17677; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd17678; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17679; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17680; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17681; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17682; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17683; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17684; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17685; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17686; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17687; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17688; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17689; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17690; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17691; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17692; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17693; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17694; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd17695; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17696; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17697; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17698; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17699; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17700; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17701; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17702; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17703; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17704; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd17705; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd6;data_in[11:8] = 4'd3;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd4;
#10 addr = 20'd17706; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17707; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17708; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17709; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17710; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17711; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17712; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17713; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17714; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17715; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd11;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17716; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17717; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17718; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17719; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17720; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17721; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17722; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17723; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17724; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17725; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17726; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17727; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17728; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17729; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17730; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17731; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17732; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd17733; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd4;
#10 addr = 20'd17734; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17735; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17736; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd17737; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17738; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17739; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17740; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17741; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17742; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17743; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17744; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17745; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17746; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17747; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17748; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17749; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17750; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17751; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17752; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17753; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17754; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17755; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd17756; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17757; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd17758; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17759; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17760; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17761; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd4;
#10 addr = 20'd17762; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17763; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17764; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd17765; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17766; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17767; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17768; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17769; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17770; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17771; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd11;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17772; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17773; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17774; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17775; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17776; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17777; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17778; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17779; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17780; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17781; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17782; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17783; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd17784; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17785; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd4;
#10 addr = 20'd17786; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17787; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17788; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17789; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd17790; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17791; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17792; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd17793; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17794; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17795; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17796; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17797; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17798; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17799; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17800; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd9;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17801; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17802; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17803; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17804; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17805; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17806; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17807; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17808; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17809; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17810; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17811; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17812; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17813; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd17814; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17815; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17816; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd17817; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd9;data_in[23:20] = 4'd12;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd17818; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17819; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17820; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd17821; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17822; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17823; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17824; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17825; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17826; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17827; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd10;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17828; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd10;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17829; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17830; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17831; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17832; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17833; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17834; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17835; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17836; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17837; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17838; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17839; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17840; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17841; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd8;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd17842; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17843; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17844; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17845; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd17846; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17847; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17848; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd17849; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17850; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17851; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17852; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17853; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17854; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17855; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd17856; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17857; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17858; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17859; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17860; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17861; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd17862; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17863; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17864; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17865; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17866; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17867; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd17868; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17869; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd4;
#10 addr = 20'd17870; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17871; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd17872; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17873; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd10;
#10 addr = 20'd17874; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17875; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd17876; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd17877; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17878; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17879; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17880; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17881; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17882; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17883; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd7;data_in[31:28] = 4'd3;
#10 addr = 20'd17884; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17885; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17886; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17887; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17888; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17889; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17890; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17891; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17892; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17893; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd17894; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17895; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17896; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17897; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd17898; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17899; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd17900; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17901; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd17902; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17903; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd17904; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd6;
#10 addr = 20'd17905; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17906; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17907; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17908; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17909; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17910; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17911; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd10;data_in[31:28] = 4'd4;
#10 addr = 20'd17912; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17913; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17914; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd17915; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17916; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17917; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17918; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17919; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17920; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17921; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd14;
#10 addr = 20'd17922; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17923; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd17924; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17925; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd17926; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17927; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd17928; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd17929; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd5;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd17930; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17931; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17932; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd17933; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17934; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17935; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17936; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17937; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17938; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17939; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd5;
#10 addr = 20'd17940; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17941; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17942; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17943; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17944; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17945; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17946; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17947; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17948; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17949; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd14;
#10 addr = 20'd17950; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17951; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17952; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17953; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd17954; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17955; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd17956; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17957; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd17958; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17959; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17960; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17961; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17962; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17963; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17964; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd17965; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17966; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17967; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd6;
#10 addr = 20'd17968; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd7;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd17969; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17970; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17971; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd17972; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd17973; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17974; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd17975; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd17976; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd17977; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd17978; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17979; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd17980; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd17981; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd17982; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd17983; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd17984; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd17985; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd17986; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd17987; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd17988; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd17989; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17990; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17991; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17992; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd17993; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd17994; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd17995; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd9;
#10 addr = 20'd17996; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd8;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd17997; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd17998; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd17999; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18000; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd18001; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18002; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18003; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18004; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18005; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18006; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18007; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18008; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18009; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18010; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18011; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd18012; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18013; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd18014; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18015; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18016; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18017; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18018; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18019; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18020; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18021; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18022; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18023; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd11;
#10 addr = 20'd18024; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18025; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18026; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18027; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18028; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd13;
#10 addr = 20'd18029; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18030; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18031; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18032; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18033; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18034; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18035; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18036; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18037; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18038; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18039; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18040; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd18041; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd18042; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18043; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18044; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18045; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18046; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18047; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18048; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18049; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18050; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18051; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd14;
#10 addr = 20'd18052; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18053; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18054; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18055; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18056; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18057; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18058; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18059; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18060; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18061; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd14;
#10 addr = 20'd18062; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18063; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18064; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18065; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18066; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd18067; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18068; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18069; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd18070; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18071; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18072; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18073; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18074; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18075; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18076; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18077; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18078; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18079; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18080; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18081; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18082; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18083; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18084; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18085; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18086; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18087; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18088; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd7;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18089; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18090; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18091; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18092; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18093; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18094; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd18095; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd4;
#10 addr = 20'd18096; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18097; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18098; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18099; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18100; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18101; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18102; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18103; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18104; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18105; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18106; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18107; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18108; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18109; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18110; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18111; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18112; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd18113; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18114; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18115; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18116; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18117; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18118; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18119; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18120; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18121; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18122; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18123; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd18124; we = 1; data_in[3:0] = 4'd3;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18125; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd18126; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18127; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18128; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18129; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18130; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18131; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18132; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18133; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18134; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18135; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18136; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd11;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18137; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18138; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18139; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd18140; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd18141; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18142; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18143; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18144; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18145; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18146; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18147; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18148; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18149; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18150; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18151; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18152; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18153; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd18154; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18155; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18156; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd18157; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18158; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18159; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18160; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18161; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18162; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18163; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18164; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18165; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18166; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18167; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd18168; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd18169; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18170; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18171; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18172; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18173; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18174; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18175; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18176; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18177; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18178; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd18179; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18180; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd5;
#10 addr = 20'd18181; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18182; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18183; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18184; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd18185; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18186; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18187; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18188; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18189; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18190; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18191; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18192; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18193; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18194; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18195; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd14;
#10 addr = 20'd18196; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18197; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18198; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18199; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18200; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18201; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18202; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18203; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18204; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18205; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18206; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd18207; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18208; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18209; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18210; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18211; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18212; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd18213; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18214; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18215; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18216; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18217; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18218; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18219; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18220; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18221; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18222; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18223; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18224; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18225; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18226; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18227; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18228; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18229; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18230; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18231; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18232; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18233; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18234; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18235; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18236; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18237; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18238; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18239; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18240; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18241; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18242; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18243; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18244; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18245; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18246; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18247; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18248; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18249; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18250; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd18251; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd18252; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd18253; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18254; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18255; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18256; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18257; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd9;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18258; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18259; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd11;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18260; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18261; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18262; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18263; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18264; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18265; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18266; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18267; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18268; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd10;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd13;
#10 addr = 20'd18269; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18270; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18271; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18272; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18273; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18274; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18275; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18276; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18277; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18278; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18279; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd15;
#10 addr = 20'd18280; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18281; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18282; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18283; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18284; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18285; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd18286; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18287; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18288; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18289; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18290; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18291; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18292; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18293; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18294; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18295; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18296; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd11;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd18297; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18298; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18299; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18300; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18301; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18302; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18303; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18304; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18305; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18306; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18307; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18308; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd12;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18309; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18310; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18311; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18312; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18313; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd18314; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18315; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18316; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18317; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18318; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18319; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd18320; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18321; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18322; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18323; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18324; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd8;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18325; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18326; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18327; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18328; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18329; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18330; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18331; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18332; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd13;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18333; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18334; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18335; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18336; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18337; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18338; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18339; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18340; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18341; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18342; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18343; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18344; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18345; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18346; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18347; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd5;
#10 addr = 20'd18348; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18349; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18350; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18351; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18352; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd8;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18353; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18354; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18355; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18356; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18357; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18358; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18359; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18360; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18361; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18362; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd18363; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18364; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18365; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18366; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18367; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18368; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18369; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd18370; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18371; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18372; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18373; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18374; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18375; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd18376; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18377; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18378; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18379; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18380; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd10;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18381; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18382; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18383; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18384; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18385; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18386; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18387; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18388; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18389; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18390; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd18391; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18392; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18393; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18394; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18395; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18396; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18397; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd13;
#10 addr = 20'd18398; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18399; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18400; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18401; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18402; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18403; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18404; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd9;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18405; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18406; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18407; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd10;data_in[31:28] = 4'd6;
#10 addr = 20'd18408; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd9;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18409; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18410; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18411; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18412; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18413; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18414; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18415; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18416; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd12;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18417; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18418; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd10;
#10 addr = 20'd18419; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18420; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd13;data_in[11:8] = 4'd10;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18421; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18422; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18423; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18424; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18425; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18426; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18427; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd8;data_in[31:28] = 4'd5;
#10 addr = 20'd18428; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18429; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18430; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18431; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18432; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18433; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18434; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18435; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd10;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd18436; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18437; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18438; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18439; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18440; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18441; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18442; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18443; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18444; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18445; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18446; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd10;
#10 addr = 20'd18447; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18448; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd10;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18449; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18450; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18451; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18452; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18453; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18454; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18455; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18456; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18457; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18458; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18459; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18460; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18461; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18462; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18463; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd8;data_in[23:20] = 4'd5;data_in[27:24] = 4'd4;data_in[31:28] = 4'd7;
#10 addr = 20'd18464; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18465; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18466; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18467; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18468; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18469; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18470; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18471; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18472; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18473; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18474; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd18475; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18476; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd8;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18477; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18478; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18479; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18480; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18481; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18482; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18483; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd18484; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18485; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18486; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18487; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18488; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd10;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18489; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18490; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18491; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd18492; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18493; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18494; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18495; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18496; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18497; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18498; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18499; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18500; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd12;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18501; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18502; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd18503; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd18504; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18505; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18506; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18507; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18508; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18509; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18510; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18511; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd4;
#10 addr = 20'd18512; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18513; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18514; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18515; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18516; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18517; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18518; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18519; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18520; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18521; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18522; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18523; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18524; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18525; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18526; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18527; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18528; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd13;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18529; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18530; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd18531; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd15;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd11;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18532; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18533; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18534; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18535; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18536; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd18537; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd8;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18538; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18539; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd10;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18540; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18541; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18542; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18543; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd4;data_in[11:8] = 4'd8;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18544; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd11;data_in[27:24] = 4'd7;data_in[31:28] = 4'd5;
#10 addr = 20'd18545; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18546; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18547; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd8;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd12;
#10 addr = 20'd18548; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18549; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18550; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18551; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18552; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18553; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18554; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18555; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18556; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18557; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18558; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18559; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18560; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18561; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18562; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18563; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18564; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd11;
#10 addr = 20'd18565; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18566; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18567; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18568; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18569; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18570; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18571; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd18572; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd7;
#10 addr = 20'd18573; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18574; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18575; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18576; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18577; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18578; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18579; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18580; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18581; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18582; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18583; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18584; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd15;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd11;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18585; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18586; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18587; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18588; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18589; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18590; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18591; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18592; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18593; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18594; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18595; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd12;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18596; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18597; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18598; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18599; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd9;data_in[19:16] = 4'd5;data_in[23:20] = 4'd3;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd18600; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18601; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18602; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18603; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd18604; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18605; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18606; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18607; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18608; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18609; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18610; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18611; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18612; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd12;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18613; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18614; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18615; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18616; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18617; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18618; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18619; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18620; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18621; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18622; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18623; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18624; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18625; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd4;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18626; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd18627; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd4;data_in[11:8] = 4'd6;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd4;data_in[27:24] = 4'd4;data_in[31:28] = 4'd6;
#10 addr = 20'd18628; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd6;data_in[31:28] = 4'd8;
#10 addr = 20'd18629; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18630; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18631; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18632; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18633; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18634; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18635; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18636; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18637; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18638; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18639; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18640; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd13;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18641; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18642; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18643; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18644; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18645; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18646; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18647; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18648; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd10;
#10 addr = 20'd18649; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd12;data_in[19:16] = 4'd11;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18650; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd15;data_in[31:28] = 4'd15;
#10 addr = 20'd18651; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18652; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18653; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd7;
#10 addr = 20'd18654; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18655; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd4;data_in[11:8] = 4'd5;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd3;data_in[31:28] = 4'd5;
#10 addr = 20'd18656; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd6;
#10 addr = 20'd18657; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18658; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd11;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18659; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18660; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18661; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18662; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18663; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18664; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18665; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18666; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18667; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18668; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd9;data_in[31:28] = 4'd7;
#10 addr = 20'd18669; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd9;
#10 addr = 20'd18670; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18671; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd10;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18672; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18673; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18674; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18675; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18676; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd11;
#10 addr = 20'd18677; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd12;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18678; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18679; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18680; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18681; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd6;data_in[23:20] = 4'd4;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd18682; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd10;
#10 addr = 20'd18683; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd3;
#10 addr = 20'd18684; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd4;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd6;
#10 addr = 20'd18685; we = 1; data_in[3:0] = 4'd4;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18686; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd10;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18687; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18688; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18689; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18690; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18691; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18692; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18693; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18694; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18695; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18696; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd11;data_in[31:28] = 4'd7;
#10 addr = 20'd18697; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18698; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18699; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18700; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18701; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd9;
#10 addr = 20'd18702; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd10;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18703; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18704; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd12;
#10 addr = 20'd18705; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18706; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18707; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18708; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18709; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd18710; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd9;
#10 addr = 20'd18711; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd5;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18712; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd8;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18713; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd5;data_in[19:16] = 4'd4;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18714; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18715; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18716; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18717; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18718; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18719; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18720; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18721; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18722; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18723; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18724; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd15;data_in[19:16] = 4'd14;data_in[23:20] = 4'd15;data_in[27:24] = 4'd12;data_in[31:28] = 4'd7;
#10 addr = 20'd18725; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18726; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd11;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
#10 addr = 20'd18727; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18728; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18729; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18730; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd8;data_in[27:24] = 4'd7;data_in[31:28] = 4'd7;
#10 addr = 20'd18731; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd8;
#10 addr = 20'd18732; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd9;data_in[31:28] = 4'd13;
#10 addr = 20'd18733; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18734; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18735; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd12;data_in[15:12] = 4'd11;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18736; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd6;
#10 addr = 20'd18737; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd7;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd9;
#10 addr = 20'd18738; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd5;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18739; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd7;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd6;
#10 addr = 20'd18740; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd7;
#10 addr = 20'd18741; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd9;data_in[11:8] = 4'd5;data_in[15:12] = 4'd4;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18742; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd11;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18743; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd18744; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18745; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18746; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18747; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18748; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18749; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18750; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd13;
#10 addr = 20'd18751; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18752; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd13;data_in[31:28] = 4'd8;
#10 addr = 20'd18753; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd9;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18754; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd11;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18755; we = 1; data_in[3:0] = 4'd11;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd11;
#10 addr = 20'd18756; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18757; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18758; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd10;data_in[15:12] = 4'd9;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd7;data_in[31:28] = 4'd6;
#10 addr = 20'd18759; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd10;
#10 addr = 20'd18760; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd18761; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18762; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd15;
#10 addr = 20'd18763; we = 1; data_in[3:0] = 4'd15;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18764; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18765; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd5;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd7;data_in[31:28] = 4'd9;
#10 addr = 20'd18766; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18767; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd9;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18768; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18769; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd8;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18770; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd13;
#10 addr = 20'd18771; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18772; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18773; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18774; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd14;
#10 addr = 20'd18775; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18776; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18777; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18778; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd13;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18779; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18780; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd10;
#10 addr = 20'd18781; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18782; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18783; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd18784; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18785; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18786; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18787; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd6;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd10;data_in[31:28] = 4'd10;
#10 addr = 20'd18788; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd5;data_in[11:8] = 4'd6;data_in[15:12] = 4'd5;data_in[19:16] = 4'd5;data_in[23:20] = 4'd5;data_in[27:24] = 4'd8;data_in[31:28] = 4'd12;
#10 addr = 20'd18789; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd11;data_in[27:24] = 4'd10;data_in[31:28] = 4'd12;
#10 addr = 20'd18790; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18791; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd11;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd4;
#10 addr = 20'd18792; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd4;data_in[15:12] = 4'd6;data_in[19:16] = 4'd5;data_in[23:20] = 4'd7;data_in[27:24] = 4'd6;data_in[31:28] = 4'd7;
#10 addr = 20'd18793; we = 1; data_in[3:0] = 4'd7;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd7;data_in[27:24] = 4'd9;data_in[31:28] = 4'd8;
#10 addr = 20'd18794; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd6;data_in[11:8] = 4'd5;data_in[15:12] = 4'd7;data_in[19:16] = 4'd9;data_in[23:20] = 4'd6;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd18795; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd8;data_in[11:8] = 4'd9;data_in[15:12] = 4'd5;data_in[19:16] = 4'd8;data_in[23:20] = 4'd8;data_in[27:24] = 4'd5;data_in[31:28] = 4'd5;
#10 addr = 20'd18796; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd7;data_in[15:12] = 4'd6;data_in[19:16] = 4'd6;data_in[23:20] = 4'd5;data_in[27:24] = 4'd5;data_in[31:28] = 4'd8;
#10 addr = 20'd18797; we = 1; data_in[3:0] = 4'd6;data_in[7:4] = 4'd7;data_in[11:8] = 4'd7;data_in[15:12] = 4'd8;data_in[19:16] = 4'd7;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18798; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd11;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18799; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd12;
#10 addr = 20'd18800; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18801; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18802; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd13;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd14;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18803; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd13;data_in[31:28] = 4'd13;
#10 addr = 20'd18804; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18805; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18806; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd13;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18807; we = 1; data_in[3:0] = 4'd13;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd14;data_in[23:20] = 4'd14;data_in[27:24] = 4'd14;data_in[31:28] = 4'd14;
#10 addr = 20'd18808; we = 1; data_in[3:0] = 4'd14;data_in[7:4] = 4'd14;data_in[11:8] = 4'd14;data_in[15:12] = 4'd14;data_in[19:16] = 4'd15;data_in[23:20] = 4'd15;data_in[27:24] = 4'd14;data_in[31:28] = 4'd12;
#10 addr = 20'd18809; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd8;data_in[23:20] = 4'd9;data_in[27:24] = 4'd9;data_in[31:28] = 4'd9;
#10 addr = 20'd18810; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd11;data_in[11:8] = 4'd12;data_in[15:12] = 4'd12;data_in[19:16] = 4'd12;data_in[23:20] = 4'd12;data_in[27:24] = 4'd12;data_in[31:28] = 4'd12;
#10 addr = 20'd18811; we = 1; data_in[3:0] = 4'd12;data_in[7:4] = 4'd12;data_in[11:8] = 4'd13;data_in[15:12] = 4'd13;data_in[19:16] = 4'd13;data_in[23:20] = 4'd12;data_in[27:24] = 4'd11;data_in[31:28] = 4'd10;
#10 addr = 20'd18812; we = 1; data_in[3:0] = 4'd9;data_in[7:4] = 4'd9;data_in[11:8] = 4'd8;data_in[15:12] = 4'd7;data_in[19:16] = 4'd7;data_in[23:20] = 4'd7;data_in[27:24] = 4'd8;data_in[31:28] = 4'd8;
#10 addr = 20'd18813; we = 1; data_in[3:0] = 4'd8;data_in[7:4] = 4'd8;data_in[11:8] = 4'd8;data_in[15:12] = 4'd8;data_in[19:16] = 4'd9;data_in[23:20] = 4'd10;data_in[27:24] = 4'd10;data_in[31:28] = 4'd11;
#10 addr = 20'd18814; we = 1; data_in[3:0] = 4'd10;data_in[7:4] = 4'd10;data_in[11:8] = 4'd9;data_in[15:12] = 4'd8;data_in[19:16] = 4'd6;data_in[23:20] = 4'd6;data_in[27:24] = 4'd6;data_in[31:28] = 4'd5;
#10 addr = 20'd18815; we = 1; data_in[3:0] = 4'd5;data_in[7:4] = 4'd6;data_in[11:8] = 4'd6;data_in[15:12] = 4'd7;data_in[19:16] = 4'd8;data_in[23:20] = 4'd10;data_in[27:24] = 4'd11;data_in[31:28] = 4'd11;
    
    // Finish the simulation
    #10 $finish;
  end
endmodule
