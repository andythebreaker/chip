`include "vmvmb.sv"

    //========== this a testbench driven by 6 data in a group from python gen txt =========
    module tb;
    logic signed [31:0] x[0:99];
    logic signed [31:0] Wx[0:99][0:399];
    logic signed [31:0] h_prev[0:99];
    logic signed [31:0] Wh[0:99][0:399];
    logic signed [31:0] b[0:399];
    logic signed [31:0] A[0:399];
    vmvmb dut(
        x,Wx,h_prev,Wh,b,A
    );
    initial begin
        $fsdbDumpfile("tb_6data.fsdb");
        $fsdbDumpvars("+all");
    end
    initial begin
    #10;
    x='{2330,2047,-49,-2961,-54,480,-1728,-1111,2214,-9575,993,4052,-3518,-3215,430,2386,-1245,1867,330,1953,-4775,3457,-2783,1555,2954,-2602,-1588,2763,-4379,6376,-815,3034,-2458,-523,-392,-2536,-1047,-1115,516,-577,12,4538,-1199,2971,-2912,3154,4538,2980,-897,1973,-2158,1784,4509,-113,-3269,-2697,-4052,-2844,-5234,-1096,-203,1050,3071,4003,-777,2778,1890,298,178,-4899,1799,-2454,5170,-3618,-5302,-1679,-123,3493,3388,5361,-754,3559,-3815,4370,-1448,-4143,-720,-1811,1986,-2951,563,1052,745,2186,4262,-846,-1157,262,249,-4721};
    h_prev='{0,7531,-31,536,5,-11,-345,-3206,655,1300,-150,-1578,545,3005,0,1619,6694,1093,-451,43,49,5,-690,2,0,-3087,0,4420,-297,-634,386,6774,253,-4078,43,-16,8,596,-6244,-5694,-124,6721,-6314,-7489,-4378,7047,1937,576,-345,-1097,7322,-7510,443,6400,-310,-1839,-3803,-35,-647,6255,615,-26,-3230,398,-848,0,-2154,7441,-576,-57,257,-7257,-25,-5635,1,-56,-7604,5018,873,-4056,9,7315,-107,-7266,0,5227,-53,1492,-638,6954,-2,-978,-278,4962,926,-3516,628,41,86,-5108};
    b='{2325,-16591,-5761,-12939,-2268,8706,-14824,-7407,1971,-6577,-8862,3022,1065,-15878,-7822,-8212,-12353,13,-2687,-8769,816,-7163,-5839,-8320,-1706,-406,-5483,-1447,-5449,-2780,-4860,-11816,-14082,-8930,30156,-7968,13271,-3193,-9770,-15302,1127,-25781,23574,-13740,-2033,-680,-20019,2381,-14257,33281,-10078,-16669,5009,13349,5454,16015,-8173,911,-10722,16494,-1926,-9931,-13828,1466,-125,-4362,3579,-21718,42,-3796,25058,-19199,-13105,-16464,-3146,-6401,-6411,-9160,36113,1428,-5668,-23535,-12744,-22968,2939,-15312,-1862,-7666,8647,1607,-6269,-16708,-11044,-22578,-25273,-7495,2443,-21816,-8652,-11708,-2158,5581,-11201,4299,5498,-12734,-22167,-13652,12119,-9165,-7456,2143,875,1092,-1405,11923,-6508,-10478,-10673,3737,15556,4450,-2470,-2175,-7202,9233,-4433,-5571,1979,-5434,-6669,-9204,10234,9111,35332,15410,14570,8989,5957,-7246,-5693,-621,3356,15781,-6186,2531,22500,10458,2587,-2441,-10810,-20,9965,-4663,-13378,-7387,13769,-17402,-12050,10888,-11406,-7739,2778,-18427,4763,-8984,-13447,-11982,-18017,16992,5170,-9428,5800,-10996,10546,2462,-520,2225,6923,18095,13564,18623,-12714,5654,15625,909,-14062,7416,-11494,21191,-10449,-3354,-5722,28671,19765,-7260,12441,921,13,4580,-3010,11337,-35,-582,-1089,4050,5527,7456,-5185,-2135,9526,-8574,-12910,12626,9956,-7827,-3574,637,-10634,-10566,481,-3547,-9575,-3740,-5263,-5961,-8510,581,3078,-10800,-6459,6196,13212,6865,-20234,-5776,-22832,-262,14921,12695,-2697,11035,-8994,12646,-1105,5795,4804,-3356,-643,-25292,16640,10166,-4919,-7661,-15009,-7006,-5561,-1893,-1473,-23085,-15087,-5205,24472,-3608,7495,-12607,-6894,5776,1760,-3903,-26796,3188,-6088,8295,-4401,5615,612,11337,-27773,-4133,-6674,9150,-2237,21113,-863,8994,-5307,4187,-18476,103,-16796,25820,1778,7016,8984,930,-6279,12656,-8710,13720,-15244,26035,-34160,2376,-1462,-34628,-2639,10302,2487,-7680,8588,-2191,-16396,15078,18701,15185,23945,-715,-7021,-25820,-26542,-5571,-11767,-4133,-7934,-3090,-1916,-7265,4565,6542,-9467,18251,11855,15849,8735,-8808,6689,-10859,13847,16093,4677,20195,6220,4038,11347,7685,26074,3815,-10781,12343,22519,20742,-2722,12509,-6474,14277,-896,-34160,6064,-659,-14785,6728,12919,7866,16679,-25976,-11464,22382,-20390,-21054,2895,343,-11220,13896,-15517,8417,16220,10205,22402,-1508,-4157,27792,-2673,24042,-6416,17197,-10869,-672,-3002,-35761,-6186,6982,9575,-20820,16318,2413,-4609,27324,-9907,15625};
    Wx[0]='{1748,-2391,-84,-2595,-209,1027,-4772,-1782,-413,-1520,45,-1872,-1966,-1979,-526,5195,2395,-995,3034,159,374,-450,-1140,861,698,3110,509,560,-3002,-2878,124,-6796,813,3708,-253,-2749,548,1571,1977,-2110,273,4450,2651,4565,8852,-3347,-1206,3969,-1697,1602,-2812,558,-1474,4772,1049,-2697,-2244,4650,-5063,1347,3984,-2482,-862,-337,-4309,-708,-5053,12568,1018,-1983,-3234,-3654,2120,-8930,2741,2115,1712,-1268,-3627,-4992,1536,-3159,-319,935,109,-3535,426,-294,182,-2978,-2978,2917,-2316,-1596,870,-1390,-2846,-197,1804,-326,1583,6962,-1955,2944,4387,-2283,4411,-5000,3989,2934,1784,-5107,228,-5942,-8730,9541,-2150,6176,2575,2617,-3586,-5991,-4536,5209,-143,7387,-4245,3369,-14296,-2315,3391,-17060,7104,10263,-8037,1678,-416,-1987,28105,3261,3913,5102,9169,-9174,2028,2015,-6606,2050,-2495,3811,9936,1859,2335,4294,565,-4707,-539,-2788,-9370,-4548,-3381,1191,-20722,3979,-2504,1778,2271,-474,2880,1074,-3071,-8071,-2854,2395,2292,-733,-841,-7021,-4082,1253,435,8632,4997,-12705,-972,6191,-2617,2043,1710,-581,1738,14316,-1013,297,-5737,6621,-5258,1318,6606,2980,-1444,-1418,-916,1661,1507,-93,-5585,-5903,-288,-548,-3378,-5424,-5219,-5625,8593,6660,-1472,-5000,-3410,-4416,2408,433,-590,-541,-3034,-3247,-9838,-407,-10341,6596,-441,-3569,2214,1781,1525,-3254,-3762,1170,-3942,-2453,-182,2249,-3850,-3728,6162,-2399,-2829,-3703,272,-522,-4211,1148,-3193,2199,-3359,-2219,-6923,438,342,2124,336,-3952,-686,166,-11054,-650,-6704,422,3620,-2998,3195,1872,-1497,-1053,169,-6333,4965,-3796,-5019,2269,-1610,8442,497,-4912,-5034,-2641,1246,-2156,2364,-1135,-4892,376,4299,2954,1356,3378,-1019,-5283,-485,323,-2773,15,2834,-2497,520,-6713,-7416,2053,5898,78,-6425,-3461,-1616,-4121,385,4965,1895,-9873,1890,137,180,-1066,242,-2509,-4313,514,-5942,1334,-2377,1319,442,-3041,-2205,1828,6313,-5771,4162,7934,2741,-9667,3291,-3044,-5097,-990,-620,-2073,4191,2719,2023,-1494,-6391,-2124,-3437,130,413,-6918,-6210,6098,-2575,6240,2470,-4121,759,4123,-1907,-4995,-8745,1820,-1737,-9316,-3542,-3884,5810,-10664,3352,1601,1304,-4602,1939,4042,2287,1691,6450,-4123,-4870,-1944,2680,-955,2553,12402,-4328,-3818,-3901,13681,-2954,5732,-4650,5253,-911,391};
    Wx[1]='{-2021,792,-446,-1254,3015,2592,-2670,-2197,895,-872,5546,1298,-979,-1141,155,5888,8510,2963,-1262,-963,1883,4477,-2131,2548,3872,3259,1389,1835,-2279,4406,17,3405,-950,2327,-745,1199,-1387,563,-1486,-419,496,-636,-720,5898,-2249,2795,1356,-3088,2056,-2056,-7431,5249,-164,-3552,2687,8447,-5312,422,3210,66,6196,-5874,2478,718,3750,833,1325,-2285,-1298,1722,-1585,-42,-418,777,-995,3562,5908,2109,-882,1676,-1661,-778,5903,3464,-875,1605,1285,4020,3762,-385,-935,5019,2602,-1090,-1021,297,-2384,2312,-1245,6396,-3503,3107,-190,1981,1885,-832,1749,1257,-3190,-6499,4633,1876,-229,142,8466,-2770,3012,1375,-2010,-549,-1965,5166,2604,3222,4072,-2392,-1826,50,-2203,-3081,5249,22226,5556,1284,-1746,1431,2382,-7675,-8666,5214,-1248,-11318,-9062,4724,3200,-7836,15537,-11865,-5478,4738,-7329,-5522,5263,-9487,2330,-12861,-374,2102,4245,3220,1607,-7065,-16474,-2941,9692,11,-3347,7983,1732,-3784,-1051,1297,-2604,-3515,3391,-1973,-15302,-8378,-2105,6596,6220,15576,2475,-4357,-1325,-3288,1268,-7397,-1754,-1472,2266,-8457,4267,1472,9252,1516,1409,-553,-4443,-5703,739,-10156,1785,94,1374,-690,-898,-2218,-10400,978,-8500,-1187,1237,1070,-5078,-4675,-13300,7060,4013,1518,2719,894,9194,100,-3120,-2329,5366,-3132,-7001,-2293,-605,-4895,3251,-1917,6298,228,-4052,870,-4765,-8183,1215,364,2303,-2277,-75,-1030,-3066,4345,-294,-6401,-304,2834,-31,-6416,-2117,-3637,3088,4890,-9697,586,1417,-3977,3666,-1117,-309,-793,1115,-7539,888,-1911,-4365,-6132,515,-1495,-430,2724,-3422,1096,-2556,2008,5507,1337,-782,-5327,-3828,-4113,-4008,3022,-7719,-1665,5292,-5698,-2814,593,5439,-5908,3576,-13242,4179,-6132,5737,-6044,-4899,1315,7763,-1192,1078,27,-4416,7861,-579,-847,3249,891,-2332,-4953,-3508,6127,-3166,-1361,129,672,5971,4274,6464,-3962,519,-1973,2169,1781,-567,-3020,-11279,-6552,3303,-3452,247,1834,-8803,-13613,4926,1600,-3669,-6113,-80,-6196,2248,-842,484,-4118,-5087,-444,-6093,-2341,-6567,-276,-2138,6889,-5424,8012,4926,-8168,208,-2314,3068,8227,1760,2575,4440,634,-3950,475,-133,245,4145,-9858,6806,-3410,-4670,620,5307,-1348,-2932,-6074,8315,3569,115,-4050,17,8076,260,-10585,-3166,6669,-13056,-269,2232,10468,6459,-3510};
    Wx[2]='{-2290,5834,-2166,-440,833,-1110,3168,5678,-485,-415,3071,-838,6782,-2108,4978,3525,-8276,4807,2937,2111,1343,1026,-4538,3178,-138,1131,-487,1563,2829,8876,-2069,8051,1767,1799,-3918,-1702,4411,3222,869,2025,3349,-2124,-185,2006,-252,-538,-2990,2185,3715,665,3513,10585,1539,1430,2192,-251,4829,-1114,3605,2968,4682,1182,557,308,-292,-3881,-632,7373,906,221,-244,3442,515,6728,1580,-930,-3356,1623,-1708,-519,2061,2727,3024,-2180,-1903,5922,-3,2474,-1386,799,3984,3173,-4641,-345,3649,2763,3300,5034,3615,3964,-555,-8715,151,535,-3776,578,10400,-6596,-4194,-1437,6889,-8388,3774,-5229,-3168,-5537,2464,2568,-1842,5932,479,-144,2440,-6772,-4191,5112,-5405,-1348,-6533,12021,-235,13652,3164,-7055,580,-5629,-1439,7929,-2988,-9238,4506,718,-15126,-3625,-7993,-2722,9311,-1068,1965,-5830,1086,-7885,-6147,-10537,-999,-997,-8012,-1826,-7270,1997,-5468,828,-18730,2934,2498,341,8408,-12744,-1989,64,-834,-1106,-242,-12509,1473,-6748,-1668,12675,6235,1617,735,-131,-9379,-11376,7543,1028,-4384,-4885,-3337,-6665,3220,10820,1198,3732,-4594,6250,1644,-1787,-9589,-5815,-3078,-17617,-2973,-838,4348,-79,-8383,1903,3754,874,-5268,2390,2006,-419,-2656,-7290,-6718,-533,-384,4052,-1183,-2144,702,5053,-1557,-6967,1210,600,-8071,1557,2036,7934,-12822,-1376,-1237,-4863,-3986,913,-5961,-3244,152,-12929,1765,-996,-3713,2239,1749,-2374,-3466,-1414,7622,1099,-1239,-5830,-307,-4350,-6176,838,-10175,-3862,-2832,-5146,-1585,3793,1702,-8242,-1738,-6992,-527,-2473,44,-3898,-2780,-9721,88,-350,-227,-7856,1391,1082,2507,-9360,-1857,4621,-3215,-9311,-1309,761,-6108,120,-2604,-2064,-4020,-4794,-17773,-3459,-797,-3776,1861,-3403,1766,-4902,9990,-878,2479,-151,-5449,-1232,464,6171,675,-5903,6801,-4367,7290,-3701,-8261,-5825,6083,-2106,1777,-2727,1304,3916,3127,-5400,-6708,5249,-2724,-92,778,12324,-3564,-6103,-10361,-4892,-3940,-1065,2061,-4770,2156,-9023,2624,2204,-2396,-1202,-753,-7001,7915,-503,-1875,4790,3154,1801,-1816,-2880,-357,-9736,-2359,2052,-533,-1429,-1816,7246,-2995,-4455,1160,-6845,9760,-864,-460,6435,-1812,-4079,4460,617,-3920,-2885,-6206,-5073,1684,-248,-6362,-1962,5004,-1857,7065,-6186,-661,2082,-2907,-3293,-3813,15185,845,-2905,-2841,4204,-1400,4619};
    Wx[3]='{-1378,-2309,-282,2299,-298,-214,1143,-1861,-3410,-574,2142,3945,-971,-3937,5864,3054,-1604,2622,2875,842,2017,2160,1865,1461,-1249,-507,2336,-164,-841,-3747,-1455,242,1093,26,6474,2692,-655,-2164,1408,1848,3530,3967,-2656,2299,-6035,1715,184,1267,-22,-454,-8232,2966,3361,-1784,-633,2434,-583,4980,-4274,-3503,2331,3771,-2758,944,2758,1129,-3142,5898,-4025,429,-892,-741,2352,-1569,466,6523,2731,3815,-167,255,402,4348,-1184,2971,1939,4001,878,-2250,1079,7675,2631,1065,1727,-3020,3574,-3078,-4484,4213,-106,3627,-977,-11533,917,-199,-3879,919,-8740,-1040,-4504,-2614,3798,5678,5615,16455,265,7768,-10937,-8652,4731,1784,-1571,6074,-1126,5966,-429,-2094,2299,-6909,-11572,-2819,207,8466,-6728,2392,3859,6884,-3774,5258,9414,-9355,1990,-12490,-4589,7426,7246,-969,16123,-567,-1239,2091,-2093,-8925,5874,-3840,1618,1334,7709,-3981,3562,1700,-1507,15136,-4377,-1738,1712,-3020,4909,5429,4680,-1998,2575,-12119,-3278,2478,614,-10009,14658,-9428,-12324,6982,-4682,-344,-5795,-2330,819,9960,-5073,-1693,401,4995,-2392,-3208,-10673,-1693,244,693,-4008,4121,-4582,3312,687,8798,1505,3642,4589,1597,6000,181,-4316,467,-1317,-2719,-775,2868,4702,-1191,-9990,7128,617,2866,2081,-1832,-1967,2434,2714,4262,-1191,2905,-70,2261,5830,-4865,10878,403,1455,-3217,-3886,249,-5600,-2423,7465,2846,2054,12011,-7626,-6494,-6635,-885,-1210,2330,1209,-4750,6240,1488,3095,2639,-5209,3142,5112,792,-4550,4970,-3093,634,2978,-600,-4750,-3237,-1166,-2897,1100,2778,-850,391,1134,-1589,-2644,-3828,-7973,-2980,1318,-8920,-75,-6538,3288,-1279,7,6254,-1126,-411,-2946,3977,2563,-1843,-7255,6333,-8564,502,4045,-2570,989,11152,-2812,199,4062,-6044,10908,-512,-1544,215,1069,69,2286,555,4768,-10849,-389,3298,1457,3679,881,-722,4484,7626,2153,8413,3662,2683,4055,4438,1677,-654,13173,2078,3303,-5566,-2412,-1442,903,3842,6289,2648,-72,5888,-3652,-4721,3127,-3146,-6640,-219,1203,-3115,2379,-8500,8056,1806,-2761,-1246,7773,414,561,-2094,-3776,2238,5400,-3522,-7993,-428,-6718,1594,-5874,604,4692,1888,4423,4973,8798,-487,-5922,-1259,-351,-1043,6914,-4313,5400,-1370,4870,3085,-1842,4897,-4536,2425,-60,919,-3164,693,-6621,3945,7241,-10283};
    Wx[4]='{-2120,1262,-1751,-261,-1295,485,2841,-2780,-6284,2010,3139,-184,-10283,802,-1137,-526,-6420,-871,-979,-1685,283,-1663,358,-1470,-5834,-240,2242,-3981,-583,-2949,-144,-2261,-442,-3454,-9301,956,-3791,-1911,-1442,4643,57,1027,-7158,2902,-2575,-4560,-4985,2219,-4907,444,4348,-451,-1375,-1580,-892,-7788,859,-1555,-220,-3784,-2548,-2465,-758,-5336,-758,990,-2415,3879,-471,-889,-3083,3105,-4816,2653,-4172,-8715,337,1502,-3498,-6289,-2471,1137,-900,-3461,-28,-8354,460,-508,-3251,-1368,648,8701,515,2626,-2976,-2495,-3339,1925,-2067,-385,1574,5048,385,3757,-4018,-267,-7280,-5039,4467,4294,-3935,-2946,-858,4577,-21406,3498,-5439,1093,1303,-1646,2800,5532,3469,-613,-5239,-2152,-578,823,1278,3103,2391,19951,12841,-4777,-3305,6528,-5473,2297,-3918,-7158,-3688,-8398,-3833,-3344,-9331,2949,-5014,6850,-9658,-4838,-6196,-10839,3894,15087,-1883,-9208,-1602,-4160,5581,1441,-2257,9536,4421,12255,-2644,2954,4982,-17255,369,-3820,-6362,-3591,498,2836,-804,-9252,454,-4160,11484,-5229,-3164,1368,-1318,-5878,-7807,-409,159,-975,-4018,-2570,-14941,-4301,-5732,-3225,-1145,-8183,-1695,2641,2161,4665,-4921,8496,1102,-2985,2017,1074,-4084,-8027,712,396,-2939,1063,-6479,-6391,-3332,1160,13486,4567,-764,-1018,4960,-1652,-4833,2663,3911,-246,-24,2133,748,-398,484,-3125,1468,-9257,849,-3305,-2207,2856,-26,-279,-3425,5810,4621,9951,862,109,-9965,-4572,-3710,-403,-1494,-5634,-4584,2724,-2291,1324,-2004,4899,-3334,8276,-1549,-1044,-223,-11367,3020,1086,-2072,2736,995,1845,940,792,-5048,-7368,-4809,-3005,-8027,-256,1879,-47,-2122,4931,23,-164,-1016,278,-2260,-4858,1860,3347,-2722,2719,-4531,-958,-6513,-858,-9047,-3210,-8051,8857,-3657,4035,1549,1693,-1374,-922,-3452,-13193,-4104,-1779,-126,-5195,-13984,373,-411,3422,6499,207,1627,-4685,1172,-5283,-2731,3786,-1486,3366,1727,647,1159,640,2990,-6645,3317,-804,2082,-6035,-6850,2349,4848,518,2734,6279,1583,6083,191,-139,-10556,-3989,3637,431,9545,-2221,-6728,-8442,5405,-7568,-3491,-9067,3437,-1970,-1343,-450,-6962,-3940,4262,2978,-8164,10566,-1456,-11884,-3278,-1367,-3295,-1588,-3208,-10410,-708,-1604,-1754,-2836,-2695,9638,2010,-696,-6469,-5322,1120,-4228,-2744,-431,3315,-9755,-3637,6376,-2648,-324,-8842,-2800,-4729,6552};
    Wx[5]='{155,2254,368,-125,-80,-1270,3820,2248,3728,-449,4257,1976,1739,-1855,3935,-3686,-7739,9492,2644,2005,-153,1569,573,-713,2048,-1510,-3676,2230,2175,135,-793,943,2517,0,742,-1204,-2374,291,-367,-786,-354,2200,-1906,339,214,-183,-3432,-275,2961,-3801,-5019,802,-957,4282,1129,3461,3337,-991,1687,2536,2854,2073,6850,-3120,-190,-2651,-123,-2927,903,-561,-6767,4199,-3103,1376,-1268,-590,6088,877,-5336,2133,-30,-6660,2026,3212,-1882,3347,-30,-1730,44,-1605,-750,-4113,5224,-2946,-3823,-1096,4470,4968,1403,609,1684,14921,1478,-6494,3996,4631,-11328,-12714,3291,-3388,11250,1951,-3222,3913,6782,6518,6127,-5834,-3022,-2583,2207,5795,5488,9628,2067,4025,2482,2944,5390,646,-3952,17382,5986,1138,3469,4233,6171,2004,-8261,-6201,-1975,-3610,-17304,8486,3442,-7441,14873,2663,3530,-12021,11552,-13437,650,-10175,4614,-1190,8330,2415,-4377,101,-1479,-3718,4477,-5668,9350,922,2690,-8608,-570,-5112,-139,-12343,-3547,-10312,-1286,17128,-7539,-10126,-2102,-6328,3640,429,-7602,-1029,177,-10468,6030,5805,988,-5102,153,-4628,-4345,-1459,9189,-2124,-4084,8125,9443,6875,-3449,3986,-339,2340,-1699,-3437,-7099,-5380,-3210,5224,2136,2059,629,-10615,-5029,-7436,-8750,-2783,-1756,824,-827,1,3708,-7221,-1063,-2946,-4057,-244,-1145,-2221,-2294,-6010,-6938,-8256,-1331,-3576,-8520,-8715,2116,-6386,1397,-10312,1397,-7753,4919,-5625,5917,-2154,1916,-1881,-8110,6269,-2778,-2819,3222,-3596,-1741,-876,5429,1823,2617,-6240,-5083,2358,-4616,-6699,-1828,-1079,4038,1080,5151,-1613,-1571,2849,-1506,-951,4707,-8369,-2119,60,-2646,-4350,-127,-1131,-4140,-4819,-79,1057,-1354,-1596,-1992,-783,-4436,-2310,-3066,-7612,-4360,-3569,6884,-2430,-7050,5473,4965,1818,-2159,-5043,4384,-5698,-4074,5185,-4216,6743,-3034,-10947,-4902,-3205,-4929,-2175,-674,3637,-3132,-3879,1383,-3005,-3212,-1976,-1947,-1768,-1472,-1082,-913,-10185,-6650,-1499,1417,-1768,-5566,-3251,-3063,-4179,4904,-3461,-1470,-4133,6679,-2462,7646,-4023,-939,-5400,-1183,1331,-345,-5947,8022,5341,-3610,-3037,3442,1485,619,1318,-8779,390,-4104,-4016,1898,-10107,1475,5449,-3122,5556,-236,-2824,5102,-5371,-2281,-6088,3234,2318,-1575,1502,2695,7539,-104,-5019,3718,913,-655,1527,-3334,-6855,-5825,17861,-4079,-8432,2614,2714,3271,-3728};
    Wx[6]='{-1413,2678,3400,-1433,1183,2570,4470,4216,-1572,-1800,-1971,1004,-307,2934,1525,7988,1459,2305,3645,-3310,-3156,-2663,2312,-330,3869,11,1812,-1346,4763,1206,506,-1147,5957,1628,-3999,-284,1291,-2031,167,5502,548,-466,6455,919,6884,-2177,3703,1334,1989,1062,2185,1505,2829,535,-875,3935,-640,-5410,3869,-1784,-2369,-3908,704,-1066,4707,-2800,201,5502,1161,-2142,1047,2500,4501,311,-4489,-1826,4804,1489,698,6381,1369,1243,-4929,2329,2631,8491,-161,4025,-823,-4204,3044,-1796,-1244,2091,-4050,-884,2401,140,294,-4421,-1602,-3527,-3413,9282,-1024,-520,7832,5234,9960,-990,721,-4672,-7797,14755,-5166,-5375,-2281,-2685,-7749,-2805,-3356,6044,-631,2229,3525,6508,1273,3789,8002,-1594,-3449,14482,9370,1241,2172,7700,-914,340,-10048,-9282,677,-7011,-8764,13251,1677,4384,1389,-9663,-4755,3593,-6259,-5209,2187,6875,-561,8041,-718,3598,11904,128,3342,564,10957,1477,15351,-164,2333,-349,-1729,-5219,-8442,5717,-4865,3833,3012,10888,724,-19013,-5415,-2880,1263,7192,9970,-2236,-916,-2944,-3137,1966,3913,-3920,-1317,4543,63,568,1469,7187,6562,2142,-4477,1036,1005,2425,8637,430,4677,-795,-4733,1865,570,-846,7890,1085,-251,984,361,-2570,10839,-4382,3066,-1813,-2407,2011,343,-40,5473,-458,708,3728,-14208,-9433,-2186,9726,2766,3364,2005,2108,-892,-189,-466,-8173,-2668,8530,-5317,5996,10546,1523,-1689,-2353,-3232,1480,-787,4279,-157,-1291,5312,4045,620,1916,-1477,-3085,1141,9331,-87,2514,-2641,-121,-446,-2322,1351,-2333,-1676,-4589,451,5097,-371,8974,659,429,-2993,6928,6508,6557,-2551,1030,-897,6328,3964,-3046,1945,-997,-2080,2221,-1040,6279,-7138,320,-1374,8164,-2695,-3740,-2580,211,5263,172,5317,-184,-15068,-11113,-6313,1472,3310,-2766,-3803,-4697,3300,3432,-539,1881,-2958,-1442,-1644,-432,2607,-282,6171,676,1220,2308,-11103,-1807,-6284,-566,4914,510,4494,-2204,1854,2343,1420,-989,1188,-4133,4868,4313,-1330,71,-461,-6015,2120,-3002,4028,-4125,-1216,-444,12470,6826,-5502,-838,3476,-6821,-5351,-686,-3405,-113,5317,-2846,307,5961,-1562,-7446,-736,-9531,-5551,10078,3173,-217,-1606,-3884,-5258,6308,8793,7939,1733,8837,-1541,3481,2485,-2641,-3957,-6406,-2553,8339,-1165,14755,-10478,-2651,6035,6406,5961,-5327};
    Wx[7]='{-2200,5971,1126,56,462,266,6035,4860,3225,2675,-1798,-4223,3271,2678,507,-2067,1276,1165,-3298,8,-1811,2648,110,1350,-1173,-5214,1523,-1113,6269,-145,1372,7841,1260,-945,-2944,-1324,-3156,2739,2403,1420,3620,6406,-2980,2656,1862,-201,-10546,1702,-4328,-2573,5556,503,-3867,1372,-1170,2312,-1494,-6777,3808,-431,853,720,3520,2305,2355,-1209,1800,358,-2932,-4587,-3105,311,-3681,81,-1606,4816,5844,193,-3522,614,2387,-2812,667,-3950,-1231,902,-2081,21,379,-282,-363,3208,4719,-1402,6821,490,5136,10634,-3808,-242,-1693,5341,988,-1838,-1341,0,-6357,96,-5488,-4572,1320,3000,5839,7680,-12519,15136,9687,382,-303,-1611,4179,-5073,1051,-8447,1407,-962,2829,-2792,20488,-2376,-562,-5351,789,-292,5097,-4775,2770,4228,-4797,-874,4680,2883,-6884,-8759,-7197,4094,2094,-8583,20,-4951,-13134,2988,-1385,565,-4787,6333,-1676,2119,-16787,6225,6523,10058,-6899,2331,-7617,-2052,196,-797,-2548,-1061,7045,12910,1459,1215,-1016,4287,9536,-7329,-883,-1243,6850,6035,-9008,14169,-1843,-1240,4555,-2768,-2910,-309,-8447,-7460,3676,-962,489,-5004,2866,18974,2348,5346,3552,-12304,1318,6542,1761,2971,-28,-9541,387,-428,2646,1799,1717,7832,-12763,9072,-1934,1134,1074,-1953,-1878,1253,-1328,2369,-4714,-1867,-2846,2126,-1813,2558,2670,4023,-4887,-620,-2072,-4536,-836,-2211,1510,1944,-1334,-3225,9223,-4880,-508,4692,5507,258,4865,6069,3276,12314,-550,9536,823,-1938,4157,-5761,3867,4006,2113,-2259,1890,-1081,2320,-617,3691,-4365,1197,-5249,1645,1245,5180,1331,477,1306,-426,-4924,2583,-195,-2480,-1481,9296,5532,-5366,1102,2583,-235,2973,4274,3205,-2004,-5488,4626,-866,-2941,1530,5400,-4062,334,-1662,6650,2067,8828,-1290,-7290,-8354,-11132,2824,80,2690,6030,-554,3005,-5424,7641,-2275,9130,2583,-2912,-13525,4912,993,2290,-7924,-203,-2773,-243,2009,-7539,-2614,8090,-2227,1110,-237,-5034,-4624,1298,-3063,3051,1639,1574,3176,1746,681,8930,585,-1240,-1739,-1156,385,10195,-123,4541,853,297,-1582,-8432,5273,-2410,-4543,150,621,-175,8217,-2822,8828,-11972,5405,29,-2357,-121,828,3820,-9008,-1634,114,3208,-5903,2091,-1215,5170,9472,248,-11972,6796,5039,4416,4033,-3391,127,3046,-424,-2719,2426,-6357,4453,-47,3151,3654};
    Wx[8]='{512,1589,1065,1262,1115,-743,-2854,-4377,1734,164,-3076,739,-131,-1416,3159,2155,10156,1095,-161,1115,2103,-221,-2951,897,1058,-2152,4836,524,-5581,-1788,2893,-5156,-8178,-4033,-410,432,-201,2573,-1513,-4443,-1478,-3864,-2927,3083,-4699,817,10878,4541,-2993,-1497,6147,-6181,-92,3498,-1768,5229,646,1679,-3486,-2126,-2705,-3479,-1066,593,-760,1652,3618,-3034,520,1223,718,-9750,2132,1885,2479,-2807,-2849,1362,2025,2922,1133,4428,2380,-1512,2961,-4506,1864,837,1246,-281,4931,-6948,-3981,-4704,-7138,-1739,-1966,-2156,368,2476,-1523,-12792,1381,-4416,2072,-1270,1207,-5878,2531,-3015,1927,838,1846,6894,-15771,-11523,-6621,4172,-1489,650,1425,-2802,-2590,-4514,-2186,-5107,122,-1328,-11748,-5947,931,24160,2207,-4252,362,4121,2700,1431,3845,-5004,2340,-4472,-13105,-745,13623,-549,3957,-7485,-1098,5117,-1165,-9838,3774,-924,7260,8520,-9370,1060,1100,2839,1138,-4042,-5048,-4328,-6035,-442,-3137,-7929,-351,1252,-5732,-11796,-6391,-8154,3745,260,-7412,-8955,-9438,-1798,-2084,1887,1396,14228,6240,4499,3686,-2573,-1680,3881,2529,11367,-6225,-492,-12080,8339,4235,5288,-2727,-760,550,2915,2663,-482,249,734,5795,-102,-4353,1549,-3156,2147,-346,-1010,5371,321,751,6401,4899,842,1475,1445,2076,3762,1433,5214,733,1412,-1173,-1205,2507,1112,2055,-2824,-10156,-1228,1542,2558,-6689,-2851,-2271,-1199,-7529,2661,-5629,-5747,-8159,1750,-4887,-4694,-6997,6586,3815,-5239,-4106,-1723,-4228,5571,-795,-4682,1231,-1267,2761,-1323,-2580,2702,5053,-4072,-212,-1888,2028,3820,-743,-4331,2612,136,4440,3183,-2700,1702,2255,-1148,1470,-5366,-3881,99,-108,1850,-8271,1076,-5913,-145,-1967,616,-34,3732,6298,239,3625,-1459,-1300,2143,3034,2966,-1208,2205,4477,227,-5004,-2243,-4331,-2149,-6293,-3085,2873,-1491,-1514,3466,-2003,-849,-2656,1555,-2509,7431,3710,-2763,2253,6958,-2617,-547,1513,-1176,-6572,-983,5205,542,6523,1702,531,-4016,-2705,3562,-3117,-1652,-6655,-10966,-1034,3488,1781,-4335,2148,1340,693,-9291,270,-1230,-3684,2539,3125,-1677,3229,-3049,-2043,-5888,2487,3073,8510,1249,7416,-1949,1204,722,5634,2119,9697,161,7519,2961,-2465,-3432,7543,1385,3088,1373,1715,-4687,-511,2059,-5600,7480,1156,-9912,-2221,4733,-4484,7348,9360,-2597,7045,-1613};
    Wx[9]='{1690,2399,1552,-796,3037,759,6308,1051,6289,791,424,1627,3354,1691,-830,6474,-2092,-1599,2351,1685,-2026,1364,-1158,3222,-687,4741,905,1348,2424,45,3813,465,-728,256,2097,792,6787,598,-2457,-172,-351,-1011,1875,-1350,8735,2590,8579,412,855,331,2705,3276,1148,2427,320,-1724,-1826,5400,306,159,-1478,3649,-3522,5971,9248,-2430,-4179,-3105,-642,256,786,1958,657,6450,2758,-90,-334,-1019,4755,2171,2291,4860,6269,-182,3947,6103,2232,4829,3908,-2756,2153,7749,3249,-2670,-6865,-545,3796,-1386,1268,1752,-3256,1364,2467,-3811,-2932,-407,8759,1520,3933,8115,-3964,-3935,-1445,14375,-5112,-2294,3913,10009,-4169,4270,692,1481,5419,12158,-481,-8813,1362,764,-200,332,689,-4086,-10283,-16162,3808,-6728,-291,-6669,1910,-15771,3945,853,-7890,-6328,-2570,-3725,205,4675,-4475,3452,1486,9492,1556,-857,2315,13515,-7841,-5625,4389,2521,-2064,4689,17119,-1467,-2095,3093,7050,21953,-3229,-1520,-3906,8989,-4167,519,-3420,-3967,-10478,-12431,89,5014,-715,6103,9877,-5014,892,-73,-2283,4638,5161,473,5219,-1706,-4831,-1978,-5541,-2308,-123,-1634,-3608,-10449,403,1801,102,521,320,-1307,5732,-6650,-3557,-6215,2226,3186,-3562,8759,3410,-11298,-9033,3818,4787,1437,-1064,-2241,-182,-7016,-4069,1840,-411,-6,-3520,652,-501,5219,8134,645,1793,-98,-7216,3156,1907,-5336,3593,91,-10849,4992,9057,670,5366,4069,1883,-2092,-2180,7573,2194,-924,-5449,-7153,4460,1545,-668,-3156,2265,-3225,6127,3159,6020,-2423,361,7509,469,-1562,-3388,-5458,-1394,-300,-113,-2971,10009,2592,-505,4230,-1429,6992,-4265,-3281,-1478,-5737,-841,2612,-3020,-587,-2651,-2583,1122,1058,11132,-769,9809,-2597,879,3452,-4465,-3347,-6967,2413,1685,-7021,2181,-3828,3544,-3430,1978,4787,1442,3471,2624,-1684,-11435,-399,-542,2893,-8520,-1154,3041,-1889,-2161,2675,-3618,806,2163,5341,4841,5986,2083,780,-8149,-502,-1697,-2702,5068,-7211,-598,12910,-2008,7250,3579,-2493,7368,3847,3015,-4023,215,1822,545,5708,-7851,-6518,-3981,4174,-5102,1444,5517,1781,11074,-3378,6494,-3210,-6708,3366,9511,-532,-4960,1988,-528,852,-5473,-1284,12500,2385,1381,3947,2927,4897,-117,6040,3347,6635,1936,3571,1234,16884,-2683,-606,1782,3208,4497,-1173,4904,87,2756,5786};
    Wx[10]='{1484,4936,-1878,-189,1380,5444,-132,-1140,-2003,-319,-6005,-608,-670,6684,-3054,7548,7153,-5327,854,-2221,-3513,-4450,-1843,-3603,68,-2409,830,223,2061,1546,558,-4165,3295,-5483,1159,-2626,-1405,719,5400,1738,-122,1573,7128,-574,4953,-432,-9213,-612,-847,-1024,1235,-276,-323,-121,4831,4025,1481,-102,3723,3891,2536,168,3662,3012,-2929,-4113,269,-1525,2258,-1724,-673,1583,6425,3708,-1917,-1186,5024,4333,-1406,-1838,-1087,-398,-290,-5874,903,4291,3386,-517,-448,1855,627,3320,-2812,414,-5869,2044,4792,-1511,-502,-3090,-6440,12851,-682,5991,4553,-1195,-226,6816,9350,3256,9106,-12744,-6201,-8720,6000,3234,21562,473,-3623,46,-4099,-10517,-978,-6679,-2103,-403,-35,6333,-2829,-9575,4499,-5239,16044,-17041,-4841,-8041,2082,-149,2308,12460,1506,10576,7148,-15644,10273,-6982,1964,6728,1342,4763,14755,-3671,-1486,6713,-1096,-1368,-662,1676,-839,-2727,888,774,-19042,9379,-14619,2309,-68,-2531,-45,848,286,-2980,3129,11181,2951,5063,783,207,6552,-1582,11347,-1457,15703,-2127,3874,-6865,-3801,4008,5014,-873,-5673,1363,1965,5317,-12109,-5673,677,15751,9482,-17089,-997,-528,-1557,1218,-1370,-425,-4426,-5166,-2241,2180,1781,-3012,-925,798,-1341,3273,11591,-7861,872,-1113,-2012,-312,-2978,-3156,-2575,3005,-14296,-3232,-4572,-9975,-4853,2531,-4526,4970,-4013,-6948,-5092,-2951,-1384,-3764,-7578,3115,2609,-6748,-13867,-9213,-4877,-7392,-3730,4833,-5795,5825,-2937,-2504,3508,-6147,-1673,-2037,-7133,624,1905,1024,1337,-4194,-4094,-3347,-3159,-3112,2255,782,2048,7822,1096,2854,-1860,2088,6796,-1682,5463,6601,-6098,3811,3637,-279,-6630,1973,-314,-2514,-1045,-988,-10507,2753,-1069,-2177,-2741,-4592,-6713,160,-7490,137,-4792,2575,-218,-2041,-469,4353,-15078,-2443,-7446,-4235,-483,-1077,-1147,2199,-114,10234,5917,-6269,-5981,-8168,1318,-3012,-1564,-3796,-3593,4619,-5654,5087,-5214,-7104,-462,-2590,-1184,-3669,-509,-2976,3659,4860,-4130,-7192,-910,-5571,5224,-4694,-5034,-7919,-10654,-789,-530,957,-8369,2521,-4509,708,4104,1848,-2717,75,-5092,14736,-4326,-2526,-10976,-386,4694,-6181,6992,11425,-7460,-9541,4731,-4501,4680,-1771,-5776,388,10078,-3132,2866,10898,-5693,4860,-6264,2683,14238,4375,31,-1802,229,-1674,-4987,-903,167,5678,-9326,-4467,4577,-1669,-5825,-4819};
    Wx[11]='{4357,557,2822,1516,-1109,853,2675,-6962,-1116,-3830,-1463,-1154,5825,-831,806,7797,301,981,-470,3259,-370,-1463,-4040,906,-377,2374,1541,-882,2459,-177,883,480,4526,-2729,7426,872,2980,1082,4978,4350,72,618,-3698,1018,1590,3090,-3823,3483,7470,-903,4941,-2670,-2322,5659,-1246,6333,1527,-143,-2463,4697,-826,4487,-1345,3037,-3164,103,3330,-4023,-2956,-911,114,4592,-5688,2575,4111,4082,9194,-378,128,274,947,7236,365,-2824,1051,3811,-1489,105,3830,2202,-1787,-2203,-883,218,-1986,278,276,-5244,-2312,-1730,-34,-6918,1457,540,-4467,310,1920,-7827,4616,-104,6040,-1290,-2817,8247,3342,-7895,3684,8579,4199,3703,-3828,-3923,8022,-3723,-2291,3293,2946,-4541,1658,-4152,3601,-5,-2111,11035,378,4255,6015,-4030,14121,4475,2673,-3732,-1838,-2575,6987,4196,-6616,-5957,3828,4028,9184,-12861,-1071,-1361,2159,6918,-3715,-350,960,1257,-3806,-2218,2109,-2469,-3762,511,-6977,1506,-1334,1246,7705,12324,-1906,-10009,6020,-5805,-2475,-1125,-1693,-2443,-1057,-6416,7138,2978,2792,-9804,459,-7280,9472,-581,10107,7172,15419,-1649,-11611,-703,1915,-17880,4079,-4924,942,9843,2274,1329,896,433,4680,-6518,-5371,-279,-1927,1503,-4123,4699,8618,6704,3991,-4106,-900,1936,-470,-2839,-3615,149,905,-3735,972,-1394,-868,834,798,4284,1857,-3593,-1547,2211,-1868,-1855,-5366,-7836,2159,9208,-1419,1524,12773,118,6547,1738,-1876,2458,-5600,-8471,-431,1907,-5820,-6406,-2293,4494,2727,-9897,1319,1613,-2181,-6635,10742,-4716,6665,-13203,-2707,-3583,-3869,3969,-3,839,5263,278,2165,1997,-1849,-2060,2143,-1741,-3859,1083,6699,4152,1239,-4995,-857,-1163,6914,2011,-3249,-3452,9516,-376,4641,-554,5239,-1036,-2144,3769,4157,3115,5004,1080,718,-6044,-7280,-566,-1396,610,740,-737,6611,-875,-2839,437,-5913,3132,1994,449,-1060,1712,5375,-2773,-530,-7265,-359,-4838,2204,557,-4108,-4301,2301,6977,4414,278,1589,3029,-4453,712,1060,4924,10761,-4047,2104,3815,6059,885,-1907,-9345,1340,332,-12001,-3432,-7534,-2349,-4699,1427,3288,-301,-1,1486,5346,1047,4924,-2319,-5947,3210,-3774,-2812,-2546,283,1807,2188,6552,-3364,-186,-6396,8671,-9218,-10898,8876,10751,-148,-3825,-700,1044,3459,2023,-1007,-213,-3635,8818,4187,6948,704,5488,-560};
    Wx[12]='{1596,3435,3120,1920,-694,870,1702,-43,2150,-773,-2768,-1557,-293,1868,2934,11250,-467,-686,-1103,1023,-1882,-286,-2470,734,-598,-3518,1994,-1896,9,1778,-44,2656,6689,1749,-1066,2322,3310,9843,811,4941,2749,5131,95,5297,-1646,1229,4775,1506,2526,-756,351,888,-1519,1226,4365,358,-62,-2215,3039,1623,-4118,477,2359,-916,-248,-4687,515,1539,-1789,-5229,-1011,1739,2208,-939,979,194,1926,2980,-1783,-4475,-2578,-2055,8574,4858,-5585,6225,16,-305,-1783,4267,370,4123,-2095,-5185,3037,-34,5170,2595,-2656,938,4997,-17138,-3720,4465,-3764,1630,-3210,-14228,-5449,-2487,-560,-1590,-6113,8354,8911,6372,6923,4648,-707,-3200,1095,1600,8427,2770,-3876,8315,569,5449,-1837,642,6054,14755,-19677,14150,5239,-6396,-873,6748,-125,2067,-5869,10419,-8164,-4709,-1613,3129,-8984,-8559,3312,429,18564,-6894,-609,-2269,-2993,7885,-528,788,-2349,2692,-3017,1156,-2534,8315,2534,1201,1798,14638,-3107,-2402,5078,9262,9736,-1538,89,6625,9111,-2218,1932,3371,-2917,9345,6166,-8134,-1983,-20507,-3266,9023,4204,1717,1319,-3393,3125,637,-12675,-98,-4030,-9682,-5966,756,-4326,-4201,3188,4562,3190,-1352,-8740,-5737,-1104,-3356,1356,-1102,3735,6367,-7788,-4323,2299,-8017,99,-1556,1395,-153,-3759,-2668,-4035,-201,-1361,2109,9418,-568,1213,5073,-5659,-9560,-1055,1763,-2558,2485,1925,-5302,-3049,-3173,187,-287,378,6899,2998,855,2756,-2568,4545,6196,-614,4970,2214,-5229,4748,-3666,94,-4702,5937,-4213,1616,1402,-3515,-3005,-3059,1440,-1990,-941,-1373,7519,5068,2165,1276,598,4970,-7460,3435,5249,2924,5664,8740,1080,-2856,-9155,1138,-216,1094,1135,8364,11220,-4499,-4819,-5839,-1635,-2133,867,-2275,-6220,-410,-1600,6157,8076,5820,-3876,-3669,-1420,-6342,3269,-737,517,3483,2595,3510,2164,-6391,-1878,255,-5532,3015,3637,-3913,-4428,-3525,-1054,-386,-3718,4677,392,760,2032,2998,-5585,-7636,-1973,-3261,713,2626,-5166,-5537,5791,5864,12470,4631,7558,-3425,-2712,6440,-1408,1613,-2956,7924,3874,645,2321,2531,-10429,487,6958,1711,-5913,-88,1588,-1314,-4790,-3999,5917,-5410,-5590,473,7651,-1652,2491,-1522,7739,2570,135,1522,-3957,-2226,3747,1738,8774,-1752,3500,489,2153,1474,-1479,-2016,2413,-339,621,11191,-2631,-11328,-1295,-6933,-1114};
    Wx[13]='{-690,7216,2331,-437,683,-2758,2795,1540,503,960,5849,-396,2420,3854,-3522,1235,1663,3103,2910,1090,-1198,3093,-2536,2313,3063,1972,3100,3942,2320,-7060,-1040,-167,5185,2235,5478,3779,-12,825,-7563,2442,4606,4272,-2846,398,-2563,-648,-1239,3481,3183,-4550,3308,6181,-704,-2407,-3808,5234,1737,5917,5283,3217,-254,2827,-745,4111,-1469,-1989,4614,11699,4211,-1942,-4680,5175,-4501,38,-1762,2626,1180,3889,1801,6059,3479,1518,9072,-3203,331,2707,-2315,1497,1215,1378,1574,5683,1513,-3620,3476,7119,1994,1184,5830,8305,-5156,18837,1055,-2349,-6772,258,13603,-5122,7900,960,-3454,-4091,7412,17998,4851,2565,7700,-8461,1202,-1127,-1148,8159,-2939,9746,7993,5405,6474,-278,-5390,1324,-6547,4453,-29218,3254,7060,-1856,12070,2897,11855,-3999,7832,-13291,-12744,2492,-13847,5639,-9536,9555,-6865,746,14892,-11914,-1834,-25,6196,-582,6650,-1564,2871,5190,3471,6210,9633,348,2490,1564,-2890,-1934,-1470,-2249,-3698,-4645,-5805,2846,-10927,2083,5971,-2583,11591,-4104,7636,13369,-4116,8427,-4938,19501,4770,-3552,1372,1412,6254,-3217,-6806,-1783,8588,-555,13134,4970,4814,15566,2687,3676,1882,6186,-850,-794,3562,5913,451,-916,2941,120,-1640,-2338,4038,-5434,-1657,4641,3090,2288,-994,925,-2360,6650,486,-4204,-1588,1616,-2133,2517,3376,-4624,-5410,-119,-9462,-3928,-4628,-702,-931,-4873,648,-16396,-2583,4226,3796,-2739,-16113,-4272,-2105,3083,-2315,2614,1343,-2897,-685,-3469,-3715,2980,10087,-2023,3359,-5512,-5209,3586,-4746,-635,3088,-5991,4919,-2770,-512,-7192,1290,-566,-1799,-5292,-1110,96,4055,-4125,1530,4589,-49,1634,-4592,-1616,-827,131,330,246,8930,-9228,5849,-2480,-3083,1791,8598,-6889,5810,-689,3457,7470,6367,1785,-3955,4877,9848,1529,8876,-9052,-1914,3095,5502,2050,-6411,-2178,9023,-1899,7958,9111,-1391,-817,384,5751,-5673,3244,852,844,12197,7998,4523,3073,-6840,3754,2626,-7612,1015,3583,296,-1903,4892,3144,2414,-1865,676,-270,7700,-3730,4716,-84,7797,2539,3564,-1370,-2355,4316,3200,11718,8183,10654,-407,2492,-2631,5107,-7016,-5390,10322,-5405,13164,14628,-2517,4680,3142,-944,-9472,5615,5908,5249,-4291,5463,8017,7246,6621,-363,2454,-1061,-3952,366,3054,8281,1717,-15234,493,-710,-10058,3623,7250,2890,3977,8891};
    Wx[14]='{3645,8798,1480,-1552,2460,914,5844,614,1738,-974,5673,301,-6533,-2303,-7783,486,-7075,2722,-467,2580,-4311,-3745,-364,1625,1246,-1855,1431,-3063,5791,-2092,-946,-1861,-3847,-594,2458,-2866,403,-2099,3930,-2070,-2269,5312,-2156,-3120,6977,-2619,-5107,-4394,-1708,-566,-4682,1485,-963,-2442,945,88,1041,4145,-1473,-762,2500,-5268,-6459,-1491,-853,864,-821,657,459,303,3518,-4558,1056,-1677,-1104,-3527,-5551,-2398,-5654,4660,-1566,-481,-1508,1091,726,-862,-2196,2597,-5214,-2099,-2597,5068,-3757,2719,2626,-5078,-2548,1293,971,-1164,1439,1871,-1008,-4897,-2077,-1182,7968,4963,-1240,-4396,4519,7670,-2961,391,9550,423,6782,-3203,-3024,5473,28,-1296,-693,2421,1347,-3017,389,2890,9086,6401,6503,2404,5175,-891,-3666,-3388,516,-4440,10966,671,-11416,4555,7958,-5996,-1289,-4716,1778,3786,6015,-194,-4333,-2415,1820,-6142,-3518,-5688,8994,293,-2851,-502,-3874,-3549,6733,-3762,6791,62,313,4594,-1629,501,881,-1507,-578,6503,-933,-2486,-3937,-6303,-3615,-2388,2998,-8378,2165,640,5566,-9243,188,3989,895,-2666,5937,7216,2963,1694,305,1826,1357,-5415,3105,6059,2445,761,2047,993,211,-1844,-1848,-1693,-2929,-2322,-2220,97,2966,5449,-5791,4243,11337,3305,-1300,2054,-2429,-3903,2810,-2011,-564,-1207,315,-3872,1111,-2216,-3825,9189,2858,-352,1627,1644,697,-4125,2280,4877,-1182,-1884,9091,-4494,1998,1490,4157,1945,5463,5468,11201,1112,-1040,6674,-3703,5444,5981,4152,-2187,-16,-3247,7958,-1411,-1491,-1605,-4240,-314,11142,870,2023,963,-133,6977,5698,1046,1690,-25,154,-5971,1883,-542,3557,5249,-3225,2563,-962,1943,-956,646,2392,-9379,4638,2998,6411,3996,168,-1442,-4499,-1999,6557,1185,-198,1115,-505,-1091,4753,-703,9326,-3996,-6533,3081,-691,204,846,-3308,49,1719,2200,-9677,731,-3354,-3862,-596,-107,1116,2514,-690,-6523,4213,-4287,-6601,-856,320,-4489,6083,-4094,-509,-7705,2320,-2648,-1407,2788,3603,-7749,-4116,-4592,1728,-6376,936,2167,-1381,-434,-1475,138,-6601,6376,3095,-1341,-1081,-523,-3974,-733,-6796,-8764,1839,4614,-2758,13681,7573,-4577,5786,2316,-1726,871,-8520,-7939,-4514,-6274,-5581,5410,-925,-5727,6938,-1391,4040,533,4453,6225,-2260,-1500,-8627,-9008,4733,4274,2186,-5776,-4172,-756,250,1243};
    Wx[15]='{-397,-9116,685,-3522,-3063,-651,-5478,-880,3334,653,-3054,-3203,191,543,-1318,-3745,-1540,-4470,1523,974,1870,-4096,-3876,-547,-2189,-2849,1014,-1437,-1870,-4362,2294,3676,-6621,-5698,273,-2305,1039,-5229,2399,-2714,-2437,-1379,2060,-3066,-4196,676,1319,-2316,1480,625,-2054,-6440,802,6279,-1162,-11103,1309,1301,-423,-6440,-737,-346,-6733,674,-1113,1434,-303,6,-4062,-4460,1799,-3559,1434,-1390,1235,610,-2685,119,-2104,-4284,1829,254,-2819,-4140,-5483,-3420,1906,-2355,484,250,1787,-3444,825,-2099,1265,-874,-5556,-2438,-3879,-1881,3562,-11904,-2397,7539,4450,-1699,567,1633,-7465,884,14228,1779,6333,-516,2452,-1778,1961,-6474,-2734,-487,-1203,-1317,8339,-5781,-2912,-2276,-2196,1297,-8447,-1235,3103,-7006,-5493,-5405,-6811,1533,-548,-2995,11757,697,2717,-2384,2526,14833,1160,-10742,-7055,-5649,-1672,4548,-14863,127,-571,-14677,-737,7641,2954,-782,4465,-1743,-120,16162,2145,-395,-5981,-92,1884,-7387,2490,1115,9208,471,3427,4565,3708,12363,7744,-3129,-16718,-3237,2839,9199,-6352,656,4331,-8881,2434,-4692,2753,83,-5361,15117,4121,1929,-7861,-7089,-2116,9228,-3991,-3532,-1701,-4689,-2148,629,2780,1140,7246,420,-4797,503,-3823,-1312,-2714,-1146,4863,5024,1842,-1774,2408,-510,2832,-277,-2514,1875,3874,-2052,-667,494,319,5776,-1206,2561,5766,-974,-3676,-3642,60,-2866,-5302,-4670,-597,3459,-3583,-953,-1802,-4113,833,-2832,4743,-1358,-4169,-4416,1022,-7465,-1674,5888,3537,-3886,-6069,1997,-3017,-856,-3342,-1057,-8701,-1650,-3083,10156,-2768,-2995,-3574,5312,4135,-1809,2805,2490,-7055,-3151,1120,-1270,3491,-10195,5468,10146,620,1848,-1358,-3813,-320,130,-2144,4604,-4807,212,1680,3063,922,4453,-3056,-1306,3918,-6694,-7895,-5058,-197,-6113,717,637,-4189,5678,207,-1638,-5620,-3964,-4118,850,-2766,1127,4658,-1400,-12363,2432,993,-1242,6240,-705,-971,-6806,-5625,997,-3869,704,-369,-10263,-3181,-455,1590,-2995,-6933,-3276,-2498,-119,705,2568,-2612,-6044,4160,7441,52,1390,-7558,-4897,2154,4870,-8935,-12333,-1538,3813,1888,-5214,1502,-2073,2462,-10507,-665,2717,-1629,-1307,-5009,-4184,3537,2470,374,-4875,1801,-1998,-7192,2199,-3068,-5541,8569,-4514,-942,6552,-14521,-4482,-1289,-3046,-3032,2291,2963,6611,-4885,-2961,-1746,548,2863,-1231,5034,-3935};
    Wx[16]='{736,2915,-1203,137,-946,-639,1292,-2744,-1357,-106,1485,1206,2800,-462,7426,-301,-4072,1011,-2357,-1416,2871,-1794,3891,3063,-1062,-144,3774,1219,1078,3715,-1789,-2495,2614,2797,936,-5913,-1336,950,3085,2985,1621,509,-957,3237,10039,-869,14951,3117,-1122,-72,4470,2553,2946,2949,-4155,310,3168,3769,-81,-663,-371,-1016,3923,-603,5615,2181,-320,1524,-2998,3710,1431,4907,-3754,1335,-627,-173,4765,3884,2690,-6,706,-188,3967,4538,4458,4645,-1578,2561,-993,-210,1350,-1181,1518,1910,1918,-2514,488,1705,-1156,2416,-1998,-6684,-2639,-1411,-262,194,-4121,9492,638,-5957,-548,3239,2995,2770,-154,4453,-9458,90,9091,-3730,4768,-5297,1750,-7128,-933,3090,-2218,-9550,-756,7534,-4309,11962,3588,216,5117,-594,-464,-3120,21328,-10468,-3723,5917,3830,-2380,5541,16757,-4367,3327,3022,-3452,-4016,10976,2331,622,2338,-155,-1408,803,-516,-368,971,11562,544,-7568,-2244,-1988,440,-5083,1917,-1571,-6826,-5126,3803,-2197,-1052,-17187,-3911,15839,1450,342,-5434,-1922,-1120,7700,5273,-6997,4189,-7172,2658,725,4724,-9023,-9555,1187,5527,3740,-12177,11474,-1348,4130,1909,-218,-2027,-2521,-116,58,-5776,1364,-17,-1201,-31,-3063,3913,1972,-10078,-1726,-1827,637,-4931,809,-823,1744,-1339,2387,2790,3522,2709,-1484,-1453,-3591,283,-3247,-3303,2103,714,-9,-1287,3554,405,-4648,3605,362,-4919,4201,-2198,-1690,1409,-1748,-930,-1757,-2973,-2246,36,-7,-5253,-2529,-6997,2714,-3713,-1865,-4023,-8793,-4436,2578,-3083,1569,-3894,-12500,-3039,-1282,-4384,-1243,3930,-4545,-2524,-13701,-3986,228,6210,-1898,-1018,-5776,2187,-4770,1141,-8432,-1925,151,991,921,-960,-1470,1995,955,2095,-421,-2275,-4521,-751,-233,5800,-882,-6020,681,726,46,538,-1308,-1237,1490,2832,-3669,-196,2075,-5502,-6728,-2529,6875,-4243,2668,5405,3635,-2,2556,6704,125,7055,1475,6171,-3486,1048,-2320,-3032,6601,3686,-3144,-592,-1818,1806,25,3430,4211,-955,-839,-4284,-2663,2626,900,-160,612,3312,-5776,3327,1188,1623,5654,2839,-6240,1981,-1209,-3383,-5434,-4370,6318,1970,7934,-1466,-10927,2114,3181,-289,2714,5507,-2385,-2861,-9140,5170,-1398,1462,-7226,-958,-12636,1832,-5478,4753,-1409,-6489,2866,-1400,-3044,1960,2241,3613,-2138,5126,486,4777,-7597,1490,-1084};
    Wx[17]='{-1833,-3581,869,519,-225,2176,-750,-6733,-1621,2897,-8520,2563,-3054,-2622,-3361,-653,-6054,1139,-1221,2044,603,-4741,-2888,-483,223,-4167,-3928,-1605,-2958,-3645,-2105,-3696,-4995,-5317,-6933,2242,-1524,573,-6489,-472,-1341,-2578,91,1184,1062,-3244,-12451,3952,-2103,2280,-5458,-15693,-4421,-6152,-5073,-8662,-1843,-515,-2980,-5146,-4958,3220,-627,-3012,-7685,512,-1353,2705,3920,-1877,-3708,-416,796,-1015,-847,-538,1127,-3439,-3854,-454,3281,157,-775,-4194,-274,-3293,628,1380,-2924,-3559,339,-6992,-2995,464,-6127,-8818,275,-5468,-527,-7104,839,-2277,-801,932,-1480,-1580,-2337,225,4277,-7719,-4541,4501,-4204,5112,794,1420,-2644,5864,-2714,157,-1286,-3696,2387,713,-4782,-4382,7758,5795,-6464,-4916,2673,3498,2427,7646,-2802,3352,-1129,4680,-9760,-6132,-5463,-5209,6357,3972,-1224,-15537,769,450,-44,6699,2697,-12509,-267,9194,-1296,-2729,1352,-285,-3305,-445,-6459,-2795,-6259,-1645,-9257,-3264,-1380,-6,-990,-2990,-7934,-2736,729,-10966,-564,-1550,15166,3110,-5151,-3100,2509,-7001,-486,-720,410,4311,-6845,11572,2479,-6152,-9599,8862,-480,115,-4296,-7861,3366,-409,1242,-2238,-413,12402,611,1182,758,2827,2775,-4697,4716,2277,-732,63,-353,-2885,12910,6865,-1911,35,3715,1730,687,-629,-3845,-3779,-447,2462,-1813,-1419,3315,7050,-893,8608,-365,5512,-1027,-1665,3466,204,353,7407,5839,15371,-10644,1553,-5874,10761,812,-4665,-609,3686,2905,7324,1912,3332,-1188,7177,5913,833,2858,-3391,-4089,4382,5131,-5034,4748,3281,3952,-5024,1927,549,1574,6069,-2412,3259,3410,1674,6259,3823,3154,3388,1239,-4667,4863,-1541,3513,-3774,492,5092,-686,1281,-54,7954,-6918,-2302,7426,-3630,5556,-382,-2272,2626,-507,11650,4370,-343,-1872,2479,4099,-8613,-3378,1306,-2452,-641,-4255,-3603,7099,2015,-550,-932,5244,1629,-2121,-3051,-4733,1116,115,-1597,-3232,-34,-3085,1569,-3176,778,3535,3405,-7670,3601,-3962,-1593,-1097,1505,5039,4924,-3967,2148,-2287,1486,-4165,884,-4963,144,-572,-5175,-9462,-4897,4951,-2154,3569,-3061,-101,-1981,-762,3256,1262,-4243,1763,3198,5512,807,4335,-3840,-1511,9477,-861,5126,4050,5126,4470,-1146,-6958,32,875,-488,1846,9257,5966,994,-2983,8876,-3957,2429,-5625,3027,-4926,2673,11816,-5302,7456,-1334,-972,2670};
    Wx[18]='{783,1519,-754,873,133,1511,3508,-1226,-687,296,-3156,-753,7260,1734,1590,6166,-1072,-2519,-504,1973,-3637,-271,-981,143,1170,2026,136,639,-3837,3623,-2749,-9008,-4487,-563,1164,2475,-1555,243,2402,-1978,1076,-3154,-297,-292,-5463,2954,-617,-1159,-1903,-251,2030,-6103,333,-1086,1701,1993,47,-3083,1785,4992,-272,-3547,-931,3503,-316,1262,-283,1059,1285,265,-1992,2392,-5629,-3681,2352,-234,1318,3308,1926,-3615,1604,-1505,1697,6928,-1977,-1639,19,1224,-1501,1945,514,4162,-341,3410,-4172,3020,13,-2425,-1926,-2551,-4121,1857,783,-5727,2917,2795,3249,-3508,-727,-135,7465,-5180,-366,-2741,-605,-3615,-82,-3127,-6298,5283,1053,-1436,-4394,2502,-3044,5312,1501,-3442,632,-3781,864,6689,-4567,-7998,83,-895,2352,4018,1216,-4772,2590,-2504,6547,-9682,-2546,-4006,12617,5004,-73,2486,8740,334,1414,10419,-4848,169,-1513,1473,-1824,-1497,-3974,9028,-8081,6953,-8203,-1798,-7578,-3786,-2810,-1215,-3125,6005,-2442,-1037,3505,-6450,10625,-598,6469,-36,-2021,-2863,-5976,10117,2534,-5864,1289,3374,3034,-3103,-2258,-10341,205,2980,-69,-896,-1816,-9711,-1347,-806,-4143,-7285,1436,3193,2478,1480,-3029,3903,3024,-112,8608,-1883,2900,-2150,-1422,-1929,-2534,-470,-1075,3415,-628,-531,3728,989,471,1115,3347,-2116,-1567,-133,-111,9462,3447,4182,3454,-1448,-1889,1211,-902,915,-2452,-710,8071,3798,-2888,-3208,-4741,-1054,455,-2470,-3906,3508,-337,-4687,-2039,-2208,-2048,3684,-1380,-9394,-1885,-1223,701,-3356,8173,860,-1323,-9370,467,2352,-4553,-1063,1469,241,2385,4455,-1550,5625,3935,-3063,1142,6635,1926,2127,4831,2037,2360,-1948,-1939,4343,-3159,5410,5400,679,-2651,-3461,-6015,897,-2313,3103,-894,-1716,-3674,1823,3867,-2170,-348,-4609,-851,4848,3427,-1345,5712,2687,1173,622,-2254,1317,6513,-3420,-2910,-1549,299,749,-2512,2021,1452,-602,-5678,-650,-5830,2780,-2722,-341,208,-2590,2131,-2297,4548,4050,-2043,-1088,568,-3618,-2147,-3928,-6958,-3835,3601,-1829,-6757,596,7241,-7573,-2100,-466,-3269,-692,-2739,-6025,-3537,-2263,-5156,5180,1654,8813,6049,-6269,-14736,4252,3391,-1751,3903,281,905,-3579,-2695,2486,1222,-141,-1807,673,2521,-551,7104,3476,1604,165,225,-6313,-1926,-2304,2463,3857,-5029,-3286,-326,-4770,-181,-2401};
    Wx[19]='{200,-3798,1516,458,-2873,-1663,4665,1318,-353,-3630,-1562,306,-3505,-4011,-861,2868,1516,211,-791,292,957,127,1074,-582,1395,2592,2327,3029,1273,733,1130,-3430,5561,2595,-4111,1278,177,-1202,1036,1152,-1170,1582,833,-3571,-1673,-2236,-1837,880,-1021,-2314,-1490,5263,1934,7968,4194,739,21,2973,265,2097,2680,2239,-5092,-2110,887,-1889,389,1933,-1860,-1392,-4387,-488,-3557,-1155,-869,1029,3061,-1757,-2590,-858,-2023,-8154,-1837,-1550,-3085,-3088,133,107,388,-2272,-6552,6000,-1408,-1553,540,-458,-3173,-40,5566,-4370,2176,-1356,-57,12978,-2939,1397,3845,473,153,-220,9199,1795,6459,10869,-5595,5751,-4460,-2070,467,2573,1285,6206,-6489,13437,1651,-9995,-2167,808,2320,-8081,6093,592,-994,-4033,-2486,-275,-1019,-9301,-5932,13740,4975,-7412,-1414,15234,11152,-632,-4924,5224,-22968,716,10419,8139,9150,-9438,-1094,-4006,5048,-2463,-356,1342,8017,-161,-6132,8666,15380,1173,-811,-2697,2580,-3232,-3395,-3854,-4482,-12880,1124,-3508,-3652,-2900,-13662,-7500,5375,11962,3635,-1845,3168,-6508,957,3840,-2963,-1468,3662,-7192,-4758,-355,-1925,9140,4736,3571,10654,-24199,-2568,16152,-2465,3818,-1467,-23,2229,4128,-460,143,-1798,-642,-3295,2695,-2631,4145,9165,-3762,160,2338,1472,-1050,-1557,-5327,-3847,-1232,-3598,-2680,-8725,5771,-1311,-6298,-850,-1523,1721,-1508,-1343,-3259,-1109,3542,-545,2768,12197,-3784,-5522,-1035,4943,894,3002,-513,-375,-947,8022,6835,3583,8500,3063,-2490,250,162,185,-5400,-3930,-5190,-1127,52,2312,6289,878,-1395,1855,-5517,-4140,5473,-3139,-5224,7075,-1403,5263,725,1102,-1881,-676,-936,769,3969,528,-1877,6318,2490,-6347,-2763,-3674,1887,-2653,-2600,-5629,-13925,591,-1490,-1590,9047,-6665,-3854,-6582,-18505,-4914,8422,5947,8173,-439,1439,6005,-1794,-1733,3610,8798,-1977,-4379,1687,-12392,-5493,-3039,872,-2358,3432,4260,-5004,7124,8715,4460,2276,-1810,-4477,4418,278,172,-3100,-1651,-4162,2812,2238,1049,4772,3059,1585,-5668,-891,-9121,-567,9077,-2100,1856,-994,-5961,188,3144,-5097,3061,6230,2435,7421,97,-2502,-1152,-14062,-2634,-1921,2130,-6640,1674,-1607,-7832,2670,-3825,-1222,5126,-1353,5087,7631,5380,-2150,483,1968,477,3583,-92,-3315,2167,585,-8017,1682,-1915,10234,1628,4785,-1846,3388,7836,-2670};
    Wx[20]='{531,-6928,-305,-2481,3520,1820,-526,7148,1315,35,1309,-2758,-1826,-2456,1812,0,-1599,2858,3134,-218,2490,4448,-2082,57,-1734,-1541,1307,2015,4130,-3859,256,5698,928,-2441,2368,2196,3369,1624,932,-1270,1142,-1367,1036,-1439,-2448,3557,-8564,-4560,4934,145,4577,1804,597,-2155,-3247,-5351,-1887,-2133,-686,1378,3,5649,-5698,498,8813,-3395,1348,2437,3208,1414,6572,-4372,-3437,-4909,1904,-40,-1020,409,5288,3225,-371,-5571,1782,-4570,-1403,-3295,122,-761,1577,-1529,797,-6025,-395,2086,936,3903,-4453,2514,-458,-211,-155,2602,1326,-3613,13564,-1744,-3610,3793,-2805,8120,-9833,-3774,1821,1352,-8974,-5625,-2034,546,5170,-433,5327,303,3259,2902,7412,-10439,2333,-1383,-3542,4526,-533,9589,-5585,-3964,3093,2690,2401,400,7529,-4475,-1113,-15957,9379,9731,9257,2493,6333,-10341,1190,5742,-1285,-12617,8041,-8403,8447,1453,4326,5239,3300,-1256,6577,7226,306,3840,-3071,-3234,-2604,8588,1063,-2318,2551,-3425,-2139,22343,155,-1911,-15146,7026,-6088,4489,-3190,5976,-872,10175,-10253,4790,1129,4548,7,322,8686,637,1362,903,-2893,2575,-5966,4404,5419,-15468,-1547,-6479,2287,4204,7866,2082,6181,-7695,-4260,591,-2041,1918,2435,-1398,11582,-4738,-736,511,1335,-5278,472,-997,6708,2060,1004,2607,-3322,4323,4416,5922,-1246,-243,-2863,-1257,-545,1923,-4658,-1552,-2495,678,6064,-6650,-8994,3183,26738,-2524,-9418,4848,-1141,3554,1291,4255,3076,-6318,1788,3142,4819,-217,-807,3398,-1270,7060,4597,-5810,-6821,-2304,1291,-1903,-1636,-2888,4509,4738,3300,-1674,3715,-1364,-2315,-2995,210,5708,836,-9956,2478,2939,-5439,7128,1517,-3281,5087,-1148,1271,306,-255,1097,-2382,1179,1530,-4968,2279,-3381,-3000,3825,181,4040,6010,5229,9316,-1965,-2778,1021,-1270,5200,-1136,5742,2014,-2580,-4982,2556,133,1624,-302,384,4428,1881,1180,-2429,-2666,3793,7836,3540,-3261,2030,-3176,-2059,-1679,1768,-3522,-29,-8168,22,4548,-5014,1740,7363,13085,-622,-2792,2336,8945,-913,5952,-1121,3395,-4072,5141,-1486,3559,1182,-1861,-2773,2308,9404,2648,4790,3020,-789,2424,4855,14248,11826,1864,6176,3757,-780,1754,4450,4624,4,-1115,7470,6650,-3122,2443,9160,-8583,5449,2822,1683,-1815,12880,58,2003,-1575,16083,5288,3322,-3317,6640,1873,3105};
    Wx[21]='{467,-5493,486,-1389,25,536,-3127,-2384,397,-3715,3564,1763,667,993,-7963,-4865,6816,3107,3027,1428,3298,-3933,-2717,-1317,1790,-1167,3439,1943,-4160,-2731,649,-2344,3178,1243,-2243,-1193,-308,-443,2426,5092,-546,-654,-3269,-4099,-7504,1162,2050,6772,827,2685,-1096,-1541,3977,415,2744,4357,-1851,4399,341,2919,-541,4223,-4624,4460,-8305,460,3059,1268,280,2954,2025,-1034,729,1551,-224,-656,3000,292,2346,-1966,50,-23,-4672,-7485,142,1881,3269,-3225,-1588,98,2795,2226,-2402,-1024,89,-170,-670,3471,299,1325,2802,7260,3261,4821,9946,-2010,-2854,11582,-1385,3376,-7690,-309,2653,-8037,6533,819,-3635,-5375,-987,-3364,2766,-8056,-207,-3784,-985,54,337,-2452,-15419,-3115,2968,15312,20781,-6406,-3566,2854,402,3159,-810,-2175,-4760,15703,-6313,-14589,-10742,-6181,-14648,11318,-398,3215,2807,10917,2193,-5732,2939,-9194,-3212,1824,6464,-2912,4372,35,1467,-4436,4521,256,-5429,-7607,450,-791,9204,-11816,-3078,2257,-2785,6000,-7841,12695,1733,-7177,2250,3508,-6796,-164,-8168,12958,362,-5507,3593,7788,6611,3159,-7622,-3498,-180,-2403,8295,-1013,10703,-14033,-1184,13222,647,2308,100,772,66,9326,-4819,2136,1580,4338,930,-11464,4116,2565,10371,7031,2193,-2158,4445,1624,5244,-4472,5478,1183,-6948,1499,5566,5488,-6479,4873,-4423,5839,-3701,-4516,203,-2827,5268,3300,-2702,6425,6821,-12744,9287,4477,-4260,-2912,-1929,3969,3811,3725,-2209,8593,8671,-941,6054,-96,3002,4838,-3242,-6113,5410,2961,6284,-848,6069,16826,-163,1623,492,7324,-10,8930,108,1468,6464,-345,-3464,304,3259,2335,2252,-869,474,-254,-556,2341,3178,1567,-3483,3767,3732,567,-449,1054,3952,2341,3808,2966,-1906,8842,35,-2797,-3083,9560,-3239,9873,1956,-253,1201,2944,-6000,-1320,-4367,-1026,3034,-2565,3876,-7343,7753,1485,-1848,-1665,-4494,4946,245,323,7880,-1586,5981,4807,-3884,475,-336,4345,6821,-1508,-1778,3447,-214,4284,388,-7885,-948,5107,5263,4753,-4238,3229,9433,7138,-6787,433,1157,-7441,7075,1373,-4116,1250,3393,6689,435,-4108,-2023,-872,6372,8261,-15546,-4985,-955,12431,2866,7495,5693,2298,-7197,-3251,1395,-4187,-2493,-3845,2010,17861,-1257,7265,-3747,6586,4086,3759,-635,1605,-1172,-1002,-4477,7763,7255,9233,-122,1674};
    Wx[22]='{-3217,-5507,670,83,-6831,-2100,2285,845,-1473,-1005,-1380,304,1271,-467,751,-1950,6542,-549,1717,589,215,1189,920,3764,-2543,2858,-2386,2103,8237,-3842,1379,4741,6674,5151,-3327,-3178,-117,-1644,1359,-1094,1026,-8330,3962,-1383,415,-3461,407,-4367,1258,1640,-7749,-3557,5585,-3750,498,-4238,241,3459,-2041,-164,1017,6445,-1545,-826,-4770,295,1607,-1036,-2534,-1009,-2298,-1307,4409,-3139,1945,1745,4831,5415,1282,-2614,3701,4907,-1666,-1533,-1971,3598,343,-1207,-3005,5000,1871,-3098,1859,-445,-842,-853,-3891,1348,5253,841,-4211,-11201,-3044,-2756,977,-436,8510,-2797,18,3239,-5327,4624,7602,629,16689,-1229,-437,-11132,8491,1259,691,6811,1627,-1795,-164,973,-11,-997,4260,10898,797,2386,8291,3398,4191,300,-1821,-2802,8510,-9301,-1608,-6782,-409,10107,1839,2998,299,11357,449,-1414,-3996,4863,10273,-2285,526,5332,12109,-6342,11181,2279,-3745,10419,4169,-3852,5825,-1082,360,-19550,1911,-2098,10048,-2266,3889,2880,-3410,874,11826,3857,-9179,-9526,-4638,-6933,4291,8945,3864,-367,6157,2366,-2407,-523,10605,-2155,-7211,-3100,4045,-525,-11513,9531,-2116,-4699,971,5771,-1893,2073,-7285,-1501,-3486,1143,843,-1778,-2430,3073,-2099,-3056,4211,-4260,-10742,3103,-3254,4326,2172,-1164,-6210,2580,4450,-2687,4812,-3376,-1492,2026,328,-17207,4372,-6772,4104,4929,-2296,-3435,-2475,-3796,5327,-7050,4711,-3269,10810,-4948,2303,707,-1766,4025,-11132,-121,1765,-4086,4643,2326,-487,245,1436,-892,1936,-2509,-6411,5322,-7421,683,806,-16689,-392,-3137,6308,-3527,1721,5107,-681,-1696,-4277,-10693,1597,-5068,-82,-6630,9282,-4787,1649,-3349,-310,105,5874,-2020,2983,-2993,5981,-690,8964,1435,-3623,-6474,-805,2000,-808,-4113,3261,-9350,-6943,-6147,2015,3959,3073,-4377,2136,-1055,1394,-9814,-7539,-4299,-2039,5512,4160,8564,-10302,-1154,-571,3537,3007,3479,2927,-6694,7500,11728,1751,-6596,3576,-5458,-1489,1715,-2022,-10820,-6484,-1596,2770,-7504,1948,-4340,7846,-8193,-1285,2244,-10302,7153,657,-4379,2519,-7475,3381,1652,4260,10234,1241,2661,1483,1956,790,4233,-6083,-2619,-7490,-10810,-11894,-6005,5874,-4274,-7221,1906,-4257,-100,-1596,-453,4228,-5014,2600,-9833,9506,-4538,-8354,-6718,-751,-1618,-5351,7856,8422,76,2819,-7592,301,5239,-1936,-2846,-4775,-4108};
    Wx[23]='{-684,5375,-1573,-1748,3486,-496,1864,12,-39,-205,5102,-779,1285,-3767,749,6015,2125,552,1271,161,-5444,983,-1196,-1170,-708,1341,-142,-2673,53,8056,-1313,8178,64,-910,-3671,-447,1704,405,1802,3786,-318,4001,202,-844,5688,2604,6875,5483,4169,3166,2778,6811,-1141,132,2296,4531,-7685,-4902,3027,5727,-5200,-284,3251,-333,8930,74,-1004,4228,646,-1375,-1068,5439,3630,-812,3054,-229,966,-599,3703,-444,1882,4458,-5566,13701,760,897,2856,-3508,1110,-927,6430,-755,-152,2575,2476,2008,3005,379,259,5502,5058,-5224,1511,-8969,-1469,657,5009,-10507,-2827,134,-9672,-6284,-8081,-5415,-7021,-7148,18671,1918,254,636,-2912,1051,-975,-5541,2695,-3107,1542,1585,4636,2531,4060,-1324,-2543,-10117,-463,2409,-774,-172,9526,-4140,-6484,18623,655,-2734,-3540,12939,-4689,-7402,3671,3054,-11630,-13027,3242,13496,-2052,-3850,-12880,765,-2076,-4367,-4487,-12333,-11738,-4741,-6464,-1032,1964,-12988,1633,-2355,12187,-7968,4545,-16767,1141,3498,-5688,9560,-6762,4948,6186,1413,-2023,-729,-671,-4455,-2126,-6333,4089,-4702,-3112,-8320,-2220,2978,-9809,7500,-2565,-2186,-5571,15498,-1151,1907,-553,-3479,-1271,828,-5649,-1263,6635,-3405,3898,596,-549,-8950,-4379,-5449,-5185,-232,-1782,6269,-3566,-3493,1252,3725,-370,-5195,-3645,-2819,2678,-4846,-1046,217,-7666,-10605,10878,2305,-67,465,-10087,-559,17,-3125,1501,-1816,-2260,-3769,9501,-1962,-1196,2397,6074,-8979,-2454,861,29,-4667,-1622,1419,-9199,-3427,-758,9702,3000,-3330,-16142,421,-2995,11542,873,-1673,-7036,292,-276,484,-1466,4367,-653,3110,-1541,-2264,3647,6928,5571,4121,-6918,8354,5551,5620,-832,3376,-3083,1055,2519,2452,4279,844,-6821,-10029,-1704,2216,2629,-1450,-3857,1238,-470,1939,-5024,3872,4992,-4172,-2709,1840,1932,-12011,2512,-358,-4475,-5874,-2841,-2224,-721,-716,-1624,788,3356,-4672,-6845,-3417,12304,-4445,-3193,-1483,-838,-5390,4357,770,-1723,2106,7861,-1751,-3337,12568,310,-1733,-1187,106,5019,-4333,2019,-2165,4343,-4594,4033,-3601,823,-6333,-585,-11386,478,-751,487,2091,9838,4077,406,8774,4621,2489,1014,-9477,-1677,1654,1968,9990,-3684,3937,6298,-1480,-786,-3757,528,1529,-2915,7963,-13701,1998,7055,-2119,2541,692,2612,6240,5688,7597,2758,6669,-343,-2457,-4211,786};
    Wx[24]='{-1484,7475,-4870,-2083,-2121,445,8271,-3049,-1505,2729,-5273,-198,-3674,-223,2736,-5830,-8168,4262,3903,-591,2142,2929,1445,1431,-552,-933,2580,1934,9687,710,1676,3193,683,-1655,-1196,-864,-4255,-629,-468,1047,2481,5322,1721,370,1923,2966,3493,-2597,-3049,2181,5546,-1796,864,2335,-1501,3149,-3508,-2131,2304,378,5180,2949,-235,-1140,-3937,3071,961,-4982,259,2468,1427,4265,-2841,-1992,-362,-2103,942,-674,941,4060,-3769,1744,-1043,-4436,-4846,2541,-3500,-33,-476,-1801,-5717,-52,736,640,2150,-1444,-303,-906,-1068,-1550,316,17460,8593,12558,8017,-2883,-10302,17070,-2247,-89,-13310,-1503,1287,-8315,-6025,-9985,122,7626,165,-256,235,-6503,-4216,247,5424,-2426,-2622,-13144,2934,788,-3344,-2302,9360,1600,-4650,662,3823,-5068,-2900,-1834,-3579,7148,4865,2885,3491,-2214,-2087,-7993,-1702,806,-2949,11875,-4445,-12294,6191,-19179,3916,4611,2491,-127,6298,-3825,8227,-7363,-5097,314,811,-34335,-1535,4599,12578,-10556,-69,6333,8315,-24589,13144,-832,-5332,6250,9887,-2980,-2462,-9565,-12578,8115,6166,2229,-4523,-6181,-1173,-3750,13437,212,13076,-4565,3256,-7646,1749,-11240,1699,-10957,-5009,3112,-461,635,6040,-1503,-5087,2604,-424,-3632,1719,-2624,-2008,4584,-2636,-3615,4975,-511,558,2496,102,1311,1816,-4572,1511,254,927,-8251,1989,-2268,-266,3564,-1346,1400,1030,-488,4912,1396,1932,437,-3046,-5610,-3774,293,-8569,1506,-1417,1853,2861,-6918,6000,4904,464,-3139,-4467,1862,-2077,2854,3117,8012,-1289,9155,955,-3068,4196,-1810,1577,-1038,-3740,-571,1203,158,1223,4709,11132,-1575,2263,-2705,-1015,-6083,-2209,-102,-5454,-6,-966,-467,3098,-3696,2301,-4504,-1917,96,4812,3205,-440,2795,4482,-1308,3156,-6435,-5922,4831,2492,10761,7055,770,-1640,6093,-11250,-5024,-869,3803,186,-4521,5288,-721,6235,-4858,6406,5092,-136,-1730,4138,-8129,8291,472,7915,-5893,-1630,-3159,-2147,3271,1795,-1049,-1558,2790,3999,-3366,3166,133,-4379,-4399,-47,3193,2900,-5742,-3354,-398,7802,7866,4418,6127,7939,8364,-4997,-3771,411,8349,-2800,5112,-6191,2656,3591,635,-1462,-1634,13955,8149,3234,-2110,3891,-3771,5458,997,3947,-1041,2237,-20,-697,-7915,-2995,-10087,-9174,-825,-3679,-890,-2475,-2254,2072,3515,-3366,-7573,-2897,286,245,14199,8759,3850};
    Wx[25]='{-964,3039,68,4521,-159,-1945,-216,2147,1508,-5639,-681,618,-541,1530,2521,3051,6782,857,1843,-1031,-1511,647,701,-112,1480,-3037,1525,-1480,3061,-1334,5263,-8872,-463,-3754,-2242,-428,566,1580,2127,-3300,1141,939,4035,-4353,2443,-869,2521,5151,3540,4003,4570,326,116,667,-307,4575,2895,-3227,3613,-581,-1348,3657,5771,-1335,581,-1236,-1065,-7929,-1195,392,-1535,-3408,2741,2719,-676,548,1346,379,4548,-2088,1660,-5820,121,-4079,1584,-662,2448,-2025,1497,5761,1857,-5302,7260,-2305,2524,3632,5874,3664,982,-1921,1724,-8774,-2199,2078,-9316,-1832,2988,6079,-1064,7778,4836,-4802,12011,12412,-6362,7568,3471,531,-2165,-808,1076,4768,473,-3171,2844,4106,168,2148,3994,6791,-550,1602,10439,-3330,-850,-8012,-8300,-1962,3000,-6679,4907,8955,4877,1109,-20253,-378,-3605,-9609,-2509,2795,-19365,-4011,-4787,10595,-1654,3134,3635,412,-901,6679,3471,8408,5058,3679,1844,-3937,4348,18818,-778,1234,1850,9648,3850,-5493,338,5288,12109,-7607,7026,-11308,-1444,-10097,1092,4909,-723,59,-488,-8261,-2612,2326,-4016,-10898,-1881,969,-2370,7016,4892,-6191,-623,-7387,-1860,1776,605,-1435,-3261,57,-1826,-5292,-4653,-1342,8349,-2429,-3608,6723,-6254,1777,7377,467,5507,-735,-587,-106,-1201,-4531,367,-4028,1472,-912,-6308,2990,4814,-10839,-13613,-8676,-4650,-574,-9091,-3522,-8784,-888,-4309,-798,-7949,5424,-2644,-5102,-9365,-3166,-219,3193,145,-404,273,-1494,-480,-10468,2180,-6010,-948,2856,195,-3435,-9663,8188,-11660,-3706,-5244,-2102,859,-1314,-6621,2442,4335,3032,-2912,-8217,-8642,-6860,-1112,-769,67,505,-2619,3891,1282,-1064,-1234,-2032,-792,1881,4201,2519,-4338,-2071,-5361,-834,-1822,-621,-8061,-8793,1256,5878,6455,-1872,1424,-6245,3251,-10039,-2973,-6562,11445,5927,5405,-2546,-8300,-2983,957,16005,713,5996,-5112,4926,2961,-407,3242,4714,1400,-6748,785,5117,6811,-3730,-11640,-9799,2418,819,-1044,-4033,-1024,-141,1395,-2283,3784,1021,2081,-2332,-8227,466,-2014,7221,-1308,-3527,6191,4829,4721,-4587,9926,8437,5776,83,-1489,3071,-1028,1293,-4477,-11650,-3493,-5156,-2731,-1260,4282,-4072,-397,5917,-132,5112,-3486,7436,5737,-3881,-94,3305,1214,-8720,-4128,-506,-3098,-413,3696,4755,6894,16757,1012,-2476,-1416,-819,5561,-10273,-6611,1579};
    Wx[26]='{-447,-125,1287,2673,-460,-1406,-3466,-1964,-1406,-3203,599,881,2563,-1958,2448,4489,-2915,-5893,2070,3464,3327,1652,-181,1114,-130,3066,12,-1879,-6059,614,-1425,-1214,4108,-4165,2683,-1052,-1212,1614,1379,-4187,758,-3503,-7836,-2768,5117,-928,7456,1270,-1084,3713,-5068,-2047,-123,3500,2021,4438,-2778,2454,-852,-1763,-2683,-2060,2817,-3281,2465,-1016,-393,3127,-1989,1824,4953,3579,4155,-5185,2360,4924,-2644,593,217,-4831,-1466,2463,438,-5336,2014,-3635,884,-2768,-1431,2656,-1010,5112,-313,-1871,25,-1304,-515,-3012,-6298,989,2946,-10986,2539,-5527,734,-1929,9995,-7612,-4709,-2805,2139,4890,-4333,-5541,2403,-5307,-2690,6889,-2751,2897,1510,2427,3449,2176,-2249,-11953,-11367,3366,-6738,-7363,362,-1425,-7885,-1257,1250,4086,-17,2580,-1271,6933,-5219,-9272,-11074,-1510,-1045,940,-14267,-3701,-1264,-8525,2469,-23593,-15,3498,3488,-2980,-3017,-866,10595,3540,-4946,-7739,-1416,5151,-5961,-329,-5986,-4089,-651,3886,2841,13798,357,11787,-988,3098,9350,-10488,3503,-10107,-8129,-1887,3205,-22617,919,7280,-1367,-5468,-3684,-871,-2570,-4626,1997,-1815,-2070,-2504,-4785,2639,-738,-7060,1040,-1030,-4001,-1501,189,-478,1586,402,-133,-1899,-1215,1201,1539,-1089,3508,480,3923,5083,7265,219,2288,-16,1365,-2254,-4648,-8955,-1323,-2517,4135,-4729,1188,7104,-256,-10097,4233,3215,-3876,1614,-5732,4782,1240,4582,-2349,3852,-3303,796,5234,-1042,1419,-4641,8330,7641,-831,-3518,-1470,8505,-1159,-5048,1917,3894,-2012,-1654,-7226,-654,-5571,817,-318,-12333,177,4665,-2375,-3283,-881,4824,146,4194,1140,3891,-2597,-2719,-1568,3876,-85,874,-1112,2678,2027,3166,2387,-6079,107,-2968,-1130,-773,-3984,-3457,1945,6743,-4941,-265,-1994,3178,277,-56,3549,-4262,7065,-5395,-4677,-2658,-3959,-1099,944,2817,-2496,-3540,-3715,-3159,6757,244,-677,-1992,-3061,-3288,2376,1446,-6748,-8286,5234,2269,424,4785,2293,-5966,-1140,533,-1451,-427,1855,-640,54,2702,-1617,-2169,-936,-1192,5747,6547,70,835,8652,-1844,-1374,-2763,-12226,4011,1845,7695,1754,-5971,1356,-1661,11435,-6030,-9521,6538,-6992,126,-10927,-1033,1273,-6870,-2391,325,1169,1068,8432,1124,752,-8076,-5131,-863,6435,3400,-1951,5009,1379,3957,4545,11308,-3251,-16318,-1971,-6635,-970,-1040,-2966,1154,-3164,4870};
    Wx[27]='{2622,-3686,-2746,-317,2895,974,-4682,-2670,5268,5766,-3461,35,516,-5703,4182,-3767,2188,1459,1358,-172,3620,-1263,-3537,16,-2406,2410,-2039,2275,-2526,3942,4479,-4101,-7177,-5234,4775,-2188,7543,690,-2397,-4812,-212,-2727,-421,-3254,-10224,1916,-6220,589,-2490,-1794,5620,-3767,-3806,2902,-2719,-3115,-1907,2668,-259,312,-490,-500,-6713,-620,-249,-3454,2103,-11992,746,-3481,-3320,-328,-383,1002,2092,-2907,-4609,8105,-5693,-4709,176,-12548,-5161,-9589,2097,5810,5107,776,366,-2878,1010,-9262,-1878,-2039,-7851,1520,206,-5024,32,-1530,1844,-12734,282,6513,4899,207,6240,-7631,1496,-98,2310,-5268,-9277,7739,6704,-2692,6225,8881,-2958,1591,2539,5200,14833,778,-3750,381,1938,-6040,3913,-234,1181,-6416,-125,-1285,3986,-820,4211,-3229,-1179,-9179,4941,-23671,-11972,6787,10664,-4758,-5043,8027,-1267,9472,4079,-12705,1447,-1520,6391,5947,6494,-5078,5986,2536,-2517,9140,-123,3000,12851,1436,2182,-4772,2268,-3386,-8085,-5854,-2890,15117,-1522,-3686,-7705,-12558,-6899,6113,1039,14560,4167,7158,3159,-12626,-463,-3979,3991,-5834,-4675,6650,-1727,1155,-1149,-10693,1650,12089,-8154,5683,226,1103,3149,-2856,3234,1922,10771,-111,334,1213,-8515,3620,-141,-1958,8461,3718,140,-495,-1227,512,4516,333,-2883,-982,-1896,2824,-5429,3010,399,186,-2832,4929,3913,1036,-1474,1925,-2802,-2971,-2565,-2497,1888,-7207,5229,-1756,3918,-4719,-1254,2890,-1556,5727,-3188,184,1170,361,-3283,-15585,5410,2587,-4340,-9287,-2661,-5268,-1795,738,-2152,-780,2641,-2283,-1597,1165,-1131,-5585,-1114,-106,2834,-5507,-4523,408,4482,4365,-2766,-241,838,2371,-3469,-2856,-2517,-8798,-5747,-959,1958,5410,1761,-92,-1032,9794,4965,7221,2543,-1000,-1356,-6708,-3813,-2377,-1061,-3378,6987,-1228,3193,14218,-7514,2166,-2175,-4133,9428,-528,-2709,-2871,2020,5053,-6689,2152,-386,-1350,6333,603,-5107,7299,-3149,2282,4780,-8081,2088,-7519,2435,1522,1102,5424,-4104,-5683,4030,-2561,9921,-4597,-1384,-10039,-1594,7055,-1494,1997,5693,-3039,-4667,2922,-3352,4396,2624,-232,2260,4721,2163,-2685,-680,6816,2812,-1704,-3769,-2266,14843,-5893,1989,-9931,-3090,3391,-3562,-12246,3203,-3029,6860,-254,-85,-3908,-4802,-7832,189,-6000,4914,-6206,1885,-6865,4960,-1055,-2963,-7875,-1337,12832,2558,2866,2812,-3601};
    Wx[28]='{2086,1036,-2094,-2707,987,3969,1832,1342,-116,-928,1945,-1751,2402,6352,-2712,-734,-286,-184,2054,1049,-158,-3305,259,2220,105,238,4360,-842,1280,-1126,2391,7133,-2486,-3186,-1207,-4096,4057,-179,-1663,-1981,2391,-5200,2600,1273,-103,225,-9462,-1888,-597,784,-5429,-5585,-2812,549,1748,4375,682,-1973,-6069,-1870,4653,1379,1166,-7299,-2980,877,-3830,-7880,2161,3432,1195,-2254,3737,2780,-3117,2810,-1831,-1040,-2396,8081,949,-9184,1610,-4987,2485,-2963,-2178,-1468,2507,1004,-3432,-4111,79,-931,3725,-3078,-457,1568,4743,-1685,-1496,8974,-2347,-11748,1395,-1547,6967,6118,-3669,4287,-8632,-6899,-1624,-8100,-8486,-9990,2607,2929,-780,2705,1531,-2697,-5727,1788,1418,-7031,-5366,4243,-808,17402,858,12304,12343,-18066,-4614,-8051,-4750,3171,5410,2132,-8188,5380,5556,-8876,206,-2243,1015,-11718,5380,-11962,1374,-2949,-8002,12500,-3115,-10439,-13505,1789,1636,3618,56,6855,3669,1534,-9174,-2641,7919,10566,-3166,-1821,9965,762,1545,-14208,-1921,7456,13437,10996,-8774,-3942,160,7993,12529,-13964,-2067,5249,2290,1107,-1412,4313,-494,4057,4890,256,-535,1607,-12880,13222,12460,2432,-2783,-3544,-1021,5605,-3273,-285,-865,938,-1909,-5683,-1722,-1214,-3127,1351,-3791,1750,1647,5668,4309,-1090,1530,-2670,-3166,-304,14,-891,-974,-1166,-8916,2653,3237,-403,-1973,-729,-6220,3847,-6635,-4536,4621,3588,-1267,-7998,126,-2058,4184,-665,-10166,1190,1168,2707,4572,-7436,-1965,-1669,702,-1943,1689,-487,-11210,679,-2387,-5234,4077,-3432,-6074,1953,-6362,-8261,3674,-1130,950,221,1560,2619,-2590,-6474,14980,8623,3781,5581,-7377,2137,2053,-2136,-5302,380,-1811,1990,5927,-4379,-1234,-5126,6865,1129,4704,1774,-1544,2597,-5239,409,1405,-1668,-4653,8193,209,-9038,-5854,1304,12001,-12148,9414,1938,1271,5156,-11367,772,-2526,6923,-2753,1285,-7583,-1850,-181,2797,-4038,-2570,-2492,-1510,13017,728,6347,2416,-252,930,-1387,-4958,2529,-8500,-2364,1956,788,8359,-3364,2150,3884,5229,-9003,-4760,-2919,-4758,2851,-1400,-1975,5092,6347,1901,7524,-5439,-8544,3007,-995,1925,-1788,-4826,-4479,-2988,-12236,-3317,-975,-1008,-6000,-29,374,4311,-2644,-4677,9902,10449,797,2897,-11425,1226,4077,-140,6943,6962,-211,-281,7998,17275,-6113,-1662,2829,1409,121,-4548,-3977,1708,1178,4597};
    Wx[29]='{863,-5468,-3239,-3564,1238,60,-1130,-3410,-447,1319,2951,-497,-2934,-7202,-5175,-12304,-6708,-343,-195,-2558,-192,-2963,-4753,-3334,-664,-2250,-1973,602,-1166,889,1912,-8427,-626,-7050,-1331,-1414,-694,-919,-2724,-3820,-3847,-2041,-5234,-4907,-3000,-2327,-9541,-6923,-2827,-2324,-5322,-4636,6230,-4628,-3886,-150,-1049,-2675,-2188,5444,-2529,-143,-2727,-7783,-7026,78,950,-6376,-820,597,-4924,-4909,-2470,651,2072,-5332,-1174,-723,-4812,4145,1144,-5556,-1932,-4445,-231,-831,-2254,-210,-159,-1127,-741,-5190,-946,-2502,-3679,-1429,-2734,1691,-2583,-8720,446,24902,1676,929,2252,1398,-5805,-123,-1793,-7182,-1989,476,-1391,4357,-7075,-10585,5034,2636,-4536,-3850,-1056,-55,5429,-10029,3505,2893,8505,-948,4064,-3439,596,8911,-5742,12070,-608,7241,-202,2008,-119,-9545,3635,3835,1287,9467,721,-1621,-1260,7158,-1757,4836,5776,-15498,-52,-2464,3671,10205,2685,-261,-3942,1451,-2139,-6362,-6440,-8598,3762,-834,-3107,293,3728,3540,3005,-4897,3581,-8720,-977,3195,-10351,17587,2541,-3027,5805,4655,-1097,12363,-1139,-8339,441,1262,-1508,309,-2805,26445,-51,-2493,-9340,-4953,8496,9321,2917,13457,2241,-5351,-1557,-847,3886,2083,438,-2683,273,-1392,893,-1854,764,-3898,3833,2841,-4685,-3642,5649,3342,207,-4096,-491,3137,1666,-3659,2978,2017,-1541,-1578,1534,-1001,-3688,-1785,4548,-28,8515,2534,-10839,2330,3452,5234,2083,-3610,4018,-4904,8505,339,-3625,2666,-5097,-1922,5668,6875,-4140,-4399,-3801,1663,-7666,-6044,-4042,-1682,6430,-1061,-2320,-2237,-670,3254,-3081,908,-3007,-6708,-4335,-8833,788,1141,1477,1552,1254,-1759,-942,-7045,4687,861,945,-7104,-853,3046,7177,1838,2807,-513,-667,-3510,-68,-5024,-5903,-2224,4404,-2861,3671,-69,4084,164,-783,16650,-348,-1827,-4089,-4721,-1535,-263,-5058,-4575,-1591,-4062,-5292,-3867,11953,-523,283,-2030,-1802,653,3127,-7314,2094,3911,-6181,-6093,-708,-5273,1986,-574,-4130,1799,-3889,7294,-10585,-5541,891,-6152,-4113,-1302,-5478,-11259,-507,-9106,-2243,1983,-2463,-5556,6132,-795,-2204,1506,-2705,-6997,-855,-6660,-180,-428,378,242,-817,5200,5761,1044,3176,5493,3576,-13369,-130,-4567,1528,-2165,-2028,-3088,-1307,2342,-3208,-2114,-7495,-2551,-3945,-10166,-563,-3022,-7563,-5576,7055,-1975,-94,-12675,-11962,-2678,9428,-1040,5253,-6601};
    Wx[30]='{2231,-14150,-1365,2551,-953,320,5644,-5390,1663,433,276,-659,454,-2783,-4028,-7587,2351,3859,292,356,1733,531,-1813,-3845,-175,-466,1402,398,3369,-1240,-816,-572,-946,-4482,2114,1503,1212,-197,-318,1303,1251,-2399,-7221,-4746,3173,3640,-5937,1196,2034,-62,-3601,469,-3342,-1951,-3527,-3806,-1790,2464,-1335,824,-1772,6977,1231,2539,-1074,-2449,2369,664,1047,2734,184,-2016,-5424,-584,1877,309,-1146,-2370,-2548,-1203,2088,-3388,2172,-166,3027,823,-1441,-3818,1572,-3112,-348,-3618,77,730,-6313,2719,-2100,3620,-6635,-1765,-1513,-137,2315,-4682,2224,-1311,256,-11464,8750,959,-4265,1846,-2604,4785,-728,3266,20019,-7114,-1779,-2766,1745,1271,-533,-1600,-3947,-8144,6484,3833,-460,-6123,3659,-5336,-3549,-748,4882,1546,3779,-3171,-3154,5268,598,-10849,-518,-1258,4113,-5166,928,-2283,3623,-1831,-3759,-2644,5722,-2597,2858,8466,-1016,-39,4670,545,1608,-4528,-3259,1109,9365,-139,-1470,6196,-3095,-68,-13974,-5253,-3486,3698,-618,-7299,-6704,217,-2841,-7543,652,-6977,-186,7832,6235,2303,-1923,-267,-725,-3488,2739,-1901,1994,573,1374,2457,2683,531,-3759,2958,1781,15468,-1172,27,3842,579,1958,-4499,-1144,2961,182,483,383,3583,-1251,-2624,6987,-179,1176,-1539,-1445,-1234,882,-2006,1494,1640,-582,-381,10029,-5610,-6176,2403,737,6284,-3586,-6870,-4914,2106,850,2246,7041,4814,4650,2429,182,7441,1749,-200,573,-629,4384,8618,1439,3696,-3994,-1988,-1199,158,4711,-5805,173,4035,-729,2919,3813,-2371,5937,4589,-1870,823,1071,-1791,805,3291,2161,1206,640,6040,-1464,-3452,2932,1678,-1860,-4077,-2298,-1636,1152,2592,-902,-697,8,6250,-4697,921,3049,5834,6523,40,3237,431,2919,13164,6206,-466,1781,5175,6914,-5170,-5932,-2670,-8315,322,124,5371,-7797,-7685,8500,4140,-4338,839,3508,668,-5537,526,520,916,-136,1342,13398,-290,-2841,2009,-4042,4460,-10898,-3188,107,-219,4345,3481,3742,9765,3510,-658,1004,-2022,2543,6342,-3872,3015,886,-5029,5078,1518,-4201,-3203,-5200,14023,1718,-3525,3588,4003,-656,4189,190,1872,6396,2907,3913,8876,2558,5385,-249,-2592,-1881,5122,4221,2807,-4536,-3559,8803,2250,-653,5839,-5141,8286,209,-2436,3164,4926,-4,-523,-3645,9594,1058,7548,10166,-299,230,5102};
    Wx[31]='{2614,3015,-81,456,-994,-2834,232,5268,469,2296,3713,738,1759,6352,-1688,3247,4172,2902,3249,511,-1168,343,-1514,-1536,3403,-148,38,2298,2888,-3828,3078,2376,4829,1922,3923,-403,-1198,-2841,-1346,-192,509,-2207,-815,526,-7729,6333,5961,-504,-1165,656,-4487,3730,-7353,-53,-8281,-5766,245,-5517,-2437,836,4045,3007,-36,-263,7968,2491,2215,2281,-2841,-74,-3833,312,2597,-4599,886,-1232,-344,2484,-3205,-607,2705,-523,1446,-1047,-889,952,-4318,-5161,-983,-265,3676,-6987,1156,-2636,7412,7495,-991,-4265,4433,2949,-988,-7597,-3601,-7167,712,3486,4440,704,-1608,1630,-14179,6391,11328,3151,2487,3962,141,3466,-1545,-4550,-4953,-3452,2792,2700,2604,1430,-7138,-3054,2440,7583,-7695,-13115,4174,10605,6787,5483,4909,-1549,-9355,3874,2257,-1584,-1717,6997,2653,7363,958,-1311,-2159,1330,12597,13730,-19257,7617,6416,9331,4467,2648,-3129,53,3359,-3388,-5815,3686,-1572,3034,-4655,-5507,4814,3513,2497,-10429,-8823,-7192,4252,360,11464,-17402,15224,-60,6835,5444,5341,11005,-632,3498,2194,-19785,-220,-9038,-8061,6157,8374,1502,1834,7182,4042,-3750,2597,1959,1997,-6318,5278,6440,1915,-1102,3430,8715,734,3610,4680,1782,2478,-4897,-991,2001,-2211,-78,3420,1300,-124,2274,-2145,4968,3398,-3840,1827,593,1181,7973,-3681,-8110,-3808,1888,-3376,7949,993,-2241,1059,1206,-362,-1168,-2023,6293,4150,2176,-7661,916,-1654,5917,12460,-3112,-416,3845,-562,221,-1079,-5380,11376,-3530,2653,9384,1150,-1420,-4541,2019,8725,-7661,-2365,-1888,-1378,-1032,401,9077,1052,4382,8164,11542,1641,-6074,2147,-16396,-1657,-4157,-4104,-1613,-77,1276,97,-3459,7910,2386,1245,-2910,-11357,3442,5366,4692,838,-453,1766,-11943,4719,-106,3078,-4299,-5439,3862,3454,11650,-2467,895,1112,134,-2597,488,745,-2897,4221,7265,2741,1674,-3281,1236,3085,-555,4819,994,-1800,-550,-4750,-5556,-229,6450,-20,3601,-2722,1390,-960,3774,2998,-2592,-9702,-1314,-7358,8535,7631,-68,-4919,509,9106,1496,-8676,-6411,119,-717,1271,3833,3547,-6010,2088,3959,7617,-4816,205,693,10976,-3925,2624,773,-1240,5000,-2208,556,14140,11855,-7250,770,-7685,-1243,4663,-7412,5244,-3732,5849,2788,-386,-8457,623,-4948,11074,-5151,-1376,-1892,-5366,1143,-273,3645,3776,4074};
    Wx[32]='{968,1072,-785,4270,-2056,997,-444,1931,-1044,1503,-11259,-1184,-1012,-2600,701,-1490,2780,-6284,-289,1439,2452,2761,3476,805,2790,-4467,1064,-476,-123,-430,-737,629,879,-1854,378,-841,-1423,916,717,2385,-186,-17,-7778,4003,-6118,-27,10947,-4370,-3212,-4584,1590,3276,1623,-1867,3149,-365,-1564,784,-1846,1652,4870,781,6166,4223,-4619,440,-72,-3835,1348,-1944,-1428,2265,-115,-2871,2457,-1752,-3208,-1081,1418,1534,134,4599,1949,-2145,1702,3193,433,5922,-3491,-261,2836,-1643,-753,-572,5107,2663,-495,-9223,795,267,-791,-10429,-1134,20,2135,-2467,-4875,5058,-1018,-1359,979,4890,-946,-3808,5087,-3300,-22773,6201,357,4707,3037,1109,-58,-791,1955,-3493,-6298,-4108,12070,7592,1306,10283,-186,-5014,895,-1616,-3359,600,-2539,-1271,5869,3862,3620,1765,11376,-4047,-14179,-305,5717,5249,866,4497,7119,2770,1091,3984,2766,2476,-4079,445,5424,-151,7504,-986,-11464,-4802,717,-8344,-437,-1130,4909,7636,1246,2944,6474,-5590,3830,6166,-12636,-1296,-731,9960,8842,-1188,6538,-3803,-1387,8256,3134,-3854,488,-2827,2088,-4194,6083,991,-656,-11250,-7158,-9052,-2529,-7617,-1068,-824,-3139,1586,9501,-4677,2814,-1229,5981,-1322,3095,-6123,4189,-3544,6040,-1951,1291,-727,-321,-2403,2296,-1336,6474,1193,-4155,-1614,-7250,7514,661,-1071,-1453,4255,-541,3349,0,2592,1457,-1210,-3891,1575,6855,5581,4799,-676,-6127,-3723,5058,740,-611,1403,5786,7758,-1693,-4750,6811,-1158,-934,-3217,5087,852,7978,3276,3786,4526,1761,7255,-1122,-922,4895,2039,-1986,6440,1430,-3657,2049,820,-709,13,2277,0,1328,6367,93,-1789,2766,-3850,5590,-904,3898,2248,-1411,3288,5429,-201,5703,-3747,333,176,-2863,-8222,-7578,-5727,2702,289,5317,-174,-805,7988,417,-4936,5180,-1567,-2695,1079,716,-7524,291,2160,1633,2282,-1436,-396,3115,-6406,6162,-2766,-5375,757,-3581,439,-1870,-1291,-1386,4882,2232,6606,-4519,-4899,-3908,-1223,1134,-3208,-5009,773,6098,885,-2802,-2832,-4460,4064,5869,839,6333,2498,-1574,3205,288,1520,-3459,2539,90,-5468,-3251,3854,4868,2983,7172,-10185,6303,-1649,-4057,1409,5214,-3195,-1502,-264,-524,472,7104,-2595,9311,5683,4355,2709,2080,-1394,2988,2668,6694,-10117,-1763,-7553,4926,4819,6542,1191,301,-1662};
    Wx[33]='{687,-2313,653,-1684,-538,908,7,-1911,-5532,-2407,-908,-2949,1148,-2402,-8837,9653,3964,-6635,-376,2349,-1147,-1293,-1322,-1771,1184,994,-1931,2220,3164,586,632,1448,-1627,3269,-2519,536,2900,-1213,-2897,-5517,1589,5439,7749,499,2059,5771,1408,190,-3798,1621,9975,2592,3383,4099,4897,7231,-2382,2042,-4023,5014,3513,5283,-1903,885,2427,1341,-3730,5449,-2924,-3728,-28,1275,996,-1101,2309,-7656,-3852,-3691,2160,-3928,-2393,76,3181,-10009,-2144,8789,-406,1104,5048,-73,-5468,-1428,850,1898,-2038,-377,5859,-8349,1666,-270,-5473,-2373,-523,-6777,3811,-1177,-7050,-4592,-2805,6542,3562,-5620,10869,-10351,2475,-1993,-2265,10048,4104,1337,567,9902,-11435,1573,225,382,-2514,-6787,-3750,-107,3024,-17832,-6494,2069,-7841,-2470,-1848,-5585,-4084,-9926,3884,-5380,7138,-673,-19169,-17617,-3493,10195,-11337,4196,9755,-11113,-5771,1365,1209,-11103,-442,310,-1843,-5395,-737,8115,-2082,4216,3366,-1931,-2790,-1859,1412,-164,8588,1489,-1735,5385,-430,-8305,-12910,12929,6953,-863,-2958,16220,1517,-12666,-1688,20878,-96,8686,44,-2305,892,5932,-7324,-448,-4826,-2941,5834,-12236,8076,-9121,-4418,-5214,-1420,2222,3798,751,1254,-122,-353,-2075,-2666,-888,-1387,-4162,-14638,-6079,-5332,-4418,-3571,570,-1635,-833,3540,-499,-6264,-6025,-11953,1011,-2292,4558,4362,-5751,-267,-10292,-4243,612,-7680,-4040,591,-991,-3481,2592,2595,-2717,-1184,-4721,5625,5190,4414,70,-6074,-2736,-304,-1187,5913,-5522,2668,-5117,5742,-1211,8007,-3222,-2183,-198,-2445,-7587,-5395,-4794,2249,-2883,-601,-1466,-2142,2927,1206,3703,98,-6708,382,-1400,-4946,4851,-4870,1674,-3515,-5253,-5312,-2990,5249,-567,8413,-1018,3537,-1781,-397,-4382,2509,-238,-2678,-3110,-4011,-941,-8261,-4787,2294,241,2442,6181,-7441,-1650,-449,1571,699,-4895,-15625,56,-4353,-13398,3354,-2222,-3337,-702,3603,-3271,-6181,-2976,-6875,-133,-4074,6430,4001,-184,3625,-8007,-1300,-1557,-5253,4975,-4697,-4270,-3552,3325,4086,2758,-129,-537,2595,9218,-5029,1624,-3244,-1915,-1186,908,-87,-6113,-1033,5224,-6069,-3608,3315,1740,-3518,421,-2531,-16083,-3471,-6948,834,-4152,1118,1920,-2086,-12753,-2731,2467,-5976,-6884,436,-2609,-7788,-368,-4299,3981,-22539,-4743,-7705,-7539,-524,-1538,-2587,-3527,-56,-1650,-1630,-2578,-1704,-7265,-7729,-22};
    Wx[34]='{-390,-1538,-456,573,124,967,555,-8867,-2900,2125,183,100,-1728,1827,-1517,-3212,-2066,2980,854,-1718,-1474,1063,-1401,-1264,474,837,1022,-1088,-3063,2114,-5209,4997,2868,4628,453,1270,-3537,-1387,5039,5605,-371,2196,-1821,4433,1179,-223,154,-1405,-491,-1270,2568,2797,1424,2661,5219,-100,3491,-913,1958,-809,1820,2500,83,-391,-3559,1385,2117,5590,-386,2092,2724,-1221,-1655,-1151,-5927,-323,10537,2252,1400,-2207,1617,4001,3339,5058,-2067,5156,1387,2309,-2844,-4108,846,6513,697,-2115,1434,-2888,2551,-6547,-1571,2349,-5014,12773,-3798,14765,-1206,1927,-1258,9096,2126,3,1197,-7348,-1462,6577,563,9907,1469,-3510,3720,-3,580,-6157,-179,5419,1407,7060,5932,-1563,10761,6752,1809,4462,4406,-10546,-2614,1950,908,-651,-5014,-3271,6582,4423,11572,3298,2917,-11904,12216,2746,-7866,-4299,-11259,10351,-5708,-3215,-1772,-16210,5859,2487,8603,957,5717,12597,7675,689,-8051,-546,9487,-20273,1557,-3544,-14287,-12861,-6420,-5458,5576,-8925,-7368,6181,-9301,993,5878,3933,3569,3566,-3415,2565,2294,-87,1148,-5727,-4489,-14091,-405,-1508,4494,-4169,6313,7553,223,-4653,1312,4804,333,-164,-1223,-939,-2119,-3227,682,4235,274,-1303,479,-5424,-176,-391,5629,-2604,2283,2958,-2883,2636,164,196,7285,574,-1068,2014,2534,-9804,1209,155,-3383,1223,7568,-1656,-3627,2026,-3957,-825,-2727,-4370,-3671,613,-4104,-1986,7451,-6796,-4560,1074,-1990,-8125,-2137,-1406,2043,6904,264,99,-5883,7231,-3229,-10673,1381,5029,7543,1063,-4104,-7915,1549,-685,4504,-1715,-1416,-3898,1284,-1608,-5688,-6840,2163,2469,-2030,3566,1982,1864,-5942,-4123,-3071,3645,3041,-4060,-4851,-571,-4345,-1838,-13320,-2254,-755,-9433,5468,214,2366,2,8691,1594,2578,-503,-3496,-2756,-1401,-186,-2551,-4379,3271,513,3476,1794,7885,-4228,-1060,4409,2467,657,-4138,1094,515,-3085,6577,5800,3759,-4890,-1906,-5888,-8408,4008,422,-1221,4575,-2663,-8779,-610,4968,54,-5654,3869,50,3596,12236,-3735,3029,-948,-3864,2783,-3959,-926,17753,11357,-3159,-665,4211,11367,392,-3864,-15283,6215,-3784,12382,-2578,1121,9604,5903,4680,-1195,-4533,-689,1033,2690,-4892,-7241,2467,3356,-513,8403,411,-3066,12617,-5434,3320,4907,4912,-4257,1010,-8149,773,8984,-10908,-5336,917,3586,7182,-3806};
    Wx[35]='{-198,-4685,-1555,-895,2097,-40,4731,-3317,-421,1031,-408,-1434,305,2521,-889,3999,-1082,166,598,2127,-470,-2956,-1912,4494,-2384,1372,-1427,-74,-14,3842,-817,9672,-1904,2939,245,6381,-2121,958,-2493,2060,866,1728,-1267,-684,3366,5068,-4719,331,3046,141,-2502,7480,-1751,1356,-2452,-5898,679,3796,-879,-944,-2493,-230,-1293,-706,2753,3361,-2602,8642,3220,-3303,-621,3325,289,3208,-1400,722,4658,1012,-2573,-2297,4833,2221,-1621,5507,-2741,3474,2199,4584,-3293,1352,3076,2744,-3076,463,-5034,3366,2194,-2995,-2095,-1560,-2086,-1296,-1063,-276,-1511,914,-3671,3557,6206,-4965,3947,-3652,523,-3435,11064,-3767,-8901,2583,-1243,3540,-1881,131,5014,-2054,-1975,-21,208,6997,7846,-11523,6040,8066,8916,-3066,7343,8823,-251,3041,-8452,-8247,4362,8330,10898,-9829,-7241,-12314,18164,-1243,-6450,9863,386,1402,7792,6528,-1968,7421,-3315,-1596,4616,3388,2354,-2800,-11835,-694,-4511,95,7368,3771,2558,-4584,-2519,2065,-969,-11933,3071,-21835,-976,25019,-3896,4313,-2216,22539,828,-7431,3395,1735,-558,10654,870,-759,-9741,5434,5742,-1968,362,2888,-60,-8334,1345,-2736,-4252,6425,-941,4833,-1275,1909,-4973,1044,1859,1085,2824,-1285,4213,-4663,-4411,1691,-250,347,-1195,3876,-2055,-539,3496,1183,3791,3417,-522,-2678,971,4748,1889,975,-671,-1062,-327,-3354,-2797,3942,1064,1467,-727,12,-648,5942,2788,1971,-1242,-3676,-3112,3500,5346,-5039,1494,639,-50,-4565,-2656,2177,641,-6899,-2919,3195,5712,-3276,143,3955,-3491,-12197,716,-6914,-1859,4277,-130,2763,-2127,-12939,-1530,-1972,-4797,5244,-1966,-31,1099,-2983,-1016,-6118,1367,-855,4370,3962,-2746,-6035,-4082,-2290,906,-1168,4731,-94,-2309,-1461,-6093,8691,-4338,2059,-567,-10039,-1816,2084,3688,-4064,3300,411,3793,4462,2556,3371,6821,-5458,1089,-4858,-3747,-3583,2734,6552,-3339,3554,-1988,-6367,4328,2388,1480,8701,-8251,-3620,6508,1749,918,1833,-1673,4599,-1447,6367,947,-83,-3569,551,414,-5371,-2105,84,4233,-4777,1555,-3393,-6113,-8486,-5278,3142,-5961,-10673,-1308,-3212,691,-1549,-167,6694,-8032,-715,-4914,-12871,760,1153,-913,-84,162,-5683,-3854,13,-425,1810,-2463,5273,-106,6381,299,-814,4067,830,603,6865,-513,-6323,-4558,14511,-405,7802,2374,5249,-3249,2534};
    Wx[36]='{459,1117,-1539,148,-646,-4135,3310,-2366,1102,1804,536,-695,2403,-469,-5214,2128,-5688,-353,-607,892,-4111,-257,4572,355,513,-296,-177,-340,268,2178,328,-7084,-2871,638,-450,-7,4174,-1171,-2377,-4257,3593,2305,-1492,-7656,6547,-6352,8520,2358,1984,-1385,1473,-562,2404,2352,1418,-4550,-167,-1161,-19,-314,237,-1459,250,-752,-1624,-2158,-815,-4133,-1049,933,642,-3322,-1958,2976,-1003,-3518,-565,1616,-1112,-5698,-433,-4291,2519,-4965,107,-3679,4135,-1848,1319,371,-1317,-957,5307,-2514,4418,-676,-347,254,-31,-885,-1085,-15097,-1585,2258,-3002,3842,-8286,-12666,-5429,4453,7153,537,-5502,-3410,1339,12939,19550,3105,6401,-457,-589,-1414,-3317,-4858,3950,-3237,-4887,915,-4157,-2156,1306,6489,1507,-534,5708,-6733,5405,2858,1416,16191,-2683,1204,-5449,3869,-7104,11484,10097,-7875,8276,-8852,-8383,1389,-4589,-2102,6435,3854,-5795,-407,6367,-664,4431,-1961,3017,3317,2117,-679,3693,-10976,-218,-1539,1795,-5820,2932,1766,-1662,-12304,-16914,6181,-7382,4538,-4555,-7573,-2841,-2954,546,11845,1496,-70,1477,-1669,114,4895,-4077,102,682,-7578,-2353,7041,-505,-8559,-691,2812,-964,-473,-416,-876,2961,-2290,-1921,-2058,2009,1862,4411,5185,-2646,9140,-1591,-2396,-1608,-599,-439,2653,396,1089,5019,7661,4255,895,-6928,-456,1580,3962,147,4707,-8442,5708,815,-1568,-3579,-3847,-7470,-210,-12333,6000,8710,-7666,3920,1826,-352,-4262,-1106,-8452,93,1638,-221,-871,-92,-4943,-2922,-886,1442,5063,-8876,3076,-1047,2156,-896,7963,2238,24,12089,-1832,4924,16,-4323,896,-474,1756,-2117,1552,-4858,-2232,4040,5385,-315,587,551,-1717,-2578,-1705,-1427,-2398,487,-601,-5874,4357,1562,-2379,1601,-3676,-2539,-2922,-5922,657,-3178,-12148,5292,-4555,1733,-935,-366,-671,2224,-2176,-1962,920,-1833,2514,-9741,-5839,-9472,3271,3073,-1258,5649,-3337,3041,-5874,447,-5141,-4677,5166,1719,-1790,2980,2260,1269,-4809,8662,1979,-3686,783,6000,5683,4191,-9008,1768,-1389,5292,-1213,3554,-5341,3476,4912,-8334,-1728,-2700,-2539,-4406,5800,776,200,-6074,-108,3449,-290,-5585,1752,4602,-5019,3364,4465,1743,-406,-5307,-1909,3093,-1578,-1434,-9008,-1656,-3601,-704,-4694,-9770,3005,5537,-1652,4282,-4682,-1043,785,3061,2829,-498,5200,-8164,-3979,-610,-825};
    Wx[37]='{-784,-660,1374,35,1210,-2098,-618,1026,-1065,2812,5117,-299,210,5268,397,-1741,8852,2060,-1492,-78,-1707,1971,-252,-527,-2193,443,527,2521,-1915,1352,-1673,-1163,-2399,-1478,-2846,-1467,1865,1734,3857,4938,-1141,1552,1601,291,7529,515,1988,1430,3691,1340,-4714,4904,-687,-480,-2209,-3337,-3403,-4367,1932,-4169,-8266,-1384,-1198,-962,5161,-65,838,6313,-2053,1767,0,7622,-140,-2387,4826,-179,2966,640,2187,5097,745,6679,-1023,-3190,-861,721,-809,-3818,-94,-2229,-2083,1030,-1862,431,2810,-1017,3862,8637,-1955,2119,-5751,-14814,1333,-1140,3728,1100,-2333,-6967,-245,-1931,-21113,-1911,-2509,-10244,-10009,3603,11621,-2467,4465,-4067,-660,4682,9892,-3337,-1682,-12158,124,1983,-7714,-7475,2011,-3703,6669,-2,2039,4477,1046,3178,-2022,-7236,4338,-6796,-4418,-5859,5810,14609,-6440,-8779,1196,-485,16,4589,-7724,7910,-2246,-4880,866,1713,9770,-2646,1622,7299,-4499,8525,-393,-3342,-1473,19892,4855,-1279,9941,-9184,-1052,-1240,3464,-5776,-2893,3576,8642,-5244,-1713,-5898,-2277,-15888,-6704,-11738,-838,-1381,2392,-4150,-4116,-2880,1652,1160,7275,1693,-1065,7016,1679,-9438,871,4912,-887,1687,2137,-1552,6674,1972,-4274,841,1401,3774,1624,891,1694,-6591,2814,787,-3781,-817,-2375,-3027,-2281,3918,-2807,6782,827,1376,13876,-491,-828,3417,247,6591,-7094,-408,-8120,534,358,-527,-1406,-1677,-1370,10898,-7651,1619,2171,2207,-2626,3698,6157,-6655,-897,-7368,748,-2292,-3532,-6000,535,4401,-3215,2565,6254,143,2086,3295,4013,-4914,-4384,1867,4384,5019,-1600,-3933,1060,-4597,-1381,-844,6674,1710,-2614,-2531,4189,-4665,-828,-9799,-1040,2929,1557,-1889,-881,-2153,-4377,2344,-192,2170,184,6884,-3115,4396,765,13574,7412,8330,-1190,-4023,4609,757,-490,-8530,4262,5883,1928,5952,-845,-899,6801,5585,-2121,4003,734,-651,-3225,971,-3264,3288,-869,1120,10751,3891,566,6152,-2524,8881,-11435,-2861,-6879,-5405,-3356,8491,3271,2382,3850,19335,829,5317,5834,-1708,-3635,-54,8081,-8974,-275,1962,-1687,4172,4033,3813,2324,-23,4152,5444,10458,7949,3857,1157,5874,5351,-6425,8452,2110,16279,-1766,10185,-1857,-960,7900,3654,7490,1932,-1807,1876,6645,1535,-6875,9584,2829,-3767,2561,5605,-2324,9521,-3269,6035,2200,-290,-2666,2049,-1030,6596};
    Wx[38]='{-501,-4880,-1663,1889,-192,-349,-1437,2294,3481,2944,-1040,5151,-2651,-981,-3181,-1503,328,2661,-530,794,678,2910,-649,-1629,2512,-993,3735,-1978,-5410,1196,-2181,-7153,3579,-6586,357,-975,806,-54,466,2199,-4707,-6367,-4550,848,-4716,2612,-3527,-1605,3251,-3583,205,-1116,-3041,-2775,-1665,-591,-2005,-3601,6030,693,-5766,-6210,-901,304,599,2722,3237,-7963,946,1701,-3308,-974,-1790,1348,173,-5913,2873,-2045,-5566,-1694,641,-14794,-2973,408,-29,-3176,1781,-323,811,1121,-780,-6596,-2653,-872,3708,1926,2819,-3078,-2393,5200,-1638,13691,-798,5429,-3171,-2978,-2177,3464,1822,-3605,-11210,-4204,341,1549,2355,12695,1679,-6694,2470,-1552,637,1455,-236,-70,-93,-240,3920,5039,1925,-1259,-939,-4077,5390,183,2149,-3862,-2622,1596,4553,-2736,11142,-12011,8867,5307,-8242,-11416,14345,-1837,-384,13291,-1538,-8857,7973,3044,-5644,-600,4909,2666,-5952,453,6196,-9687,4875,-2770,96,-4296,-213,5083,1906,133,-4069,-9873,2832,9072,2381,-11132,-5932,-2553,7216,10195,2137,6430,-2832,-2115,-2749,-20078,-7807,-150,2032,645,-197,-6669,-4726,2393,9399,2102,8208,-3435,-2167,-1210,1350,12578,40,-2436,-1003,400,3173,5830,-1384,574,5961,-6977,3996,5180,961,10566,475,3959,-3168,-2868,-1057,-2487,375,3518,2094,6503,-1420,-150,2768,3308,-1939,7646,2802,4907,3547,602,-2927,-4116,8139,4184,5019,6923,3732,224,-14316,2398,-9575,-3251,482,4997,-3027,-4191,-1245,-3381,1650,-4853,5156,2479,434,-3549,629,-1240,13134,8159,-1988,-2221,1076,4353,1872,-819,4958,-3000,-22,4956,715,144,-4968,7592,4895,3674,1651,-7299,224,10224,3420,-835,3710,286,-3869,4345,5087,1550,2480,2110,-3464,-5830,2573,6713,2609,7817,3017,5009,-4277,-3461,2680,10009,2912,-770,-2010,-9282,-2390,2172,2050,193,483,5161,8159,-3100,-7294,736,4882,213,-1501,145,4599,1473,3125,4057,3889,2314,-5166,2049,-2396,-3225,4086,3112,-301,2436,6840,-1336,733,5126,-2595,-8237,-10478,3676,-2441,-1494,3588,-2893,42,-5512,-5053,-2692,3764,-226,2332,9360,-181,3908,1093,-1071,2324,6523,1147,4323,4707,1767,6699,7578,-7387,-2341,-689,5175,986,3559,-3576,4157,-4291,3530,-321,1279,4931,8876,8823,1544,6401,579,-3369,-2653,1511,6674,-2219,-1937,-9047,-2727,2125,9428,3457,7460};
    Wx[39]='{52,2357,1258,-1104,205,694,-996,1374,-170,-2656,1164,91,-3745,-852,-1431,606,5620,-3068,-295,2873,-3286,4816,3857,2387,2191,-1256,-1023,-1235,-5449,-2746,-595,-12412,-3354,1196,-159,4096,-3847,1929,-4841,-6127,-4160,-1866,-53,-2963,-7275,-4909,4843,-2385,4299,-2343,-5336,-3369,-1011,-4687,2266,881,1008,-1530,-1276,-784,-3457,-6752,2858,1232,-4536,-72,1108,1010,423,-1452,-2407,-1798,-3940,5483,-1492,-408,825,14,-577,-1279,250,2600,-597,-5195,489,-4978,619,-65,2531,4912,4377,5786,-98,-6713,3759,-960,626,403,-3845,-3913,-3540,4621,-1901,4719,2464,-3176,-5004,-12666,2080,5893,1560,-37,-4975,4780,489,-5522,3847,604,1369,1322,-3249,2700,956,-1472,5087,-2191,-2707,-1292,1721,2406,270,7866,-1247,2138,8,-2729,4743,1315,8925,-6181,3603,8188,5395,4602,4914,-872,859,-10839,2905,1948,6425,13085,14521,3762,2006,8051,-7690,2958,7773,3156,3879,2470,-7436,-1838,7045,1789,-3164,-2462,-608,-1201,-3676,8198,1440,-2486,-1927,7963,-12519,16318,-5102,4797,-5068,1934,3730,-27148,-5683,4519,4169,-2432,1778,9316,-3586,-17031,-336,-559,-5805,-3046,2475,-10107,-1811,-2790,-3364,3903,501,-2702,1104,-274,9326,-5922,3686,800,1549,-237,9223,-242,4938,4719,-3806,-440,-792,1748,-1700,-1679,5258,-159,760,2145,-2998,2587,175,-2429,-1997,12148,11289,7983,-798,760,-1289,-1324,6748,2141,1156,2551,1080,3999,4477,5209,1306,4501,-470,2790,-5410,8041,6538,-4838,1575,-1755,-1761,-447,-2237,2951,2277,2237,143,906,5942,-3562,1804,-11542,728,1217,2651,5581,-2403,7124,-600,4760,5693,1026,-2592,620,-2016,-5888,-3635,6630,-3791,1403,220,3969,-985,2045,7900,-3652,4172,-1010,-7036,-1954,5820,-5615,8359,2449,788,-175,-4819,-2463,2666,10742,10351,-3991,-246,-1993,-10458,-6269,7553,1496,-426,-5297,-1779,-2165,1379,-2221,-2531,-1989,3034,4362,-651,-1039,-2476,2368,-2556,-582,-1248,3410,-3957,-1291,5844,-344,5708,521,-39,-2437,-2634,-693,-2827,-487,-1169,1755,6484,-1286,-2685,-938,-351,273,4221,-4687,7514,1134,-626,2592,-7832,8574,1668,-3862,-4648,-1129,-2741,2795,9555,-3366,9140,4711,-4511,7636,4069,-1794,951,4411,-1927,8603,-5131,-3823,2004,-1044,-7558,4995,990,1623,-97,-421,-3947,17714,4636,-7436,-1198,4809,-5244,-595,7617,5527,1883,2924};
    Wx[40]='{-586,-165,2381,492,-830,3239,5913,755,3110,-1773,-4555,133,-500,3957,3244,5034,-2297,-1275,1021,-2264,-2177,-917,-449,-2425,-2763,3088,3183,2526,3493,-527,4326,-3056,-1934,-5908,4753,-850,2783,1412,-734,-1961,17,1658,-4970,2034,6088,-233,-3527,5375,-5903,570,6279,2587,1883,-2337,38,1041,106,-610,1078,96,-60,3000,-546,3024,2058,-3508,1211,-5742,709,-656,4025,-3264,661,5322,1812,5942,2180,5971,4929,-3286,-1796,-6166,369,-4257,-2973,1148,295,-4406,5390,1251,5507,328,4770,3657,3264,-3168,2680,4645,-1233,-2985,7968,3820,319,3251,-2042,-783,-14296,10966,-4416,5888,2656,9765,7036,17587,56,-5053,24472,10488,-10058,-4956,4841,-13203,6958,-1781,3908,-450,2719,-7451,-3559,798,4104,612,17148,-214,2543,-5322,3066,-997,-12177,-1915,-10000,11289,-13544,-8217,-6625,8588,-7055,9311,-7382,4069,4670,3425,-2259,7553,751,1229,-11181,-1900,-1036,1882,466,-6357,-15498,7294,-13681,7231,-982,-2386,-1934,609,-4338,6674,2475,19980,3071,-9155,1394,-1459,4401,-2117,-3007,-10371,9741,18164,4162,-7045,466,-5434,-1530,4084,-6972,-15478,6499,3979,-12646,-13437,175,4274,-5893,5605,-2020,-4152,1005,-5122,2866,1228,-11376,1303,8740,2156,5048,1501,1088,9785,-4521,-6713,2338,-3791,4836,-3283,1002,3986,-623,-6103,-4296,3681,-4091,-967,-2536,-3808,-5595,3640,-4240,1940,2685,-136,486,2161,1586,12197,3535,1022,817,-4538,-12470,6079,4221,5649,-1993,-4575,10195,3586,909,-5922,-2103,8842,-639,1752,-3281,2646,731,3564,-4326,3828,-6264,-1732,361,2484,3386,3017,-4760,8164,1282,3820,-1325,-3881,11240,-874,-7519,4079,-175,119,3476,-1781,-4050,10449,-700,-2751,-1009,2883,1012,8432,-4809,7192,-4816,4462,-2595,8369,6064,2482,1269,4418,6240,6918,1445,10839,3708,10312,7666,10078,-689,-750,-1789,11728,3149,1959,-6782,9907,-1141,-5834,3811,9326,-4135,-8115,-315,5317,-5532,7451,3864,-6948,1925,635,1434,1226,2358,2668,4511,7416,7539,9438,1258,-3166,2695,8681,3737,695,-4465,9335,8291,5883,11474,2927,8989,-831,-10136,3459,-808,-10107,-4997,2602,-1439,3010,-881,681,14033,5209,-7338,5488,3205,-10429,5302,-234,-3833,148,-5605,-4726,5957,5708,5122,-3493,2408,-1986,-13886,2634,-6640,14609,-4160,-509,-1787,-9843,6967,12656,7338,-5195,1128,6093,4924,-8120,147,4660};
    Wx[41]='{1949,1076,-2386,-3083,-1027,-2474,396,1508,-463,215,-1459,118,-1297,-4768,-3164,-3325,-3471,2098,2683,-3532,715,-3950,-1061,-2600,2563,-2342,-2059,-791,-1030,3376,2663,-3198,-3881,-4223,1650,-2379,-2443,-4277,11191,6166,700,1561,-3723,-4770,-2480,1663,-9326,-2286,-5966,1146,1217,8076,2412,1551,-3449,-2034,-7,2917,-342,4919,2622,-1866,628,-2198,3623,2235,1372,-433,-3388,576,-1507,-28,-1518,-1844,-2132,-1694,1864,828,-3076,2604,690,-1257,-2885,-1436,2998,-4875,-2626,-22,6,-1303,-1870,2132,5556,1962,-1092,924,266,1595,3911,-1943,252,10361,1313,1641,4252,1334,-3183,2298,-5029,-423,-4006,-3129,3845,-8520,-15449,2220,-646,4165,-1706,-2678,1652,-5737,4333,2351,-4262,7163,4335,812,5859,7685,-1343,-1529,16181,-3757,3461,11523,-3876,-4226,16171,-6479,6757,14111,7744,-3505,-14697,-1601,-4682,4084,-6606,-3415,-1446,144,290,-6958,1213,-4763,6196,-3227,-8666,-733,2883,8911,-707,-1929,-17724,724,3952,3303,4868,2076,-13300,-12363,-5649,1597,-3222,9628,-12744,-1390,1461,5981,14970,-138,-7431,7685,-5151,9584,6655,-1663,2932,1267,-7304,-1967,-12685,-3537,2648,-1564,6811,8032,9775,-3093,-880,-2917,930,798,-30,-506,-517,-5922,1251,1878,-2988,1689,-243,-8403,-6074,-4006,5683,-3535,-2126,-374,-141,1320,-1986,-1967,6118,83,-5776,-3168,-9453,-4045,1370,-12324,-2846,-3439,-4189,3395,-2111,-445,-6904,-1284,-597,3674,3967,-1137,-5834,-6113,10205,906,-3203,938,408,-13232,880,-4047,-1634,3552,1298,-769,-1616,-9121,-521,-6723,3774,-352,4248,1557,-1876,-8759,-469,77,-6772,-4177,-2244,-2366,-915,411,5009,2490,-80,-305,-341,-2330,-971,2145,1201,-5175,-4121,-3359,-799,872,-4064,-8217,-6010,-5458,2349,2924,-6791,-2358,420,3503,7353,-1712,-8247,5493,1800,-8164,-10927,-6044,2304,9443,-9111,3696,-7490,-5322,-5390,-681,-6323,-2056,6274,-2456,4626,153,773,-1505,7495,4052,-2286,-478,-22,-5170,5234,-8300,-2675,642,5639,3024,3027,3723,-1221,5688,2729,4802,-2016,3081,-5703,-1387,5966,6953,-3264,2541,-1514,-828,13828,4599,7089,6230,818,-9824,1035,187,-2373,98,1439,3837,7788,611,2629,-6459,-29,-134,5698,-10156,2119,-1218,3684,-170,6025,-4423,640,-2198,1700,-6181,2318,-1643,-4223,-9287,-364,-7158,6665,5566,239,-2829,460,6088,-12285,802,-1128,-5117,2580,-3725};
    Wx[42]='{-1068,3452,-4758,2030,-770,1817,3779,-894,-722,-3166,-2780,727,572,-6967,-354,1269,-10195,1241,626,1856,1147,-344,-60,-1573,236,-1076,2186,-3068,-984,-2446,-1519,-8481,-1029,-5117,1319,2670,-308,1879,-543,-2797,3015,-3613,-544,-1677,5439,2127,-3637,-1882,711,129,-1141,-5522,1323,1892,-2998,-2878,-171,-2131,2541,-2453,-7006,40,4152,-1756,1062,555,1558,-8994,1437,1131,1048,1041,-2990,385,2081,-5478,-638,824,-764,-1044,-2382,-7451,-3957,-1430,3950,-4208,726,-2288,-4167,-70,-3664,713,-1135,-1618,-1938,-20,-5126,126,-1791,-6411,-989,3847,1690,2504,5864,-3012,-4741,-10761,-3063,-3952,-4355,-1914,-355,11796,10478,-4089,-2235,-2495,342,1788,3422,3918,5292,-3188,-3920,2103,-412,-8535,-6206,-1002,-1741,-1934,-22109,-10341,1757,-938,-4003,4904,-5273,-16552,-3874,-13574,-3337,1871,3007,4499,6064,-9409,-4111,687,-4936,573,10673,16855,-1981,8774,-438,1640,-381,1187,2629,9160,5429,-5249,7797,-3259,-5053,1439,-1618,-2871,1577,5605,3754,-5209,2907,-6489,7988,-14208,740,-4770,2478,-686,-4809,-5317,-1318,-3173,3911,-7592,1727,-4829,-592,-1098,-4040,4868,6313,5483,-8901,-13632,440,-22304,-668,1531,-3361,-3244,4824,-513,8203,5981,-338,-2209,-4372,1500,2968,8217,2113,-654,5947,778,-740,492,444,650,1353,-2751,5288,-3186,5307,1287,4980,-5761,1406,5385,-2205,5458,-2451,-134,-1459,1006,-6958,7475,4440,7631,8310,8779,-14560,-560,-1604,-799,-1805,635,-5117,703,-288,1397,-3115,-1890,463,627,-285,-8901,-5595,3376,1233,-2176,-3215,-3835,874,-2407,-1363,3,-3786,-208,-325,-3442,-26,-243,-2612,7485,-4145,-5048,-115,1170,-6577,351,7260,-1993,2944,729,6445,1425,4541,537,1018,1705,6718,-1514,-1462,-11718,-782,2854,-1809,6210,-6845,-1217,7285,144,7202,6523,-4370,-1934,-9501,-3869,-753,8696,-5229,-7275,6166,4052,2949,275,4907,-114,2407,-1953,8872,-3366,3149,-580,49,619,-1459,2763,-5458,777,3737,-3176,-185,4519,-235,3986,7099,-1756,3435,-624,-1437,-1955,-7963,-10000,-2861,-136,2680,-6972,4899,4750,5756,1953,3093,2238,5678,-8691,-2038,1881,-3378,537,-7309,-755,4106,914,11220,6621,-3593,3354,-1501,837,4550,-3461,515,2020,-3652,-7543,-3327,4375,-3044,-5532,-3566,1657,3115,645,-1531,-5571,431,1041,-6850,8940,3139,-5839,-2631,-1464,3308,396};
    Wx[43]='{394,-1755,-3083,-1658,-6074,-704,-5585,-2905,671,3210,-720,1778,-4360,-658,3530,-5136,-6313,-1887,-3498,-777,2416,451,-1545,-324,-3100,-3571,757,2421,-351,-1516,3168,-7709,3190,-5449,125,-2142,1164,-1523,-1577,-2131,-4184,4506,-351,3393,-615,-2663,-814,2089,-1921,-580,-545,-5664,-1575,2893,1817,-4816,1024,3896,-2968,-3220,-642,1956,-1362,-3706,-4084,1517,-847,-8916,-2011,4323,602,-1163,872,1909,171,3056,1303,4077,-1217,-221,-1470,-2663,-4748,-1278,-2519,69,-367,-1052,-354,-1245,-7651,-4692,809,-1441,-5195,-2380,-6176,1073,-1655,-271,757,-2712,1844,-6464,426,636,-4289,-14541,-812,2602,11982,8544,-4423,-5434,-21855,-7543,2376,4694,2275,-2003,2421,-809,7338,1558,-2714,1936,-2117,-5185,-7280,12812,-6972,-6782,7246,3850,-3203,-5986,-410,2248,-3225,5175,-8041,1571,-10703,10039,18281,-2802,-5698,3984,3876,-16308,11083,2612,-3210,-11181,-4987,406,5371,-1298,-3500,-2058,-7128,-3020,26035,-9082,1254,-608,3447,1024,-2141,1135,3408,-8334,2307,-11914,-3520,2849,-3425,1085,2055,3637,-5434,10566,-13300,16816,4279,-6142,-2678,-5913,-3278,188,4555,3920,-3605,-2070,-5170,-1845,-4562,3464,-6337,3913,5712,-9462,-5610,-2102,-202,-1447,3696,1116,-7719,-3449,-1768,-1133,-3569,-2941,1073,-4521,-7363,-867,-5532,-1696,2371,-125,-6347,3395,-3217,-4494,3149,-1791,-910,2452,5849,-3137,-12490,-2451,-2519,1146,2437,3300,-6948,-5209,1202,-10751,2597,-9394,-14599,1240,-2070,-3544,-1408,-5346,1024,-4472,2717,3515,787,7006,-7700,1750,-5654,3308,3337,-3071,-3891,5385,-700,-271,-1414,-5473,-1256,3559,-1833,-2188,5751,-4399,3535,-1636,-2900,-4465,-6835,2111,-1940,-6708,759,-2231,-505,-7641,548,1483,-4462,-1860,2215,2089,-1056,3190,5415,-6884,-5634,1588,2124,-3715,9550,-16845,1397,1304,-3698,31,6406,266,-2272,2734,-6005,182,-7280,-7612,612,-1972,-7666,-809,-6196,8037,9223,3022,-208,3386,3703,-1392,-737,4348,864,-1135,6113,-11923,-9931,687,3613,-2795,-2580,2634,-2304,-10712,-4228,-5800,-865,-2873,-4645,-4648,-7265,154,-606,-2619,-6186,-3488,10751,2983,5883,3483,-1527,3496,-1019,-3977,-1927,-5200,-6616,-1025,1755,4389,-3801,-12099,1939,13037,2602,2462,6689,-49,-301,-625,-4985,7246,5351,1252,550,-4123,2983,-10634,-1652,-3500,-2468,-4616,1889,6152,-2370,4609,2780,-9638,10224,-8276,-5781,-9912,2091,-7543};
    Wx[44]='{1169,5332,172,1384,-1635,606,5708,407,-478,-848,-2026,1743,-2021,-3044,-4599,-1247,-3232,-2497,-3024,767,-2446,1258,4570,-1778,1782,-469,776,-561,-1555,1287,330,-3708,4755,222,-4790,-1896,283,-670,414,-6503,-339,-3037,-2741,-6474,-4802,1932,4216,-6962,-1843,-21,7124,1376,1350,-1811,2929,2990,-2941,-540,577,-22,-66,-207,6469,-1284,1843,-428,-708,-4353,-1062,-1258,-5415,-2155,-1860,-1573,-284,-253,-104,-2856,-1110,4064,-386,-2474,-562,24,4489,-711,630,2856,4257,2087,-1730,1596,162,1739,4616,-2275,-1063,5449,-1848,-2416,1190,-6708,957,-7211,-2565,-482,-2744,-3491,-220,1936,3955,1630,3041,-6459,6259,-1124,-12519,-2236,1949,1401,1635,-83,-3791,2900,1146,-3181,-1942,-1418,-3198,-11708,3886,1850,-9741,2780,-1287,-3615,-2968,-3305,5610,4289,4838,-16826,-1965,-4921,-11298,-3898,-3447,-6943,-4082,-7685,-1198,571,-2453,6875,-2504,6450,1105,42,-4667,-1495,4140,474,6616,711,2174,-2490,-1624,9448,-566,-6513,-5024,-1480,2592,-3666,1428,-16552,-3107,2471,514,3977,-1362,-10156,2858,2746,-468,-697,-1699,1816,1544,-1887,-2900,-18925,-2430,2619,2071,-2768,2653,19052,-5908,2561,638,7934,2463,-3237,1163,110,-5576,131,-1262,869,1840,-1636,-4255,11767,-9589,6831,6323,7456,-5634,969,-556,-4892,4965,-7695,2088,5249,-2246,822,-4389,-5786,-1840,7875,5483,-2675,1262,2873,-1566,-24,5019,-3190,-2252,-2829,4355,3432,-2961,-6445,5268,1568,5747,3288,-992,4353,-1649,12861,243,5258,3955,-1213,-1329,1950,-5068,787,4003,-2622,-2324,-3271,-3430,7631,-740,1475,513,2236,736,3986,2753,11396,187,5009,2081,-1643,-309,-5976,2524,5385,1923,2486,2316,2956,-4370,1666,1678,1358,2127,4296,-1036,1798,-1232,-6059,3542,748,-1865,12958,-2766,1276,2335,1860,-4448,-9975,-5366,3850,-9824,-4257,-3176,-2053,-9790,-2229,3208,1093,-6127,1961,-5781,-1695,4133,-5708,4868,3278,-3767,1145,-3190,697,-7968,3010,-1705,-2744,-6713,1934,-1903,4465,-1125,-5917,-1281,-2368,-1621,-1181,-1396,-5185,3100,-954,4040,-9,5839,-5161,2834,5717,1015,-4726,642,-3259,3872,-2069,-10146,1372,3547,187,-856,-7651,1999,-113,1892,-7709,1296,-6210,-8388,-1262,-7172,6337,4187,28,-3706,-407,348,-3825,-4150,9672,1567,6689,-4724,8530,-1425,-3254,4108,2443,1643,3652,2353,5874,9150,-6923,2211,1666};
    Wx[45]='{-29,-5000,-3706,-3371,1628,-345,-3059,-1054,761,2893,6708,3715,1241,-464,1760,-520,835,5292,2056,-3818,937,-320,-4331,1167,-2359,2335,2430,2384,-2512,-2264,-65,-2449,-2468,937,-1029,1285,345,-296,-8950,5209,-755,2919,-104,2543,2856,-3007,662,8618,1050,-2362,-1947,-850,-55,-5234,2331,-6342,-830,-1612,2141,-1947,1857,1658,-2132,-3811,-2858,-600,-610,121,6835,3388,-997,2573,2497,1607,2165,2514,10097,12,-3505,-2797,1011,3510,-1994,2561,160,1516,157,563,-2619,-408,-1773,-2071,-184,-3417,965,3789,-3020,-1999,-1057,3918,1618,-1467,877,837,6528,-1091,2631,7065,214,-237,-773,-6264,-1296,-11113,-3881,-4841,2775,4111,3190,-5576,-2966,-5698,-128,-8710,4020,-1179,-546,5083,-3774,2016,-3051,-10732,11474,-11816,-1319,-459,6191,541,-19111,640,-4689,4064,-16083,-623,-5053,19287,13457,4721,-3933,-8935,-2279,2088,-4353,7587,-2834,-12070,-5136,4565,-3874,125,-1922,-5561,-4289,-3576,-2044,-764,2246,-3237,197,-2414,9511,-8701,-2863,10390,-1961,19990,-529,8437,14833,-7670,4257,10585,9658,-9008,-6254,-417,-3979,-6831,-3798,-1436,4108,-11044,9067,1900,9755,-7954,5688,11464,4787,-88,393,11357,-3078,998,-2279,328,-3615,5195,4587,2431,-2783,-2006,-2812,-7954,-1151,1838,4956,2504,-2578,-1006,-371,2792,-3251,4531,-1021,-2897,-4509,-1315,1201,222,-1641,-3405,3591,-1496,-7412,-5878,-222,-97,-1529,4777,-900,-1840,10732,-52,4619,-26,2176,-2812,-3298,-3640,-9462,-5644,-5327,-6064,2548,3703,-4655,-1480,-2404,3933,-5073,-6508,429,-3930,5888,-5620,-600,5610,2954,-489,-3745,-5937,2778,-4328,-6665,-955,-9858,-262,2137,-908,2476,-1422,-5698,-9912,-5292,-733,-6005,2192,797,286,4143,2305,-7143,1940,3579,-1328,988,-4487,408,1245,3002,-2709,141,-206,-2766,6132,-9033,11562,6254,-6542,-3581,-2425,3149,-9184,-9790,4797,8754,1713,-942,1856,-296,-3105,-7797,1215,-1171,3078,-2144,3415,-2709,3103,6665,235,-540,7412,5385,-7294,244,3652,934,2399,3930,675,-5122,-7060,3942,-2479,3750,2398,1270,-4040,2839,-4409,-6684,-2025,8222,-4309,3327,8164,899,2097,1235,-334,-1181,4641,-6875,914,800,-1264,25312,7036,-6640,-4465,9868,3295,-563,1087,101,2770,-204,-452,832,-2149,-2305,-19394,-4711,2464,-8247,-106,722,4367,2592,-5366,-6533,-960,-4758,-3542,-286,-251,-5209,6938};
    Wx[46]='{-582,-491,310,-1315,-1761,2119,1201,1461,113,-1035,490,-865,1442,3713,-3476,-1486,-1977,2252,-1729,2822,2895,2298,-569,547,-410,-1931,2792,1302,-36,365,3041,5761,4975,2626,3718,-1322,-2553,401,-1651,-1013,503,2624,2263,-2395,1070,4001,3984,-4643,-269,-2937,3825,4155,3640,4382,-1402,-11152,3229,5361,-106,-901,-2031,2044,-933,1958,1217,-382,2497,3073,-1006,-1900,-1420,944,4748,3471,-205,5195,4130,3256,-2673,3942,1112,4301,16,4174,541,5063,-14,2509,1765,4003,-1068,4357,-814,3916,169,-3386,-2275,3830,2229,-6010,-2861,-9453,-726,3666,1928,-38,616,1343,-21,-2951,-4313,3562,7348,-2438,6025,-836,8256,3115,530,1878,2395,1003,2043,-4550,-3127,1197,944,6230,-13496,-1781,1080,12246,8134,12070,221,773,1489,-1481,-5234,-14628,549,6835,-14550,-5253,-5625,-3669,-13496,10351,-6088,-3142,-7460,-7978,5102,-5424,-373,-14160,1502,-7031,-2900,-2910,-863,-3928,-8710,-2369,14541,-1505,-2161,7734,1247,-7485,-8969,2885,3623,-15117,1934,-1555,-14335,-906,-5776,-3229,2305,6801,-1802,-1794,3867,-11474,1090,10126,-55,4575,-2115,-9448,266,-70,-7265,1063,-2093,9370,-3833,2344,-787,4978,1069,-41,1657,-1533,-6450,-2086,-1949,2780,-4013,-689,-2337,4130,-8413,-1616,-4838,397,-1040,-1223,1560,-2133,-1547,-4660,-2056,-3959,-1148,85,-2607,-4589,-6630,-5170,-569,-415,-2465,-3806,1873,1170,-1665,-1617,1297,-8916,-4421,1295,3398,1679,-9086,-1563,-1663,1151,-6435,7021,1254,4570,394,5151,-2288,654,-2988,4511,-2299,-6274,2514,-1550,-3759,3066,858,-4238,934,-3334,4699,2170,1644,-1520,1682,-1021,3395,3984,1059,2519,1955,-496,7309,-8779,-660,-4777,-2893,2239,-5297,3195,-4152,3198,-5234,-643,2519,4567,2744,751,168,2678,8198,7016,-194,-2534,-3103,4348,2717,-1198,5595,-928,-3005,-1378,-735,4335,-3586,-2885,-3625,-2402,1436,-1157,3310,-2553,-2197,-2666,-54,-2900,-1623,1635,-3835,3359,-2277,967,-3999,427,-5771,-1551,-3955,-6635,-6137,-2072,567,-1745,-285,-2301,-949,626,5644,481,2105,-3386,-643,4768,4882,2670,-11435,-6191,-57,-5932,-2011,-630,-5170,-2775,3947,1385,-3974,-5009,7055,5688,-11074,-5468,4812,4562,-2534,-4279,-3896,3515,563,-962,1938,2661,3928,3034,-2868,6401,-833,-1069,-1586,-2524,-6284,6191,-7275,-4248,-1145,7133,9829,4223,1922,2687,946,2702};
    Wx[47]='{-2420,-7260,-2692,1049,-1883,1707,-4045,-6572,1113,-996,242,-4003,-8618,-3469,-4599,-5517,-9838,-2347,-5815,-623,76,-1933,-549,-4348,-2949,-4174,-7954,-6572,-8334,2661,-1965,-7153,-3776,736,-7338,-4580,-3566,88,-2543,-2122,-4118,2213,-3930,-2357,577,-4960,202,-5810,-624,-955,-8427,4345,5092,-2536,2430,-17998,-2001,-2211,-2639,-6503,-7817,-4726,-2121,-2819,-1405,-1677,-2553,-4123,503,1087,-1479,-1306,-844,-286,3261,-4501,-8974,1585,799,-8671,-4406,-4899,-3867,-1296,1630,-8925,2097,-2949,-3825,858,-449,-8442,-5722,2309,-7451,-6210,-8159,-4687,-4816,-5947,5107,-5219,-1606,3806,-2868,-1563,-5229,125,-4191,5346,3850,2597,-2460,0,17861,-9770,-6699,2773,-873,292,-815,938,7436,-334,-4807,61,-6723,1390,4572,1082,1093,-4746,-966,-963,-2221,-12402,-4458,-2863,-5517,11230,6064,-1029,-2546,-13583,-2459,5820,-10429,2822,-5395,-5830,-551,-870,-5322,13535,-1944,-3295,2507,-262,-2226,-5791,2534,-15322,-7656,1741,1738,-1611,-89,13320,-3496,740,4416,4045,6250,-15224,6967,-12792,936,-6972,14667,1983,-1245,-2697,16552,-6484,5952,-7968,-6547,-6069,-149,-439,-7602,2148,5034,3020,-17548,-12968,-3471,-16591,-12636,-810,-652,4003,-2587,-2666,-1735,2052,-6411,5581,2827,-1937,-11,-1206,3359,1351,-2883,3986,1425,-4382,-2384,-443,-2032,-2736,1312,-1395,1870,-817,6069,241,1057,-4465,-2492,973,5327,-3488,4575,-3757,4670,-293,-592,7109,-629,3586,4157,2055,6137,13525,5654,545,1232,2712,5673,3566,825,1230,-424,8037,-53,1331,-135,1661,-2792,1123,3054,-1329,-10449,5009,265,6621,2283,6635,-3444,3652,-2016,1898,922,-53,1497,2521,4260,-747,-306,1218,453,5180,7695,-1427,-994,2734,3293,846,2517,8583,3867,8027,-5073,180,2084,-4609,696,334,3872,4699,3469,312,-1276,-1026,-2376,4943,-3928,-1103,-9858,-6782,-1311,-1328,5561,3793,-834,-12578,-3012,-5678,7758,1379,-6411,-13437,4521,-3645,-4113,-1636,-5004,-1956,-3022,991,1776,5434,-1221,-1997,-2971,6152,4775,-1778,-3918,-2012,-922,5263,4909,4040,-4760,-162,8281,-3410,1341,2463,5693,416,5063,-4548,8178,-190,-3916,-12421,-1606,-2236,8593,-3679,-7158,8437,-4265,4470,7939,399,-560,-7685,-12041,-4326,1335,-6860,-6660,-1002,-1745,-8959,-2915,4987,-8403,2065,-1744,2360,-2768,-859,-1168,-1343,-3745,-1696,-1901,9550,10527,3850,-2053,1135,-1619,-8354};
    Wx[48]='{-537,-2158,2563,398,-1657,-793,2030,-173,-2357,-2795,3591,593,3439,2617,57,9716,-2098,-3781,-1480,-2888,916,1032,503,-848,3044,-294,2188,788,-346,-1281,-385,-2751,6850,1406,2285,-562,4228,3059,-778,-1458,-869,-1089,6762,1450,338,2978,10429,1583,-1158,2375,-1004,3803,-956,-957,-1113,6665,-109,-1561,297,-1408,2963,5356,4863,3710,6762,-1590,2844,-1025,-2609,-2944,3779,2321,3483,1665,-891,1110,6962,1740,-1204,-219,1613,8076,1997,1759,-7641,1614,-1697,318,-1433,-515,-50,331,3496,2138,5791,-2658,1794,1979,2770,1072,7250,-2208,820,-118,2114,322,-6855,2568,-4792,432,6962,-1395,5571,8027,-3273,513,425,5092,1517,-500,1867,1511,-4716,-5820,-649,5346,-610,3,-9589,-6147,4221,9116,-2,-7836,-6489,-112,1353,5366,5742,-8085,940,-13232,5317,-7294,-13388,-10615,-7333,-1766,-5629,4094,3886,3701,-1730,-2697,1683,4992,-1669,2963,-5107,-1372,-6074,9482,-3569,5439,-10878,81,-5991,7929,-258,283,-3041,-5659,2580,1986,-1400,8652,9384,-574,10917,-3034,-3188,-4230,1168,2790,-7460,-22929,7597,12265,1862,817,-1983,-3630,4182,5297,-6079,-68,-4672,3542,2479,-13134,-1553,-8208,-1669,-1668,1667,-93,-4809,-12197,364,-459,-6015,-80,-2661,-3950,-3901,-8588,4934,-8325,3708,-1590,1006,-880,-1658,-2575,-6406,-2639,-596,-2275,-4399,-5927,-5688,-8525,-8227,-10478,-8842,3593,1566,-1546,456,-2288,-3881,-2692,-7426,-9326,-10390,1701,7983,-4384,-541,-3432,3103,-2183,-4709,-5405,-5200,-1512,4265,-2309,-4929,5581,88,-4284,-690,3854,-13457,-3195,-1799,-2060,408,-4653,-3801,6010,2592,-429,-2568,-7158,7861,-10498,-8281,2592,2968,4108,-8598,-3417,-1689,-1317,-3225,-3830,7500,2495,117,-3959,-6596,6440,3586,-4731,-7045,-6186,-8955,-10410,-1098,1762,161,5893,-1033,-12968,-83,-4714,1583,2534,4736,452,2396,348,-6713,-1106,-1051,2176,5380,-1734,-7402,-520,4711,-305,4396,5590,-3525,-4716,-473,-4375,1794,1582,104,1227,-2678,3833,-5708,-2829,-4101,-6660,6547,-1156,886,4721,-5981,1894,-7065,-4824,-2883,6567,5717,-7216,-5683,81,-9135,502,8139,-3032,4057,234,-87,973,7246,-3647,-139,-7622,-422,-3107,-5185,-6191,3693,7475,2095,1333,-2381,-3603,1505,3076,-3732,358,-1535,4975,-5029,-606,-14785,4055,-11884,88,3208,-4355,7080,-35,-2978,9819,10927,-6376,-1503,-13271,-2666,-3691};
    Wx[49]='{145,9926,-215,-316,2229,-1645,-361,-175,-143,4741,12080,5556,-3552,-2841,-1688,-3129,1463,6220,-1087,-2753,3732,4167,-1826,2729,974,-2868,400,-849,1645,335,-2054,1309,4785,4567,-4411,3264,-5517,-3769,1169,-349,1903,5805,-6308,5083,-6181,485,1987,7026,1844,-994,1052,952,2103,182,4782,1894,8037,4455,4074,-2810,-747,1311,-4338,-191,1743,-1391,4174,1694,745,4025,-1529,-45,-4499,739,-192,-761,-129,1092,-2238,177,3518,5317,3620,3110,4633,5361,-1098,1287,-695,-222,1049,6005,-659,-1842,4648,1010,-3808,4208,841,2340,-1419,14179,2207,4750,-1925,1610,-1205,-5678,-850,-7651,2668,-4389,-5249,14082,16582,909,4672,-8159,2646,2290,-1678,-1097,-4003,1062,-2152,1401,-1093,-4069,-1458,-2100,-481,-3959,17861,-9291,-1370,529,8208,2452,-1600,12001,456,858,-18623,-172,15253,5043,12578,9150,-1091,226,3972,-2415,7749,5488,4133,-10517,12412,1149,-206,446,3693,6523,-9555,-3664,8608,-2514,3110,-10234,-2141,-49,706,-15859,-5903,-1522,-558,-5053,-4919,5825,-3701,1336,497,1680,-4479,-2531,-2270,-10625,2875,-4321,-4321,-2291,-975,-5566,-10732,-1422,5825,-8764,-3974,678,4174,-2675,-3398,9731,-2012,838,-2215,-158,6718,-759,1224,6826,-6318,-168,1560,-2646,-3825,1241,-502,1511,-1345,2595,1445,-1657,-1000,-4294,3129,-3918,-2778,1055,-990,1896,-3242,-4775,-5859,1475,-4335,-2025,-1571,-4836,-7231,-914,-4501,-5258,1437,10673,11357,897,1462,-4714,-3049,-418,-11992,-7338,2261,4504,-2619,-4702,-5429,-1046,-938,7475,162,-6079,2944,-8935,58,1762,1329,10048,-1843,5195,1666,-2609,-2493,-1623,-163,-4375,-7446,-7275,1304,-127,-1499,2883,1682,-2795,-750,-6684,1142,-3012,-978,-2059,-1141,-624,-3994,-2607,-5585,-730,375,-9438,4489,1372,-4404,9023,4050,-4970,-7636,5878,3666,1765,9057,4787,-2169,4042,386,2724,492,4099,12363,-7509,-3808,-831,9980,-4709,-3266,1145,-527,22,1114,2340,1163,2878,-2279,6982,-3522,2636,165,-4436,6025,4245,-2017,-6577,5200,-487,172,-1247,-3759,1038,16132,-3066,-2059,-3063,-603,1658,-4914,-1328,-114,3476,3374,4978,5024,3271,3093,-1013,-254,1356,-1087,2619,4672,1849,6166,8798,7133,1314,4792,-66,4387,1331,1647,-4667,-1708,4741,1058,7197,3630,-5161,9277,-3376,4721,-6459,-59,-1774,2218,-3149,-4548,7949,-4064,971,-6821,13779,2685,6059};
    Wx[50]='{-8,5322,-4401,2883,2114,941,5688,5224,1192,2961,10195,-2517,5620,1824,-2866,-1058,4118,2137,-853,1126,-2476,-126,1749,214,1844,1560,-208,-800,-622,1145,-2770,5048,-4086,-569,-1245,4462,4770,1791,-2861,188,2795,-447,-242,-3125,-1821,4433,7187,12832,419,-731,33,-619,2073,739,1550,2580,-2032,-5463,1552,-6308,-5346,369,-2498,1032,-3547,3278,961,-974,-157,-1851,4099,3066,-4946,2364,357,-2169,3818,4025,1150,5839,-171,7792,-3352,5156,2453,1325,599,-1324,-1094,4160,3090,327,2285,-52,4653,3361,5390,3464,1052,2407,-2670,4145,1856,-6083,-1932,2529,-1340,-318,-328,-2478,-194,-1538,-3969,-3164,11845,2963,11396,1953,4985,2641,-154,-4672,875,-7563,1507,-4938,775,-2778,-2047,-8720,3986,-2946,-5283,14785,5166,6030,-698,5053,2778,-7631,3161,-979,-7636,-1512,-5000,-7304,11601,-5961,1330,-4008,8330,1578,4792,11640,-3352,3176,-6660,3166,3283,4426,-2254,728,8212,-6655,-12978,531,-2058,12792,525,-2370,3796,11279,59,-9804,1878,-1750,458,8569,2885,3178,-2744,8032,-3603,-5986,4770,-2934,2958,-3864,5664,2307,-5761,-7377,-3981,2087,10234,1159,-902,17031,-1223,-5068,-228,-21074,-2324,787,-5571,455,3208,-1663,2286,343,-4873,4975,-1083,2893,5771,-6318,8305,4365,-302,5869,-2033,-1023,2880,-1658,2393,3496,5458,1784,1525,-4399,1842,-2778,-111,3430,-1754,6313,-5590,55,-8603,50,892,5961,5439,7861,7524,878,-3952,-697,-434,1180,-1512,-2062,-2836,8417,1248,1159,3212,-4816,1430,1038,-3728,4479,5317,-892,-5947,-572,-2685,-3740,-1221,-1791,7919,-5195,1061,-1455,1406,1871,-933,6650,5991,6923,-5092,-12636,2451,554,4584,-6748,1279,-814,1781,6215,-1927,-4306,3872,-5375,7587,-2308,1132,-27,2406,2707,354,-3330,-6987,3308,-6567,-377,149,-755,446,-16,3571,2973,-140,3742,4880,-3598,1677,14423,-740,2631,-798,2093,2111,3364,191,509,-942,4028,635,-2166,-603,1028,9399,4814,3505,1707,3588,-3547,-2047,3874,-1857,12236,961,4770,6040,1441,-3112,664,-1922,886,-1975,-3676,1522,4504,928,-858,1673,-8208,1091,7368,-1285,1994,500,-1705,4589,4797,-5913,1147,5219,-1345,4445,1883,1262,10039,1240,-8256,-1389,10117,378,-5356,-3244,-2391,-7656,4013,8657,501,2012,-6474,-1802,7954,2697,6967,859,-5512,8759,-9301,6289,-908,1508,5786};
    Wx[51]='{362,-661,112,-1336,-1534,-1273,2604,899,-311,-1596,9018,1429,-3205,1763,1442,-5639,-1306,932,-664,-1667,132,-1317,108,-2081,3662,-1251,-255,-1227,2995,2517,3166,3605,2687,-2448,2205,5239,-717,370,-6513,1981,-446,1838,1115,971,1108,-1662,11923,2697,-508,-1452,1278,382,1270,-1884,-1379,3562,2568,4467,3750,797,-236,-1434,1411,2403,1553,3049,-583,10429,169,493,-2137,2359,-4494,3657,-714,-4516,-1566,-94,-877,3354,-1456,10410,4277,10341,-1745,-472,2534,644,2269,-23,-1553,2839,-809,2827,2156,1024,-260,391,-1029,-483,1132,11718,2873,-679,-7167,910,2290,-2167,3854,-8476,9233,3781,-781,7465,7387,-12919,-6259,-3513,-7792,258,-4143,3547,1938,7119,1224,-8447,4916,1657,5874,-2341,115,8715,-9785,2293,548,4414,7524,1230,-5844,7490,-2283,-1834,-11230,6240,-10068,11728,-952,-4033,-5791,4846,10634,3940,4794,-3229,4843,3312,14648,742,7490,-1091,262,5668,3405,-1876,15771,-3684,-749,10458,228,-904,-12773,-2709,-20,-12734,2775,11611,-1320,2491,-15175,5468,-734,17412,-1202,-398,-5107,-8959,101,-7646,-640,1673,-3063,1572,-4626,1728,-4543,2432,3002,-6381,-4973,2004,891,-982,1824,4897,252,-1589,3166,-1441,412,1387,-3215,1949,-2281,-4460,-117,-2402,3691,4328,1533,2036,3139,-2756,-3537,-3955,4301,2517,5029,-886,-3254,3205,-890,-542,6430,3295,5351,-3552,2358,2983,-1622,-3806,579,-10156,-6611,5102,-9418,-5239,-14482,3125,-2080,-1793,637,1978,5839,-12197,-8173,-7783,-2871,3686,313,-913,280,5996,-619,-5869,7133,114,3518,1990,-2152,-56,4851,928,-5317,-7207,-33,6591,420,6196,-4543,-1383,1043,2915,-270,-1588,4978,-2683,3081,6738,-3688,1844,4812,718,2741,258,-4,-2917,-2617,13310,-2492,2741,2437,-1945,-8115,-643,-372,-622,1755,-2089,2430,-5454,-244,-1350,-864,-2310,3291,-1666,6191,1418,1262,2932,9741,-2131,-1173,1424,9184,-339,5976,4262,3571,2010,-4138,2382,7519,2778,3591,-3186,1152,7788,1279,-4052,1020,-3754,-2583,565,-4326,-9199,3422,858,-6196,-2648,-478,-1951,-5073,-2709,-2347,-1368,-1907,-8334,5302,-962,-4414,-2807,7055,-3669,770,8037,89,-110,-3408,11337,-2314,-1159,5917,-687,4162,3632,7397,384,-6635,1114,3684,379,1003,50,12636,-8525,9433,-1159,-3146,-3500,7514,6401,-4,17177,2243,-469,6083,9375,2551,-3002};
    Wx[52]='{-1489,1262,-2768,-1322,1990,-26,-5673,-7514,-2502,-2702,-2851,2541,-2114,-2399,-3547,-1708,459,-2854,145,1162,4914,-626,-1444,0,767,-1756,2150,887,2797,1683,410,4375,-295,2351,-4116,-3049,-2412,3471,2897,-1290,-1018,-1817,2492,2133,2198,3691,4279,-8540,-1051,895,-4697,4777,1979,1334,1883,2003,481,-367,-1577,2543,5029,-4904,4003,-1323,-4379,-2349,-2509,-1842,253,-18,-1000,-292,7177,-3415,2380,-1668,5600,1303,1914,534,-1373,446,1910,-1531,3881,346,2153,3476,-3049,1038,-4841,-8559,-4536,4729,-91,-208,-1052,-2873,-53,-1253,-1950,-2199,1093,-4421,5361,475,5991,-12822,165,-3657,-2692,-2922,277,-11718,5097,-16582,-11845,5961,4067,3217,3635,-4245,6171,-2602,-949,4294,-8652,-624,-14580,6748,-185,5014,-13242,5209,-2355,-2170,-5131,4089,6318,-5712,935,-1734,7836,903,7324,-7597,-15644,-8120,4252,1257,-3679,4809,6269,-5039,5659,-2381,9086,-2653,6035,-4416,-6772,-16376,6030,-6469,7958,2125,-664,-7524,-1627,3642,4138,288,1962,19667,390,-306,-10517,9985,-2116,5883,-10458,-9370,4333,14560,9916,-5830,-1347,6660,2502,-1790,15107,10595,378,1867,-11806,9082,-9687,-8168,-6718,-3132,-3107,-13564,-2590,35,-158,1296,-4401,-1220,-1300,-2039,-8710,427,251,501,2346,-4042,-181,-1558,-1878,-445,-21,1524,-7114,4672,-2937,-4531,1511,-673,961,-2966,788,-1503,-2985,-7431,-1205,2739,498,1716,-202,-6997,2680,-3823,3752,-5922,-199,-4887,3388,-1234,-1396,-3764,-2170,-8085,-2182,-2249,-3708,-5092,-971,2724,-6323,-183,256,125,-156,4978,-10136,-4699,-2060,-9311,-3332,-755,4777,622,6225,214,1408,2915,-2785,-5683,-2624,3120,-565,3400,5092,1903,-3286,2731,2341,-3034,-734,-1916,-606,1933,-1868,2131,-9501,1424,-2636,-3449,-1206,-5063,-2177,-143,-207,1726,1182,-559,-254,3381,-4399,-1651,-1551,-1915,-3366,-1566,-4550,-5185,-8613,7622,-7421,354,7080,4033,-5161,-2990,4223,-4724,-3269,-3771,-106,-1796,291,2266,-10458,-10146,4138,4667,1319,3547,-10048,-10878,-5517,-10185,7089,-4326,1469,-4763,-4650,6005,1307,4240,-9951,-7773,2724,1655,-826,-663,-1237,5463,-4365,-2556,2697,-7265,-3459,-4697,-12021,-316,-10146,1569,-847,-11113,-3876,-6650,4504,-5043,-1580,4892,-5595,-1671,2517,-2075,1610,-5439,-1137,331,2438,-6152,-4858,-7504,-5478,3813,1531,7080,-5693,-5346,-2340,6015,-194,-8144,-5449,-1710};
    Wx[53]='{117,2116,-330,-1658,1151,-2064,-4123,-3442,1547,455,-5747,-922,-1849,1729,1118,-7744,3833,3190,-503,1308,1293,1194,974,1538,0,-1531,1596,-1490,-3002,-3256,-376,-1127,2941,3300,-3781,3112,1282,-2093,-4396,3608,1751,2712,1437,-3347,-900,368,-3522,-759,1525,-3039,-820,897,1721,-2807,405,8823,-128,3493,411,3291,79,-2032,-675,1964,-2934,2258,-1136,-4909,3215,745,-6918,-8247,4416,-2683,-2851,495,12236,-1370,-3781,1462,-2432,-5893,-856,2878,3725,4555,-1781,-1386,-2498,-1407,-5649,-948,-137,1158,-954,-1262,2047,-939,2126,4260,2045,20371,3244,-2000,4428,3349,-1502,5126,1995,15,-5043,-3083,14,-2194,9394,-2707,-7910,-3251,388,-2758,-4,1650,143,4064,-187,-769,2088,6284,-23984,3640,-244,12099,-6840,16572,-535,-3251,-2990,3500,-5117,-4592,-1843,-17880,-13066,6215,11806,-771,373,2448,10507,14677,-11845,-3120,11240,7031,-2519,-1541,7011,25,2186,1034,3845,7070,-8691,-2758,8139,-1495,-2427,6762,1502,130,2012,-4877,-2568,2222,-6376,17900,1334,-388,6567,-3791,327,-5131,-5717,3071,-9213,-1,4533,-20449,2075,-702,3305,-2954,-4001,1216,3994,8530,-1754,-6152,7963,-23867,-3295,-2332,-1627,-1126,-3166,-1444,5498,1282,-3081,378,-3806,3659,-1849,1685,9663,-7236,-10058,4650,668,1213,3046,953,-1128,-916,-3049,816,-1213,1839,-535,1243,-6777,2451,9755,7773,6372,-2509,-299,2741,3669,2685,-1,7216,-4797,4094,9912,-1810,7060,6982,-2080,7905,-10683,1646,6860,513,2792,-2497,3771,4394,340,-4594,634,2302,830,-4050,15380,3481,2319,-1953,-709,1845,3439,1490,2734,53,-2077,3386,-4338,2902,1713,-5883,861,3640,-2712,5664,2110,-8564,-3991,4858,-3942,3486,3347,-276,-969,5903,7050,5332,7207,-12822,3769,3864,65,-392,-10429,2272,-3005,-3203,-481,6513,-2091,-6821,-4772,2012,-5893,3034,4182,-3930,2089,6127,3305,6611,6181,930,-7890,304,-6816,-2142,-352,4299,2521,8798,-2344,3881,871,5942,6176,-2958,8188,3891,1944,676,4953,3330,-3110,-9589,3801,-1453,7729,8476,-3791,-1657,1329,508,-7949,-281,-3430,-273,4279,1464,-265,1901,1258,-1579,7866,-3168,-6347,-4536,-319,-1086,-5976,-2230,-1357,-3352,7016,-1553,-2222,4248,4162,5415,-4750,2089,-1495,5341,-2595,-1920,-10136,1734,-7954,6381,-676,9868,2187,-470,-5664,-4499,-2756,1905,4604,3586,5874,5283};
    Wx[54]='{-2885,-5112,-1523,3850,225,-3244,1015,404,-3740,1507,-3132,-1119,-3059,2944,-3444,-2553,6269,1665,1030,-177,1083,1724,4492,899,3398,4597,2052,-997,1361,1887,-1149,-829,-3085,623,1937,255,-1185,-1683,-5771,3107,891,-1448,-3945,-1188,2095,583,-8173,841,2609,-1191,9956,-1624,5351,2125,2597,7358,-2478,478,979,8935,-513,2238,2780,2800,-327,1420,-976,-834,-1322,-980,-4125,2012,1932,1888,1107,-2105,-1734,243,-6357,-2673,-268,4682,-3920,-6147,2316,-6147,97,-1247,3796,2344,228,-3295,877,-1589,-2932,-1759,9033,-3754,-911,3681,-399,-4475,2124,521,-8208,827,-8789,-5292,5546,196,-9790,6567,-6928,2009,4086,12412,9799,-633,4770,4914,-2095,4814,-820,-3105,657,-116,-3215,1026,11464,3571,2489,10117,-4765,-3669,2705,-4174,878,4250,8642,-11181,4814,-6806,146,-2792,-17460,-6899,7314,-13886,8217,-3103,5595,16035,10087,3925,-4912,4704,8530,-1726,-10253,-1044,964,1412,17753,7377,2211,468,2022,-18701,2368,-3066,4746,4401,7114,-8789,-3395,-1058,2648,1032,13808,-3127,-4240,137,-1987,-14375,2149,-6323,2445,-1303,4816,1359,-6181,441,-3891,2257,1210,3383,4343,-1370,-3393,12089,2543,-2524,-1263,-9018,-2447,-1098,-964,-1506,3408,-2556,-4526,2199,2646,5283,4704,-6459,-10771,-1226,-3710,-382,976,2352,-2602,-2795,-3752,-399,2427,-3137,-4743,5170,734,1239,2111,-8803,-5810,-4472,-3642,-2883,-2070,2736,742,7929,-3122,-3483,1293,-9213,-6660,1057,1462,7216,-3720,-4409,4089,-5361,3796,1547,-4362,2536,-2590,48,-560,-1922,-5385,1137,-520,-191,-2683,-4929,588,-3142,14,-5664,-2756,-3295,-1821,-6865,-3935,-2360,1986,-2490,-535,-9160,-71,-2053,-293,-9062,1843,5112,-4802,4067,-4660,-12519,-5688,4594,-6259,-5239,2690,1396,3266,-2374,2083,836,-41,-5556,-3510,-694,3830,2812,292,-10957,-9848,3615,-901,6928,2135,-2500,-1973,3200,-5566,-4042,-5058,3056,1931,428,-1546,-2861,2149,-6918,3535,1907,1911,2239,3627,-7636,248,-2773,-3239,-5527,1497,9057,1049,5541,-2089,-7304,6679,-4172,-4020,-4812,-1844,363,-826,-9970,1206,-5034,2824,1361,-4260,-5942,1256,-1027,-1359,780,-382,719,-2271,5126,-6684,-5869,6586,-5336,1506,-8110,3090,3115,-5424,-133,-1333,-3420,-897,-3403,-3220,-829,3366,-4228,4086,-4565,5537,4680,2624,6630,-3256,1386,758,-5683,-3974,-1279,8349,3979,-2778,-560};
    Wx[55]='{-334,-960,667,1856,-2719,-3935,1132,-3737,927,2570,4230,201,-242,-4494,449,2421,-2973,-1025,-2373,233,-2131,137,-3686,-62,-1538,-812,-5224,-2000,-5722,-1093,-128,-3627,-936,-1689,-5937,5981,-5151,-2585,-7397,-2993,1186,-3281,314,-505,-1839,224,6733,-4650,-1939,-1557,-2458,-1502,-3498,2937,2893,-3955,-100,1845,3332,-464,-3830,-3657,-3537,-4824,-83,1712,-1644,-5693,-5058,-2155,60,-1015,-2238,-3571,-2462,-3576,-5737,-3867,-2238,-2080,1113,4077,2934,-4775,-6181,679,-102,397,720,1647,-1572,-1170,-260,-3315,-1579,-3022,-2802,-1028,-4841,-2578,718,15283,-1741,-1215,-5517,1927,-3745,9248,-6577,-5810,14033,5332,-1012,-15068,5668,9096,-6416,796,2690,-375,-928,-2135,2100,-3464,1965,1973,6376,5229,687,-1022,884,582,-7099,4245,3049,3527,1242,2321,1927,-5214,4025,616,-137,3107,-15576,-3151,5483,-1811,526,-6474,1971,-8198,-12119,9272,-7246,6835,3881,423,-8310,1172,2995,15117,946,-1478,-8461,-1654,-2213,-138,1232,156,898,-5205,-2705,-5405,-2012,3674,1264,1644,13564,8906,6000,6816,-3952,-1605,-79,15517,-3769,-2648,-521,376,-1574,-5502,-4577,-2061,804,-14941,2160,-2293,1318,4208,1922,7368,-1759,1084,1129,-1697,4147,8403,-2988,-1956,1918,-2624,-718,-7358,2917,-1787,1519,1566,-2006,784,-2541,-3527,-828,-793,5527,-1209,3408,-1492,2479,1890,-2476,6782,-2438,2966,3659,3654,-2171,910,3574,8652,-4077,-6225,-253,-5185,-2310,-617,2934,5034,-2407,3559,2971,3181,-6845,1983,-778,8686,5332,-653,680,-5878,589,-9516,5786,5009,8056,3891,-2404,18378,-480,1466,-4853,883,-2624,-2766,-1461,2047,3315,-1680,1004,-593,-289,2587,-4226,7607,3740,4555,-955,3637,-5039,895,-2285,42,-3471,-3540,9936,4455,-4050,8105,-1871,5727,-496,-2174,-5864,-1938,1167,-2861,-2900,1352,-4580,2270,-6416,-3361,6347,-1483,1994,-1518,3793,-5112,3188,4160,2166,-3930,-3708,3334,2592,494,-2758,-488,-10839,-1870,-401,5898,924,-471,-5380,3547,2381,1827,3896,2121,-1723,-189,-7729,-2280,-2287,5693,12529,96,-1518,1239,-1514,1229,-9487,-572,-571,9067,2687,1538,5507,1439,-4453,-5126,1783,2897,1190,9096,1850,2788,447,3239,2038,1541,-6015,858,-2915,2215,3408,-4382,-6982,3300,-4562,2834,-2158,-1715,-10732,8339,-3295,7885,429,-5390,1511,5454,-3029,-9658,693,2006,-4602,7763,-5000,1170};
    Wx[56]='{-4067,6372,1017,2,-1558,739,-2320,7436,-746,-2919,-4890,-1329,3691,-4963,-4714,4206,-7753,-5166,2213,-369,2558,1186,-2480,-3369,1412,1511,-374,2252,-1936,1417,2185,2281,2100,-2763,3266,-1378,5795,669,2087,-6225,4509,-7172,1838,2265,8686,-697,2810,-1519,896,-1959,4301,1293,-4401,795,1517,-1816,2558,2431,-5205,4794,-1856,-142,3796,0,6157,-3420,1505,-689,-4235,-2841,-1619,-8105,2180,-5219,2254,1906,-11250,2929,4326,-2902,-1417,-5644,1466,-2100,979,5737,-853,1153,5507,965,4089,2174,-2386,-1314,4670,3818,784,-8466,-4401,621,1439,-18535,-5083,-3503,-170,-1322,7700,-8056,-3576,-1101,1748,-564,4543,604,11074,9902,-6787,-18,-1212,-1706,668,2897,15322,5009,-497,2316,-7817,1702,9311,7104,-292,12021,-905,-13789,4409,-8217,-1016,324,622,2069,3452,-10742,1672,9365,14169,-9326,-5253,2983,-6499,-1034,-744,-13974,-4296,-4125,54,9370,3972,-1364,-2066,2556,3918,5258,-7700,1523,7875,1634,-1365,-6166,2165,264,8242,1601,-3779,191,-246,2115,-788,14697,290,9428,1017,14160,-12031,3227,303,15966,4047,132,-1667,330,3391,-348,8002,1734,-1440,461,-9589,-17500,-9775,6142,1041,840,4638,-245,3549,-1680,4116,7539,1976,-3984,374,-1810,-74,1982,-80,3664,1464,436,-2995,568,-385,1872,864,4521,2084,-183,-1182,-4311,-1064,2312,-1065,-3486,6123,-7368,-837,-2905,-2690,2423,-6020,-3569,2484,-1656,2442,-1206,-11435,-6914,-4252,4465,5439,-1224,2108,-2159,-914,-8051,2932,2824,-1196,2163,-1157,-4025,2070,9814,19,4401,6020,-4216,714,15927,-2346,-1451,-993,3564,-3364,-1311,6362,8388,-3608,-8286,4179,2183,969,-6450,4006,2609,1162,-1800,2211,-835,277,-233,6455,2371,5517,2205,13447,1385,-1392,4458,4582,8466,1472,-2797,243,-6162,7944,12646,-117,4511,2191,2481,-9970,-5234,-1815,4680,6596,-9741,662,-14228,1402,-855,5175,-1238,-128,-1441,2888,-2749,128,-8339,-1207,-132,-3300,-3967,10273,-12509,1939,-4958,-1072,6430,-2379,-11464,-2081,-3679,-3623,3010,269,-7187,1549,-1353,3881,-663,3811,-1071,-252,-3684,166,7060,-1794,6611,-2683,-2373,-1585,-2058,-423,-4240,-2406,3996,299,-2274,10947,3583,-8720,1052,450,-11757,5380,-399,-437,-9355,-3142,-2578,8129,-1793,-3837,3083,616,-4980,1093,121,3342,235,4396,-9765,-570,6596,7470,7612,180,7841,2067,3090};
    Wx[57]='{-2132,-4680,71,863,760,9,841,1237,-1582,-282,-8784,-1182,2602,-1617,7524,-7084,-1363,-3073,-2213,-3540,-2166,3894,841,-3566,1799,1828,-2624,-2138,-6206,3410,397,-4047,141,-1872,1202,3222,-848,6240,2446,230,-1715,-675,1948,1481,-2115,188,9819,2447,-1155,-1561,-1076,2188,-1313,3957,-715,744,-2316,-5009,2255,-1639,-3889,-5458,8354,-2426,-4421,-1462,-1939,-8276,-2164,1162,1622,-1685,-3093,5205,581,3518,-2080,187,3496,452,-1795,-867,1250,-3049,-2817,-6660,1405,-1596,-946,-727,2915,1910,761,-5708,-8583,-300,2089,617,-2958,3002,287,-5600,722,4707,-3686,-411,-9067,-7309,-181,1767,10029,1340,-3310,9926,-10771,-4101,-3701,2432,-285,-2617,-723,3889,-5214,-1320,1470,-3415,3203,2156,-4096,-13593,4667,4858,-4018,3427,-4604,4045,-3554,2922,-9570,-1571,6635,-6586,-1555,7109,-3254,2495,-2335,-4516,-6313,-688,14189,-7788,1756,4499,1499,16035,-10419,2534,-1796,-897,5034,-4841,-6284,-932,6806,63,5195,-5346,-1274,-959,196,-4479,2156,-14902,559,-4357,-7353,-2185,4401,-526,4033,-12216,-5468,-4350,915,10146,-1639,7880,-4848,1860,-3591,-3408,-6464,-1324,-4841,2758,3725,12578,-781,-8754,-484,-8906,-2536,-6489,-1416,704,-1998,3957,2841,-1276,-3498,10,3015,-6518,-295,220,-1596,-3764,1748,2108,-443,-2775,955,-2949,-5454,-86,2147,625,10908,-3479,1291,3801,-1173,1483,-4064,13,2702,5419,3830,-3295,3908,-2829,689,-2058,8022,4238,8598,-667,-3049,-5854,-3100,33,-704,1751,-1145,276,-3981,-4233,-5551,-273,911,-691,-2465,4216,-662,3000,3854,34,-332,2420,-3747,3505,-10224,-7119,-903,1180,10244,-4797,2563,363,2038,1787,-2183,7187,134,-5136,1077,1417,-1859,-980,41,-4506,-7421,-3684,-9799,-4484,2617,-3215,150,-6142,-30,3610,7568,2580,-2714,-1405,-683,-3525,-4809,304,-14677,4440,4389,2524,4958,-5014,2546,-681,4455,-6669,867,-2418,3405,-690,-2106,-4409,2849,-2749,1148,5732,845,1154,8925,2866,6630,1593,-1557,1870,4360,-3701,4755,-1383,-4111,9521,5981,4125,-9326,-5073,2927,-115,11240,257,2208,5991,-556,-1110,-5551,-4689,-1036,919,1885,-1324,553,-212,386,4453,1507,-254,811,-3918,1248,-3740,-9614,-3129,-762,-3864,1975,135,6337,66,-296,8486,-679,10693,-2932,-3232,-1678,8491,375,700,3320,6352,-7006,-5278,345,-336,3195,-8422,-5336,2863};
    Wx[58]='{-912,-7055,1208,-1329,-1910,-1749,4938,4689,-2121,3974,-1154,4016,3452,1095,3041,2116,-1583,2152,4072,1871,-1608,2563,-78,-804,-2580,2548,2124,953,739,-3046,-3666,2408,-1912,661,-791,1536,-3269,4133,6,-1420,4560,148,1138,1080,9257,2927,1479,3549,4565,-606,8432,4882,700,1577,-355,65,4348,4665,3300,3166,-2402,352,9697,2301,2259,2143,-813,7294,-685,-471,517,-2631,-2352,-247,-314,446,3586,-2980,273,3508,2023,272,1998,-263,-5102,3366,-1838,-424,-359,5375,1281,2276,4316,-3684,-330,1538,-1716,-4279,858,2128,-1436,-136,1391,-336,3395,-41,-6616,7553,3630,715,-1190,-1246,2619,6479,2229,6821,-11259,-3388,164,-1380,-143,5039,3320,8310,4526,2807,7802,821,-5327,-3710,6728,-1091,-5229,5043,-746,13085,-4797,1871,-15810,3835,442,9379,9013,13740,27832,-13037,11728,5136,2900,-2841,1441,-15244,1929,-258,-5400,4152,-2365,-4108,6015,4765,2805,13925,-5366,5131,-240,869,526,11093,5004,-1898,-5937,-7978,-2033,-1712,1995,-5249,1235,-7690,-11064,3276,-7485,-5527,-14453,-3569,-2080,4165,2932,3449,-1986,6123,-591,-14013,-8608,-2578,-7666,7265,2333,-5419,2110,10351,661,-7436,1770,1469,80,-1645,2080,-3906,2531,2436,-864,-207,-2575,-6064,1078,-7773,2156,-1207,2198,6147,-1468,-2331,78,-1608,-223,-3002,-602,1267,1463,2922,13,-4362,-5390,-2536,-1485,6713,-1850,2592,-5639,-5107,-4660,-8969,-2033,6254,-3291,-1705,-14853,-6054,-1126,-4497,-7534,-6538,2172,-1511,1715,-3403,-3652,2360,954,-7270,2902,-2978,-3947,-85,4106,3759,-4230,-6669,-3085,-6616,2517,-406,-6196,-3366,-650,-3945,-8066,-4616,3979,305,-2216,-1638,-4399,-5092,-3037,950,404,-1203,725,2966,6674,-1453,-5776,-8110,1873,-116,-549,-6606,5800,-1791,-1142,1888,-1260,-5747,-1232,-1846,9257,-6210,-1120,7597,2983,6445,5048,-506,444,-4826,8886,4580,9912,7065,-8432,-6894,462,4228,-6235,-1430,1192,-8198,5825,4523,-712,-3571,-5385,-3735,1986,4960,-5922,-4670,-14101,-2656,4626,-2553,-2656,5483,-3974,1904,-2695,4279,-8178,-167,6416,2128,-6254,-6547,-661,-4355,-7167,3312,-195,1787,3234,3715,-2069,3181,-508,-8198,1329,-5620,-3352,-1872,-1717,532,-54,-1726,3513,-2392,-3789,1163,3303,5166,-728,2531,1906,1661,-7216,-5507,-32,3237,1248,6909,11269,-2087,-1956,12324,-3339,-6025,-8471,-1613,2058,3081};
    Wx[59]='{-1990,-8383,-4753,682,296,398,2171,-2347,-740,2670,-1413,858,-2491,245,1243,-4548,11953,4902,3640,-1254,746,-1566,-2680,-2086,-2449,-962,2517,1026,-2141,-3566,-2409,-5761,536,-3962,-8164,4135,-2154,-3383,-3225,-198,-2475,-9570,-4570,289,138,-2476,-4335,3100,-1300,-1396,-2651,-1649,-181,-1169,-3781,-5854,-3552,5000,1680,-3034,-7763,8759,-3413,-2033,-875,5234,132,-7055,-1353,3532,20,-9931,727,-7329,-78,-2083,5532,-449,731,2215,5986,-1239,1407,-4453,-1506,318,-662,-2673,-34,-2895,913,-4702,-1833,4013,-2459,-3811,1741,-5229,7143,-759,-3547,10625,3166,5522,7597,455,-4047,-996,3430,-2424,-9702,-6982,2700,12216,1210,9765,845,-6801,2038,-4663,1220,-5747,1262,4274,-5971,-2775,5820,4907,-10498,-3229,-3212,-618,4155,-10781,-2229,2595,-4055,2648,-4299,-1560,-3750,5273,-10332,13095,1665,569,692,4675,823,-9570,-3508,-7299,-10224,3408,-7124,-8,7851,368,2565,-3964,-617,4670,9775,-5317,-2430,-4140,-2036,1307,5922,735,-1124,-9936,-6352,6923,-759,11201,13144,10927,5566,-1816,9726,4433,-8046,-13964,-8886,-5556,2924,-2729,-5244,-253,-10810,4936,-8574,2233,16767,-6582,4694,431,6347,-8676,-1087,1942,-2824,5302,-394,1376,8398,2197,351,10107,5776,2117,-2343,3544,5122,61,-4033,7236,-1268,-363,1671,35,-3188,-7133,-29,2268,-2741,3449,4699,-10039,-507,5971,4187,9116,2408,1588,-3078,-1490,-827,2890,-1079,-3183,5844,449,38,-1134,-4655,461,-8037,2196,-9702,4206,2727,6230,3364,2583,2493,809,2988,6376,720,-3525,4194,-2380,-6503,3269,358,1291,834,4206,-31,7363,-3110,-2746,-1654,-3869,1232,-1237,7939,232,-933,-6513,-621,1071,-7934,5405,-5673,2783,1102,-22,-2768,-4902,4865,1470,9809,6230,-1951,-542,1413,7807,-7250,944,1452,1013,-3300,-6127,12871,-2062,1611,7001,-2089,3061,-7348,11826,-2127,4221,8881,7333,11572,-939,-1484,-678,-2474,-1507,-9633,2607,4296,1064,-761,-287,3105,-1501,-4309,3676,-5009,1264,3464,-1050,-2998,8041,3708,1806,-462,9204,-755,7241,1461,9370,-9550,-1945,6362,5878,3547,1893,7998,1579,899,-4755,5712,569,-3403,5693,-2680,827,-2692,-4545,11318,399,-5781,5927,471,3605,2592,-989,12031,-2454,-2072,3674,-1779,-154,3059,9252,5864,1138,-11357,-1614,-4072,2312,-5585,967,-141,-4123,-5131,14951,-698,-723,476,3933,4318,7216};
    Wx[60]='{784,-1481,2177,1282,-458,-2575,-1320,-2836,4060,3269,5385,807,-2496,6435,-3925,1126,-6489,242,1693,545,489,-3681,-5859,1672,-2272,-1125,1768,193,1824,1054,-2156,-2369,1262,-141,-1932,1982,-2700,1755,-2073,-2220,-1842,-3225,-3327,1231,-1827,2583,2270,-480,938,-1405,-1033,-4113,-5141,-4030,5341,-2264,-1006,5937,-2073,-5800,3850,-1063,-8945,-142,-676,3415,-367,-3957,-46,1555,-4030,-7656,1245,-1298,-736,-1010,-1373,-4025,-4855,-3796,-510,555,-5810,-2031,-3110,-9648,-3125,3051,1345,3293,-2233,1921,-2390,-4138,-6391,-2305,-2442,-4182,3945,-3911,-1043,13798,-3088,-3403,-1001,4990,5297,1369,-2467,811,430,7275,-721,7475,9565,11406,-3757,4108,-1271,1878,-1121,-1892,-423,9770,4313,-5131,-2358,-1483,-1842,-4357,7026,-10654,-32,1593,-4943,-2109,5146,-387,-2326,8413,-4130,20625,-1213,4570,11386,-13115,4584,6875,-6455,1547,-7353,835,5180,-6538,-3989,-7177,-789,-3757,6528,6342,-181,5039,-18603,-4582,10468,1412,-2805,-12275,698,-2851,7299,1683,-5131,4509,60,14960,4440,-1754,-7104,-883,-1618,5024,8378,12636,-5234,-3024,2421,4438,-646,-1778,-3586,-10195,401,-99,22539,-6572,-4318,9750,7333,-12861,-822,6323,4353,1749,99,-2370,5175,5595,-8076,2141,5683,-2418,367,8173,-4301,5639,-200,7470,1243,-80,4614,57,-2081,1090,811,-354,-2476,1157,1815,3024,-3244,1210,-673,3647,-2565,1801,-5288,-1694,10917,6542,1966,2052,2041,-2846,3269,1917,-13671,-7353,2442,2917,3686,1455,-639,773,2561,-2322,897,4670,-6308,5976,4250,3662,2546,5610,-1434,921,-968,-125,3498,817,4572,2448,3771,4645,-2492,9116,8354,1872,1885,-8227,-4633,279,447,-2154,-3195,4609,-3215,-4523,-5312,-1357,-4294,7460,9633,-3786,7602,1342,-1757,-778,-393,-1990,-2070,-5942,3295,115,-1745,-12255,2524,-4555,3344,5156,11005,-1014,898,3637,-1719,5581,1043,3837,-12294,498,-3098,-2086,-7622,4348,-2363,3208,3022,3583,-2915,892,-1160,-5151,-11425,-29,5605,5317,1777,-1497,-3852,2678,976,4880,931,6640,1203,4567,-1152,-1337,-13408,-132,4333,3471,-6191,-3837,4938,10244,-3093,10087,-1105,651,-661,-3298,-2137,7890,1304,-1781,-2766,3215,-507,-7006,-5639,-128,901,2851,-86,2514,2541,-92,827,-2420,1095,6889,2447,-8579,-7485,774,-2108,-457,458,1088,1981,4570,1212,-2846,-3798,83,-8168,2802,5888,-3779};
    Wx[61]='{1846,-3222,1066,1682,-1350,972,-3073,-2454,-8085,1235,1353,-765,-603,-2304,-584,4721,3012,-1729,-4743,1927,585,-924,-1295,-4272,1904,-315,-3056,2761,330,3598,4794,-5439,4309,805,2656,-991,544,-2512,5668,4704,2105,3227,3608,-465,7553,2695,-5473,1574,-4375,937,-2235,-2066,1782,5053,-520,567,3500,2320,-115,-54,-2832,186,-575,1050,2683,-2888,-2369,1392,989,299,-1927,8598,-5800,996,-1467,-5405,2438,407,75,-2575,-2030,-7416,2243,-3254,-1289,-2800,288,3728,-1021,-1001,-1013,-1273,158,1520,809,11,2113,7929,419,-88,-2980,11718,-2291,1051,-3388,-200,-5766,-12001,841,-834,12636,1801,5898,7299,1102,4006,9101,2015,2225,3701,-989,5410,-3291,2663,-5981,4072,-900,-9106,7988,-7031,1610,-6196,1429,5800,-680,-2335,1160,3049,-11621,1160,-4372,-8427,-6420,-13007,1416,673,-6674,4160,-2171,-10908,15498,-495,7329,1501,227,975,9858,2199,-1461,-7509,1165,4636,1817,-3139,6865,-2932,-1090,5932,-466,847,-6782,-6962,284,-18818,-3815,-17041,-8554,4641,328,-3127,-3671,9809,2888,3342,-2692,5952,-1159,10644,3610,-1656,-1253,6381,-14404,-1735,-6362,4836,-2481,-1807,950,9946,310,-7299,170,-5029,-2093,-1106,856,-4174,-1915,-4333,-4033,1607,-2839,-4992,-2517,-9370,3378,-7729,-4272,1624,1566,813,-1844,-7719,-5419,-4406,-3549,-379,-11523,298,-930,-6455,-1474,-8325,1055,-3515,-5234,812,-5458,-3137,-4780,11210,-8945,3522,-734,-1596,-1873,-3500,640,-2912,-11582,-1895,-2,-2880,-6088,932,-5112,-4514,3381,-5361,-9,-5717,-4091,-4128,-11503,-3928,-148,-4082,-306,-1832,-2580,7968,-1373,-4824,-3979,-11416,-657,-6538,-6772,-1751,-3291,56,-276,-1013,1633,-3789,-1839,-5151,1667,-902,5825,-679,-11494,1170,-1846,858,-1254,-10781,-5058,-2700,7998,-575,-4431,-3850,-6054,-438,-4738,9838,758,-138,-2401,-3122,4636,-211,-2670,2416,1899,2102,-5112,2338,3447,-257,3918,-1943,1220,-684,-6323,3808,2423,-106,4765,434,-336,-136,-1373,-4816,2773,2722,-706,913,-4533,1943,9985,5498,708,910,1091,-3684,-7182,526,-1524,-11035,386,-269,-4392,3767,-3635,-8779,20,2305,-3408,-834,-1070,7231,-779,-14443,-3127,205,-3549,-1497,1154,5454,-4885,-9291,-4763,-7431,4689,-5981,-1280,-793,-4897,-4523,-6503,-4746,-5463,6113,-272,-1512,-879,-4372,-3928,149,-8095,8725,3771,-1857,-786,-8662,-3940,-163};
    Wx[62]='{1567,6640,-4350,-4843,932,1246,3288,-3261,1307,729,429,-1517,737,-4445,3046,-3073,-1122,1180,545,2418,704,1232,-3110,-2263,-1026,-961,793,225,3203,-794,681,-1866,3020,2983,-803,-4836,-718,-1904,-3825,-2414,260,2683,5532,-2658,-2978,-1303,-7412,-4294,-6923,-3056,-4753,7822,1441,520,363,-5175,-7216,1184,2565,-1724,-2366,-59,-1655,-1643,2758,1690,3310,-2379,-4467,-984,1885,-7622,-1634,6074,87,-188,-12255,-1319,-2451,-4621,-975,-13466,-3395,-5708,5449,3764,2020,-1414,-623,1920,1390,-623,-1547,-1353,-2702,1740,1585,-667,-6396,70,4995,15273,3959,-3007,-1268,-1975,-5019,11210,3349,-47,536,-4113,246,12792,842,-1555,20761,2509,-3178,456,-2073,-6049,10185,-2304,955,-2318,-3315,-4589,17871,-1923,2277,-1422,3474,-1635,653,381,3571,-11025,1762,4565,15751,-1473,5039,-794,8750,3981,-4626,-3444,1613,11992,2312,14384,19033,2770,6240,-642,13388,-307,9541,-2106,4155,-2077,-3076,-332,880,4792,-1414,-11513,-4389,-1447,-7636,440,-3327,426,4165,-12939,-9780,1033,-19765,-5136,3105,10097,-7895,1474,2846,1756,368,-9287,-810,2403,-789,394,-14121,-1137,-8627,-10566,1909,-7675,-4265,-17519,4499,3356,-1596,-4807,-757,2302,4770,4016,397,-2944,-9008,5942,-1939,-1499,-5541,2277,1285,-1035,1049,303,513,-578,561,-4614,-3117,-1494,-6953,2111,3571,-3942,-5024,-8144,9418,3198,-3862,-4453,2229,288,787,700,991,-7968,-1582,-543,1182,1865,7788,-6513,2697,-661,1484,-2188,5107,-1287,-1862,2895,6215,3666,-12519,-243,-4621,-4411,-2239,-7407,1831,-1398,2976,338,-3291,971,-5278,-1354,905,-3378,1644,839,-3828,2954,-1551,-6635,590,152,4545,2539,-654,-4846,-320,-111,-1589,4750,6347,3798,-1212,1994,424,-227,-3256,1730,5083,1845,3352,2687,-7822,-1378,-5078,9716,1137,-4584,-3098,-797,-15390,131,808,-8266,3728,-1967,-256,-4970,-3879,-14394,-627,223,-5703,-5776,-272,-1263,-3115,5288,-1790,-2521,-4821,-14140,3510,-1413,-1779,-6821,-2314,7475,-1807,-1807,-3198,-11210,-2729,552,-2810,-3579,-1685,-9125,142,1932,-1549,235,-3388,-1965,-4633,-8154,-2469,-2059,-9130,-4602,1778,-6948,-2155,-457,1871,5722,3999,-1280,5786,-8916,-4987,-12021,802,-7412,-71,-2700,-12177,-12314,-648,-3427,1063,-8066,-11113,2983,5302,-5229,393,-2929,4523,1016,3598,2468,-3251,2346,-596,4211,3759,5375,-1552,-2939};
    Wx[63]='{1256,2656,51,-3034,2639,3413,-2587,2415,-919,-751,2502,-1591,32,-1087,-1894,-278,-4631,-505,-1406,-996,-3186,-4201,-3618,-6215,-832,-5556,1789,-944,-1595,153,750,-5537,-3420,-1408,2348,-588,1052,-3847,-1865,1892,-1605,1119,-2188,-1385,-1496,2303,-7924,95,-5361,553,-7939,1402,-3061,1579,1096,2673,-962,-957,2077,-6713,-821,3002,-6757,-3459,-4890,-3610,-2819,2568,-451,1069,-567,-798,4345,-1708,1216,-2995,-6933,-971,-901,-972,1320,-3369,-3823,-2739,2648,-164,918,1890,2159,-3093,-681,-3618,-6840,4721,-4938,-9584,3254,3732,-2230,-5791,4948,4746,-1161,-3886,-85,-1381,-2434,-1311,-2912,-575,15644,192,892,-2966,-13603,-5747,8261,83,-2712,-1962,-1662,-2204,3520,2512,-8920,-5092,2012,2165,6958,-1777,304,-4755,10830,5322,-3859,4025,-2259,-4643,17109,-7592,6479,2061,5854,-3488,-17919,-601,-23808,6489,-5078,5180,-2980,-14208,-544,3798,2824,-5053,8613,985,-17167,-3725,-6811,4030,1121,-3693,-1348,-1740,192,6352,2183,2995,-2089,-6777,-2070,-4272,-504,-603,-11035,-33,12636,2391,8466,-9062,-10234,12255,6088,-15214,-1876,6914,1168,1441,-3618,9296,-4353,3376,-9921,-6074,4724,4270,-3623,-9594,60,-5175,275,1291,1541,79,-4572,-5000,-1933,-1921,-1713,-2060,-3234,2795,851,8505,13017,-3510,1646,-502,-1868,-2773,2414,-162,-3527,-957,-9028,-75,527,1077,335,-4965,-4514,-3498,10273,-5253,1837,-1175,-7153,1600,1540,6210,-5043,-7822,2878,8798,4028,600,-2524,1257,13496,576,-2800,-8481,-3869,-8168,1765,3107,-10292,2475,1791,-1091,2541,2064,-11650,1367,581,547,2279,1252,5678,2027,1302,-2301,2059,5703,4680,1749,2534,6064,2631,-2023,4824,-989,993,5424,-898,1414,-2166,2371,-720,4912,4172,9619,-99,3720,3078,-1168,-6547,438,10087,4143,6582,3994,4731,6372,-4826,-2761,1350,1162,-5649,1071,-3864,-3640,-872,-3366,-403,-7558,-2329,-7851,-4694,-1249,-2756,-7397,-2183,1704,-8818,3022,-1265,-4711,-786,-6875,5000,-2001,-1934,-1552,-2399,-2731,-5415,-4968,-1485,-538,-3251,-1237,-2524,5688,-2983,-672,1540,-1580,-3383,-2412,-900,748,-125,-4182,6870,-5981,-5908,-899,-2973,248,-4055,3188,4768,-3869,2624,-7836,5019,-5981,5502,-2480,237,-2331,-439,-49,-1246,-5971,-4233,3310,1348,-3535,-5014,-206,-754,6352,-760,-460,1024,-4670,-2282,1124,-838,21445,21250,-1763,5820,-1065,-6684,-186};
    Wx[64]='{894,5019,-1356,-1984,-650,1312,5263,339,-4267,-242,-4074,-4704,-8369,-1722,1329,-5527,-4982,-1105,-552,283,-622,-3083,-5205,59,-3757,4404,845,-1023,-1706,26,-921,5966,-5527,-1209,-6489,2639,1859,1205,-122,665,66,763,6811,3161,-4575,-4230,1400,-2641,-2827,-1992,-712,5791,-2431,2084,-1821,-4548,-1490,2268,1893,-6108,-5112,1372,-3002,-1794,3903,-3210,-152,-1436,-395,-219,-2797,2941,-5913,222,-1688,-3483,-4870,-3093,-1077,584,-1330,7514,4130,4074,-855,-9023,-3344,-3256,-5014,-662,426,5825,-4848,4345,-5615,-693,592,-4394,-3552,-3723,802,6547,2541,-7294,3376,-643,-7265,-2512,7172,-4643,-11318,-474,-9350,215,5410,4072,3920,2204,-1450,-141,527,453,8100,5971,-2086,-206,-213,2331,6791,-14570,5087,21562,-934,1237,364,4892,9067,8916,-6176,21777,-7329,5566,6499,-15654,6899,12333,3369,-1816,-1959,-2180,16044,-13408,-364,-4619,2174,-657,-4187,-3974,8159,-4782,-4521,14091,9301,12578,-18212,2075,-2858,1474,-3127,2252,-656,5537,1483,3366,2281,-4389,-6801,-443,7104,8750,-2067,-14628,3583,-4938,-47,8032,3984,11933,9863,2211,-2775,180,3369,2344,-6733,-2551,4309,-6884,1142,12988,-445,-7680,-983,4199,-2578,1359,-1580,-2374,-553,-2919,4848,4143,-397,4255,819,9990,11621,2949,2321,-231,304,-838,-622,-2104,1695,5751,2543,1578,5966,-9755,2375,5551,7866,-1605,1514,1677,-988,3686,3562,-794,3376,6953,5048,-7358,4338,3801,2028,950,-4934,-3305,6074,-5,2622,2327,1937,-2451,1848,7446,-5649,8569,1334,8984,-549,-3386,-1307,-1844,3056,-207,2049,2524,6225,-2309,-3071,-1693,1773,2971,11826,10566,-3012,919,-4016,3630,4243,-468,-3024,8706,-1315,2171,-1157,-514,-4597,4084,958,1337,-2064,-6655,349,2939,1400,4873,-6357,508,1739,8247,624,6674,6948,-5771,-2624,-3461,288,979,-2270,12695,7563,5043,1408,2670,-3015,-9355,8457,-1549,-2447,-301,-4201,3527,4086,529,2155,-5932,-3308,-3493,910,7314,-5092,5976,-3249,2729,3908,-924,-6992,7485,939,2180,1361,-4108,-1678,-3830,-1914,2038,3256,4975,8017,160,1040,-1340,1193,-723,-4455,-4406,-3320,-737,-4001,939,-1912,-4453,5502,8789,-64,5874,-617,-1771,1673,1638,-5122,3029,12001,219,-338,-2371,-3706,2768,-2106,3383,-2890,9321,-4460,90,-2641,-9418,1154,-962,1516,5219,-725,-4123,4536,-1147,-1868,6123};
    Wx[65]='{171,-2905,-655,4196,1851,3647,308,-1613,1400,-90,2282,847,1962,5888,-301,-2434,6835,2391,-2170,-1197,267,165,523,1500,-3522,-2460,1785,-3715,-1606,-1342,-996,240,-3837,3725,3774,788,1614,-4,3991,-925,745,1834,-2607,121,5595,-584,7026,-1795,121,3,-2512,3251,-142,2861,-2717,-6313,3334,87,-921,-2915,-2839,-2181,3359,1002,4091,-3435,375,-1417,2438,-2692,1964,3112,368,158,-2131,5097,6665,3957,3493,994,1485,9511,1322,7792,-2344,-307,-414,317,738,-2768,-202,-1834,-427,-125,937,-2692,-560,9135,-288,4501,1306,1162,-2370,-1955,-1424,-5317,-7880,-5693,930,-4335,-8950,-10712,4577,5869,9228,-9589,6650,5805,241,1600,2061,-6630,-3188,-7636,-1962,2583,-1116,-1774,-2814,-2406,76,-7177,1203,12919,960,-6049,8422,-3366,-294,-7309,-71,-13652,-7153,-8515,-15087,-6250,6796,-580,-3403,-2131,-811,8789,-842,-12597,2604,-9086,-5942,2060,4995,-2036,-2509,-2861,-11533,666,-6020,5473,-1001,-384,-2929,-304,5708,7280,3200,2646,1038,11386,6567,-6435,2692,-6645,-3188,1004,-145,1065,-1256,5502,3869,-1069,-1770,701,-495,-11005,5371,2442,-14599,-5434,-864,5517,-1166,-7934,594,-5380,-312,948,-2358,803,-7724,-10937,-2368,-1556,4287,-1059,-1939,-3117,1895,5854,-207,3969,5327,-3200,805,-1204,224,1743,385,-3195,1760,1632,-2154,3149,-2066,1713,100,-564,-6284,572,-1552,-3010,671,2403,3649,-8793,-6269,-2260,-7495,479,8037,3017,2912,-333,-3210,2164,-2529,-195,-4382,-3808,5278,-3913,2421,3134,2514,-704,2072,-9770,-13281,-3913,1898,7363,1928,-1602,-5332,1928,3718,-894,-2763,-5258,-2263,-8720,-2216,-623,-2619,368,5371,-3159,2176,-3139,-985,-5776,-6240,-1234,2536,-5375,-4602,2309,4724,2587,160,-2944,-3405,-3503,3520,3039,5234,4675,-4895,2851,2619,3417,-6127,-8618,5458,-651,-5864,2117,-2617,4233,-4853,11171,787,1145,-4226,-1154,3195,-2690,-458,-2707,-5874,-2678,-5947,1970,-15,6909,-14628,394,-4157,-3706,4130,-2993,2044,-195,-640,-6528,4887,-2299,-2052,-1420,2778,4458,6406,3486,-2810,-5527,1287,-337,-2135,-3271,6147,14130,-902,6308,1003,-2266,3352,-4831,555,-2753,-7641,4401,-338,-8251,-2178,3547,950,-1739,-4069,-5463,-12890,-3063,-2004,-6269,1295,200,3039,2512,1572,2437,-1345,-4338,-3142,3317,-1257,-8251,-2700,5327,4235,1427,4589,712,-11181,-4589};
    Wx[66]='{1850,-1746,-1229,-2398,3195,-1928,-4069,-83,2237,4680,1414,-2573,664,-8422,6215,-1937,6220,-3051,887,979,118,5419,4050,2602,751,-3247,1854,-1845,-120,-4995,964,-5839,-944,3754,1647,3251,1499,1571,-5380,-4458,451,2073,2386,3090,1119,-5659,5815,-886,1716,-1325,-1262,651,992,-20,6445,4514,458,-2296,2302,3752,1768,23,2507,3291,1649,2375,-417,-7333,313,-2521,-214,-3457,1247,-5297,2315,642,-4899,-3537,-423,-1525,-1205,1835,2875,1910,2729,-3750,2963,2232,1342,-51,-1849,-852,-2005,-4711,8134,884,-2076,-4741,-1979,-2941,4804,4948,849,7099,11503,-968,830,-4067,-7050,-583,-12421,-858,1013,-10419,-1694,-6293,-11318,4604,-3232,-1856,-512,2469,3000,-1143,-453,-216,-2376,-1066,916,2890,-3737,-24121,-10957,-2175,1430,3249,725,-758,10156,1000,242,5834,5083,4580,1066,9375,-3835,-6396,7011,6318,-9155,-1036,3173,908,3244,9916,5043,3305,-3217,2792,-376,1760,-2834,-6118,-398,-1169,5952,-7612,1783,2866,-786,8305,5371,-4006,844,12148,-5019,1051,925,4775,-5991,-4274,-2385,-16240,-980,-20859,-228,-1448,-5214,-547,-3391,10371,4575,-1776,-12949,1505,2281,-11162,-3769,-1511,1866,-766,-4909,1864,4133,-897,943,-6215,2988,2763,-6298,-2849,1412,1771,5063,-1810,-4104,-7832,-527,-3435,-1307,163,361,-2224,-303,-5639,-2371,-1949,6147,5903,3012,-1446,2558,-4121,6386,773,955,-1262,-7626,3771,383,5371,-5346,2271,2922,-188,-2888,352,883,-4514,1248,-7055,848,3300,-5571,-7709,1179,-3420,-6679,-5644,5849,60,-2326,4062,-626,513,-2221,10722,-3205,-3605,6196,-6035,-950,-5102,115,-4851,-9116,-6953,-5043,5375,-4216,-11582,-1217,-4802,-1542,-11503,-556,1033,5859,-2238,3686,-5605,269,-2055,-4216,686,7841,-544,4499,-3093,2880,-2900,175,-2893,2883,895,-2680,1300,1490,3781,-8671,-541,6108,-190,-148,949,1977,-8745,9912,485,4855,2663,-1203,-1678,4101,-9389,-1403,879,-4072,849,-1014,-506,-1091,-3764,133,4758,6083,8095,-9003,-4655,6474,-912,-1032,-7490,-588,-2739,8647,29,1950,-1719,-4921,856,-9047,-2054,1306,-1022,2739,-668,-993,-1641,1413,-1389,2583,5776,-9946,3220,-8935,585,7324,-7294,241,-10253,2476,-2644,3752,7338,-6132,-698,467,8447,-3217,-2736,2032,-14062,-4335,-13339,48,502,1710,4035,3518,-9023,-476,-10283,-4274,-4011,4672,8032,616,-528};
    Wx[67]='{-890,304,-2296,-1171,243,233,-1962,-3945,-1751,-2924,-2452,107,-1882,-1562,1619,-1007,-438,-4174,-5327,1624,2739,2517,1652,-1056,-1649,2448,-4184,193,68,471,930,-4204,316,0,-5800,-1230,-2277,466,1264,-1379,-236,4035,3457,-3732,2934,130,4055,484,1849,897,-1542,3112,2575,196,2136,4296,3664,-2071,-1232,-1171,-1008,6137,1533,-3327,-3134,558,598,-5043,733,2387,6616,4458,-2136,-1926,-3532,-2519,-5468,1292,3789,-5737,-4465,3461,-446,-3166,1481,-2763,1072,2368,466,3647,-1915,823,-681,486,-2629,-742,-256,3845,-1733,-2180,-2039,2365,-2912,9926,2685,-2248,-192,-10556,2434,4577,2150,956,-953,-107,-3745,2248,-10634,4521,-796,1682,1533,-2570,1260,-175,-509,946,-975,-3476,-3962,3842,2196,1161,-1058,7890,-1479,-12080,-1245,3276,-20566,-6704,-5141,-6416,-9541,-6103,1225,5483,-14423,3598,-5087,-3325,10839,-10419,5576,4284,589,1802,3098,-3093,4621,-844,-4279,5668,8940,-3830,12890,101,984,-14277,-887,-11,-11777,5395,4755,-5405,-103,5244,-4660,-2194,317,1346,-2415,-6533,-4250,7905,3059,-3725,-1962,2403,-4660,1582,3193,-19707,9423,-888,-13583,8627,-8442,-3684,-4257,652,1115,-7666,-619,-2590,2661,457,-1644,-632,-5761,-1505,-3605,-708,285,4460,-2305,-132,3876,3325,3090,-2653,2519,-3103,332,1751,-2379,-2978,4978,-435,-3664,-9594,1441,358,567,-4311,4118,-4418,5883,1309,-7973,-1812,2070,-1000,-3105,283,7954,700,-1545,-321,68,-3881,-3032,-12753,4091,-3454,311,-7553,-7519,1961,-1103,1582,-1428,-7788,-5029,-498,524,-3881,-258,6093,4682,-1094,-1401,1477,1987,-2032,-593,8784,-4077,309,-6362,1385,-1074,-6118,2956,3002,594,-3889,2170,959,-1544,-1472,2963,5380,-1473,2048,-7373,-5620,1218,614,2191,-4743,5693,-1785,7968,-1301,4245,6665,-1478,-1602,-8823,-2949,-8886,-518,2519,7543,-934,-812,-2121,1658,-5625,-2946,4973,-1665,-3381,352,-2297,-434,-4606,-558,-6889,-1925,51,-4118,-840,-5942,-13798,-4187,-5512,891,-6718,-13242,1805,-1693,-1106,1181,4536,-2486,-9492,2076,9814,-2663,924,-3186,10390,-1542,8164,5395,-6357,4938,1170,-1359,-2880,-3937,-5771,-1374,-2529,7568,-2500,7910,-1428,-5546,37,-2531,-7602,-5444,-4504,-2758,-5639,3974,-5654,-1021,-949,1728,5449,-2719,1645,1833,3325,-399,-2364,7153,-1842,6884,-7622,-6967,3801,-1981,-339,-1480,-147,-6254};
    Wx[68]='{1229,-4042,-192,-2424,938,-953,5932,4494,1971,2152,2734,-1038,5410,-541,4338,5981,5458,440,308,-2775,-348,-366,1042,80,1077,2086,3100,589,4086,-562,1580,5541,6591,5766,1374,-4477,5473,-3122,734,1667,3120,14,2707,1257,-2844,4052,5922,5107,4675,2795,2773,1492,2290,363,-125,5585,1351,1479,3017,4951,363,787,-1564,750,14462,297,1716,4660,-196,-2043,-1494,6904,3806,-5864,1242,487,1018,3090,-185,1668,326,1907,1071,6401,1145,3879,-811,315,-920,2998,3525,-530,-3781,2973,5590,-455,1740,4838,3293,6499,344,6577,2780,-5317,-9218,344,-1826,3825,-1381,3054,-5053,-2756,2797,-16162,-883,-1257,-13330,5126,-122,236,-855,-3293,-1428,-3208,443,-2739,-4377,-302,-1734,3010,125,-1326,6684,-3662,1734,-3403,-3408,123,17324,12363,-1063,-15546,4282,2551,4877,-3769,482,-249,10703,-5532,-16025,33,-2054,-9741,-998,3640,3977,357,692,4040,-5371,711,2454,-4008,-4394,-701,4353,-3127,2724,-2270,5512,1944,-681,-7211,-659,-10458,8657,-3566,1052,4755,-4411,-2934,13574,-698,-1346,-7124,-1300,-5878,-792,-3979,-7353,-2729,13662,157,-2441,4392,227,18300,-5004,12578,969,-5273,936,-582,-2427,-416,-3540,-3659,-1232,-698,-2946,1739,-5678,583,-1160,-6875,-1079,-2386,-1301,469,-1882,-274,-5751,7397,1601,-709,5209,2749,3518,-7416,5756,-63,4020,-5493,-3693,-1352,-3906,-2271,-1124,-7602,1212,162,158,848,-9599,-7416,-10048,-131,3798,-930,-354,-8691,1739,-4291,-1713,-8325,-624,128,-1536,-7329,3234,5786,-3869,70,2514,-1199,841,-1273,-888,-3627,-6645,-6503,2399,969,1516,-1937,-5747,2624,-2507,-1666,-1367,-4331,-413,-7421,404,-691,708,1386,6743,2238,2426,1406,6103,4201,7275,-889,-1171,-3159,-4807,883,3847,-859,2529,2435,-1170,-1635,-3234,-4104,6879,-2250,6694,2043,666,-2788,-3098,1407,529,2509,1707,1531,-9697,3420,-1787,3054,7094,588,4753,-3188,6499,-7519,-584,2470,5195,628,-7900,-1824,-978,-5585,1111,3251,-586,1353,6044,-3674,77,-3522,-11611,3244,-621,-1163,-1030,-4584,5830,-456,-4753,4060,6713,-571,4804,-7055,-1441,2600,-4553,1353,3413,4970,3483,1330,12666,-4060,-1495,-8896,3522,3259,2749,-2369,6440,4274,-7973,-373,-2209,201,4184,-9399,2607,-1271,2836,-2971,1097,-4853,6840,-671,4367,-3791,1270,-1185,3120,1445,3933,-3515};
    Wx[69]='{-1447,-2595,1517,-339,-855,-330,427,-1160,-2905,-2519,-7836,-125,-437,6538,-2399,57,-3576,-6059,-3203,-3046,-1901,1741,-3049,-964,1519,-2734,206,-2629,-3151,-916,-1187,-7768,-294,-3618,-4645,-192,1062,-2922,2224,-1887,-378,-1593,-550,10878,-4982,-2336,9335,1341,-4738,-2656,2252,-10205,-4692,639,-3422,-6953,1710,-2241,-2836,-1007,-3476,-3852,1840,-5581,1207,-4587,1271,2319,-1293,891,-659,619,134,-2456,-414,-3178,2626,3815,-1358,141,1527,4638,38,-1119,-4819,-5893,-505,970,-183,-375,1089,-1391,2731,651,-4558,-3356,344,-7651,-3920,-1793,-1319,-741,-5712,-1271,-2573,1728,748,-2374,-3447,-1850,-1185,-2225,1473,794,-2766,-572,5214,9750,-3200,1577,-2644,1801,3239,-6303,-4960,6596,943,-419,-6445,-536,1507,4780,11191,6845,350,2814,284,6796,3093,-19433,-4392,595,5834,381,5698,-13212,13671,-557,-7998,2885,3093,-3146,-1611,-9443,-3549,17939,-6899,1350,-8095,4233,4414,9345,1162,6875,7329,4096,3928,5917,-9,250,5263,14726,2609,3483,341,-2120,5986,-3996,-141,-1229,-38,-4541,6147,16660,4604,-4599,2365,8691,-2052,289,-7246,11757,12666,-45,-12382,-2408,-1839,-871,3269,8701,1857,2406,3615,-3095,46,-136,-234,3527,1268,-5849,-869,-1413,4621,-3708,-1771,4450,814,-7690,2729,128,-1519,68,549,5610,712,-888,4672,-1364,4003,-5024,-764,-2770,-6689,-8676,3999,-5649,-2108,4260,-406,-438,-572,-3916,2370,-5576,4328,6459,10361,-2492,325,-1772,919,6811,5888,-11601,-1068,-4072,-6845,2500,-2447,-2059,1943,2666,-1612,5048,-6748,3200,-1503,-4191,-4035,-95,-3559,-8178,-2800,-2480,1019,6372,4211,-956,-4750,9072,1040,2780,4257,152,-407,-2105,1802,418,-907,-2937,1561,1604,-1444,-1525,-6752,75,2663,5678,1202,-4880,6152,4179,9638,171,25,9013,2198,7309,-5864,-11630,-4978,-232,-1545,499,-6860,3911,-5312,2978,-642,-4587,8701,2386,5117,2496,1567,1378,4213,-3027,-691,-1159,-2585,-6967,2514,-5273,-1435,-1499,5317,3254,-5151,-8120,-1468,-7861,4829,-3393,-1986,4755,-2171,-1821,1257,1937,-2050,1821,9296,-4187,11640,119,-6201,3759,-185,-3232,-6806,-5751,-3762,-5078,2440,10703,3098,5346,3291,-3000,3229,-11044,-6513,664,-3381,2697,4655,-4016,2081,3051,2127,7177,1495,4145,-3735,-1983,-5253,-541,-4360,1052,7270,-51,-1233,-3337,-1578,1413,1365,-2553,-2067,-5014};
    Wx[70]='{-1296,8701,1584,-1429,974,786,1901,5195,1984,632,1364,1093,1166,-300,4636,6860,9340,5214,1804,-479,-809,1562,40,-3483,-1157,-372,2375,1258,-20,-1947,673,-3593,-3874,2469,-1033,-126,-1848,-721,-5927,-6186,3344,-795,-2449,-2043,-2260,-1674,-620,4948,-3427,826,3073,247,-345,-1857,2929,6948,-587,1230,-581,353,-329,472,-1448,2014,2890,842,-241,1917,-2048,1645,972,-4631,1866,-4487,1424,3212,-5410,275,-2500,1333,1512,-1853,-563,3190,-5454,3413,-1555,-2008,6801,-3862,422,-3840,1881,29,-6386,-1676,4067,-1734,3439,545,2343,11103,1137,481,-2191,1491,-4501,-4951,-59,141,10351,-3796,3803,11318,-13808,-222,3713,3757,-4360,430,-1733,607,-228,10869,-172,4980,4638,-9511,-13906,-3059,5571,-976,1560,14472,-2396,3525,-1138,-1002,2839,-7587,1054,24433,-8833,8696,1348,-3901,27,-3134,-2476,9018,-6611,2471,7006,1407,-2895,-770,1109,-1202,-5800,799,-2705,548,4780,-3515,2753,2048,-3918,1329,3864,-3559,3498,-17207,-7407,3093,-829,-6293,3618,-6601,-3337,-1459,1417,12939,-8085,2819,-2990,-8056,903,-3691,-7802,-75,-2104,-1706,-3640,461,4880,-2331,-3781,-9873,-145,2717,-445,-4316,3596,-3037,825,1748,-4301,3710,-3076,3452,-1015,1722,-7348,-744,4655,3266,1607,874,-1492,-1446,168,3767,-46,-1268,-7841,-4240,-8315,2486,-2032,-2220,-674,3510,9414,-95,-4602,-6049,-3051,-1346,5981,2851,-5537,-588,2546,6416,-4309,-850,-781,8984,396,4873,-1346,-5083,-263,-1232,813,-63,-6235,2546,-3786,2817,7373,-3562,-7597,2081,3474,-1606,97,-4013,-950,1605,-1914,370,-545,1254,1154,1275,-919,-2717,-2673,-3791,2165,-6191,-3845,-6264,-3105,6425,2871,1203,-11093,-2242,-5581,2592,3210,1462,315,4106,-6918,6718,273,-4931,2778,634,-198,2995,-2333,4013,3315,4172,2524,8740,-3322,2673,-1661,-6625,-1392,3969,3344,4172,-2276,-3815,-4655,3322,-230,-2548,-7358,-1439,-2131,5122,-1549,622,477,-5126,-532,-4147,-13398,-5000,-1881,-297,4467,366,-1206,-3876,4077,4626,3112,-4555,-2578,925,3591,738,10087,2570,208,-3010,-880,4980,-1136,-85,-8417,-2561,1141,-3364,-4851,8671,8935,-9809,-808,-6845,-10332,-1702,-4904,-3937,2502,3957,6254,-5424,-3522,-1737,-3249,-2675,5986,-1398,-2768,-4624,-10976,6264,5092,4365,476,-7192,-2805,-2797,5703,-309,-4094,11406,-3239,-874,-683,-3093};
    Wx[71]='{-2653,35,1745,1099,-666,-1396,1441,4685,-260,-4392,3310,3212,4643,-314,-4768,5107,546,-1110,1529,-518,1224,1694,23,-358,4699,-2504,1036,-1386,4895,-5532,-1875,4492,911,4887,-2590,-4716,2291,-845,-4477,3437,551,-4313,-3557,-2144,-5419,-3225,11953,-1956,4680,2687,4189,-2307,543,3173,-226,3691,2895,-1989,-1894,3850,415,304,510,-4313,5048,1545,-1723,7304,1749,874,4121,-1737,3422,-5444,2714,3710,4223,-5029,-201,2043,3305,5625,-3933,-2736,1542,6508,866,3161,1562,3200,977,-8642,-71,1165,186,1458,3000,-4265,4440,3076,213,-6250,-683,-8740,-6508,-2396,-2507,-3288,-4855,-5141,-12431,8730,10283,7675,8046,992,9624,2322,2949,30,205,9165,-5107,4765,1795,2276,-7529,-575,21250,2636,-5537,-353,-4045,-466,5117,1584,-571,3337,3164,10527,-3127,9794,-3298,3388,12392,-9482,-3857,-14248,5366,-11015,-15703,-13242,-9511,-5693,-4309,8891,-2626,1441,1140,4040,1549,6508,10849,2495,14697,-7729,7944,531,-2890,2120,9604,4445,-1196,2680,-2232,-6381,5595,-1801,-4462,-3825,-6557,-1365,4458,-11132,7495,922,2094,8457,-5800,5073,3054,33281,-7055,1205,-2111,-1649,2258,6933,913,6289,974,-821,2205,4206,-905,-1773,4392,2939,436,-3750,2071,351,-784,1317,-992,-5908,-9042,-4729,3112,-2467,-1059,1928,2995,2961,3146,-3547,4636,-74,-7583,8808,3159,-13085,-4753,-4775,-5463,2238,-1633,-874,-3032,-6313,4062,-9667,3266,-5029,-621,1773,-2951,357,5815,-4365,-6953,-11455,-1689,-481,5688,7954,-742,-1058,2293,-3991,4692,3273,5146,1608,16425,-1536,-4353,2778,-889,-2773,-2396,-9331,-3691,-1663,854,-1456,-11396,-2646,-2573,-4050,5512,-3842,-1267,-13398,4494,1158,2332,-1904,2668,-3032,3950,-4580,-3339,5449,5893,-7534,2375,-3859,3427,-6811,-6972,4194,5742,-9619,217,-3151,2739,1124,-315,-8969,6538,7299,733,-8046,-2980,-4431,-3251,-9370,822,-2875,-3994,-1889,4724,2812,-291,-4995,7397,-4526,4902,3630,-1057,-5039,1340,1030,-1942,1188,-2305,603,-7617,3212,1153,-6542,4057,-5234,14,4001,1223,-7036,346,-4533,-4504,-10908,1944,-1203,9301,7138,-634,2302,-960,-542,1984,3706,8876,2570,5390,-6269,-3986,1216,1475,-5639,-986,-418,-1322,603,7729,11074,-2147,-3771,2817,-8149,3420,-58,-10585,797,7338,-4709,7504,-876,1557,-10078,5649,-3537,5463,10947,-5854,-8139,-268,-1171,2824,-10585};
    Wx[72]='{24,-6411,-2768,-3674,-1595,1599,-6235,-4274,-2519,2233,1074,-3791,-1362,-1372,1982,-6982,-4389,-1723,-3200,446,-1306,1788,-1882,-3366,-2824,835,-1639,-2011,-4084,5117,-4023,-5122,-3730,-4389,1425,3586,178,-3625,-2242,-535,-3718,-6259,-2810,941,-1394,-4794,-1845,1450,-2169,-932,-1356,-7246,-1425,-878,1263,-12031,2119,-2641,3449,-3925,-3256,-2651,-2320,-745,-1723,14,1021,-5517,-2768,779,-3339,2099,-902,-766,-2127,-1950,-4306,1412,-15,695,1992,857,1063,1458,2077,2281,584,1895,-2763,-3796,2121,75,-2264,-1766,-3757,-5761,-2595,-9003,-4531,1121,-949,18046,-1894,-1350,4411,-167,-7221,665,5024,-3754,-4943,-4006,178,-1064,-25449,4709,-742,4211,-1024,-2037,-2443,-8022,-3427,-5825,1391,2423,174,7099,8002,-2687,-1524,-7939,-461,-14345,-2106,2238,-5468,-11748,-3364,-6254,11201,12529,6137,-2340,-5097,-4916,-922,7753,-682,1591,-4587,-13642,-2415,-11259,-1373,-7119,6376,5688,332,-6069,2768,11054,-6533,-6440,-16621,3210,691,-11435,1107,-433,278,3918,-3076,-9746,3759,1713,-15380,4760,2276,-1938,6914,17451,-338,-2722,3342,-15029,-2113,-10,973,-3315,-8500,-7436,11611,114,5649,-5756,4306,-4497,164,-6420,1340,4287,-407,-3173,2028,101,2203,-2644,10273,-653,6381,918,2856,-7729,3266,1364,2293,-5668,600,229,-673,-1342,4235,906,-1914,1058,-4291,-2961,4860,-6210,-270,-2773,5678,5263,-6826,-3049,344,3693,5156,3496,120,2365,-631,81,-2861,-1838,-165,-252,-1750,2863,401,-4135,167,-6870,-3139,13447,-1062,-1876,-9624,3239,-3476,-4201,10917,-447,-6064,1412,2199,-16201,1557,-1520,-5219,2609,-3840,-4313,-167,471,-151,-443,3391,-583,50,-3117,-197,6538,4350,2290,-1170,1212,477,-281,-2492,692,-7578,758,-7001,3369,-187,761,-2683,5190,10849,-4819,-66,-2709,6845,9077,-4694,3769,6899,2790,-4084,-4714,1654,-4365,-1751,3747,5805,-10205,5014,-4689,6738,-2420,2536,-232,-4672,-4218,-2976,5581,-4719,-5781,2200,-2376,2963,-650,4956,49,3996,1654,-1136,2692,-3466,-6044,-4838,-7641,-1749,-646,6865,3852,-1146,-427,36,2778,-6000,-3728,1805,6040,-2739,-4663,-4729,2036,-4758,-3977,-1092,4848,629,5722,1084,-5175,607,7128,2174,-4699,-1723,-5971,1929,-3281,-308,-6079,-946,5332,-1605,1845,27,1485,10185,5371,4606,-508,-324,-1350,-755,-7016,-6269,249,-10498,483,886,397,-4536,1008};
    Wx[73]='{1799,-900,-4531,2817,2966,1423,1738,-2990,1622,744,9580,-4528,4265,406,8417,871,6518,639,2644,1767,-973,-1791,-3374,157,-2687,-1954,-3754,1937,-879,1491,2114,10576,-877,-1779,2362,5957,4812,1700,4365,6250,5781,8911,4160,-1829,1762,3701,-645,4428,2415,-48,-1721,917,-1141,4079,-1994,-107,-1943,5239,-479,3356,40,-583,435,-289,864,55,949,4653,-4099,-3178,1357,3518,-2934,6010,2863,5053,2541,2902,2910,121,1427,4167,1191,4345,-1450,-3034,974,1113,-3427,-798,1842,3229,1470,-5004,-2252,-2030,-203,4853,-4509,3112,1716,-16904,1618,-10849,-153,-525,-9736,-1772,1375,-7495,10019,-1159,-5668,5849,1850,-10185,-4418,-2590,7016,-1760,-2932,-1496,-1520,1290,-3054,-2003,5458,-7290,6831,-11650,3247,-3339,-2687,7880,-1806,495,4331,1066,7133,-5024,-2272,3430,1408,-4482,-13505,6875,15703,-1910,-5195,-3415,11914,-8071,-219,-5195,6152,17441,-812,-2165,14238,200,-7275,-6445,-1054,-4321,9921,1202,1962,-639,2415,-2685,-2153,3515,3811,5927,289,-1160,-8359,2219,4726,-1771,-2268,11835,-1088,-22050,-5463,4274,501,5888,6621,3642,7758,9057,-1206,-1191,-786,3354,-6254,-734,286,-3400,1920,7353,-5380,3149,3090,-606,-1562,-9130,-4060,335,-6933,4270,5107,-4475,-2841,-10244,3967,1176,-2116,-645,-2187,-3059,-380,2150,-5371,1861,995,1607,-327,255,7661,-5244,-5029,-93,-3627,1618,914,-2727,-9770,-4587,-1343,-667,-9165,-4455,-8569,-4094,4853,-6743,3869,-1293,-6708,-1270,-6884,-4091,2780,-6396,-2185,1628,112,-2944,-1594,-2971,-3520,2558,-13710,-3774,-2939,-331,-2148,-5214,-471,-4260,-222,-7080,-770,-3688,1259,-530,5498,-4948,-3195,11396,-9199,601,-4140,-5234,-1246,-3630,2420,2624,1940,-1459,-1033,-6933,-2629,-3991,-4370,-336,-4501,-787,1201,4519,-6552,5546,2963,-2097,-726,-8105,-2929,160,-653,1661,3745,-4782,-1354,-4995,4604,310,-4782,526,2705,-130,1973,256,-3112,1597,-7216,-789,6923,-955,10585,1278,8076,2971,-7475,3933,-692,-3271,1893,7124,-2312,3122,2495,321,3388,-5185,-3193,1823,977,-1619,-670,-1568,216,2437,-10683,5698,-2313,5375,245,5952,9208,-2722,6425,273,-177,917,-10498,-241,-7011,-1696,-1109,12304,-214,107,-3840,1613,4978,-1551,2868,-8808,-7363,564,-1928,5410,-13085,-8564,373,-2440,6665,2687,-6059,3581,-3989,-2788,304,-3464,-8354,1101,-6972,2641};
    Wx[74]='{702,5625,-3049,759,1800,394,61,1231,-4592,-1390,-253,-2419,1702,7060,-1276,-4418,-3146,-1518,1401,-1701,-1296,2038,2326,1481,-2287,798,-2849,-1292,540,-1978,2326,-5336,-883,4226,-5219,-3017,3950,-522,-5156,-5097,1557,-9995,6381,-1119,-3540,-2454,-4160,-6132,-2297,1774,-4682,4577,-3652,-3957,-1473,-3415,-1145,-1682,-2966,-5234,-1223,-4174,-474,-2646,-2595,235,-3271,-8159,2019,1822,-718,-12363,3911,-3454,1335,4941,-8417,-4379,3437,-3723,2739,-8730,-337,-3515,-874,931,-4228,12,3112,1420,-789,-6728,-3935,-3698,1328,1226,1392,-4785,899,620,-1475,812,-2276,-16669,1704,-1274,4870,3632,7084,6088,-13505,-1535,4199,-4807,14658,5346,2066,-9379,-96,2871,1619,4699,-13505,-545,3017,2558,-8110,2783,10097,1477,-10712,-4992,8593,7846,-2802,1170,-1988,-2381,-10517,3339,751,-7089,5112,218,-10566,-9287,6904,294,4665,364,11748,-5869,-6079,3388,-2819,2489,-6713,-1639,-5966,429,-1356,-1154,4929,6791,-8876,-70,-874,9125,2369,-814,1630,5268,-2127,5361,1313,-6855,-7119,1624,22187,-3549,4853,-2219,-9394,-9877,2462,6884,-1229,3828,-753,5996,-1335,8779,-9018,1950,2197,-13300,5922,102,-1845,2512,-4174,-2951,1875,343,-5195,969,-6679,-2548,1024,-1252,5146,-7285,-440,-2069,-3037,-1506,-4787,-2347,944,-2404,-1893,254,445,2641,-852,569,-1694,2010,-4729,1,2685,7158,-5952,945,4887,7070,378,-2415,-8876,2556,1416,-8076,-6308,-9155,-7324,-821,-5488,318,-475,539,2309,3608,-6899,-3100,-527,-3393,2012,2325,-2181,-1499,2011,2897,4204,8574,2203,6459,-2138,7626,2279,1229,-6611,2658,-297,4050,-1489,-3847,-4660,-38,-5292,-2963,-835,-3559,-4675,4355,825,-8862,-4375,-5336,-1564,4050,7373,-5253,5761,2624,9882,4123,1563,-9194,-332,-1131,-8833,-1221,2524,163,-443,2656,-3925,-5390,-6093,-186,-491,-903,-3918,-2034,-6254,-4916,-5576,-10917,2543,1639,2512,-1690,2761,-5507,-6108,6303,-3676,-2902,-9433,-2406,-1345,1618,3518,-772,4719,-1691,6323,-2333,-2590,-2236,-3576,-12138,-1195,-4274,-7133,-2122,-1488,-3012,1752,2175,4953,955,-1911,-1435,693,3913,3403,5390,-658,6230,1221,-2274,-8286,8237,4577,-919,-5625,270,-17988,-3293,-6020,-3864,-6577,-1756,4509,-136,-2175,2343,2719,-4587,-3315,-1233,-4384,-1939,-8735,-6118,-9252,-3715,-2683,893,3332,-10634,1064,1184,714,-3312,991,-9140,-1265,-2583};
    Wx[75]='{1287,1462,-1331,-3156,856,437,4851,-1466,2785,-1788,-6977,-2235,-3457,8579,3178,-2071,-4243,3708,2366,-1923,-983,-838,-3100,377,-2883,-1611,-2973,-2277,3752,2341,108,9199,-9345,-316,-3864,2624,-5166,-389,-2753,-225,-2570,-2165,-1756,1105,-3259,-4409,-5664,-380,-813,2463,2119,6137,-2081,-3376,-2731,-5566,-2741,-6005,-2880,-4458,5112,-2985,789,-1655,-5546,-239,-3952,-2883,-102,-1651,-496,-4682,4980,3911,-5825,-4404,3364,-458,-1643,-2910,2248,2641,-4477,-287,1550,-696,-418,606,-731,-2028,480,-5849,-2059,-1798,-10605,173,-1915,-5996,634,201,-2807,-11953,-1838,1357,1185,805,1008,-9433,5664,4685,2386,-2047,-3271,3166,-4179,-7680,-14853,-6948,-4587,-5410,-969,-214,5322,5249,-2626,-606,-3896,7509,4680,-4291,3422,6840,2059,3242,-2946,7846,-3928,-4455,-1098,-949,-4042,617,8432,3303,-5698,5375,8730,-257,-4101,2230,-5947,23125,-5107,10732,418,941,-5195,-3662,20,-1651,-8666,4077,-6303,-520,7719,2705,5317,-510,75,-3513,1218,-5917,-901,4770,-2666,1092,-3571,2457,-4265,-144,6416,-5478,-826,9833,3652,1685,1531,-3730,-1264,-2304,-4052,5937,4353,2297,4936,3601,12714,-6547,-1574,-3149,-93,-10898,2731,-1236,-2379,902,-3808,-489,-3117,-3188,262,5190,1103,-119,-411,2985,8432,-3107,-874,3161,1210,3103,-3750,1771,1914,-2595,-489,-4143,9189,-2500,3740,10751,1788,3278,3017,-47,2121,2939,6611,-380,3225,-8818,8784,-3522,4558,5581,3669,-6196,-2954,4340,-2641,-8237,-2663,-690,4172,1156,-5971,-881,-4663,1557,-196,-127,-1895,949,6586,2316,2519,9472,-2075,-965,3967,1098,-788,-4982,-4755,643,-469,4816,5634,-2249,2413,-809,-1752,-1223,571,2512,-2412,1510,-7221,-1215,-673,4267,-6948,-2326,-6308,422,373,3315,-3352,3142,-4619,-9794,3146,2731,-3181,-13720,-380,-8515,-2832,-2617,1275,744,-6484,-5620,-4523,-62,4519,3937,650,-6811,-15039,-600,-2563,1198,-1303,2565,-346,-10097,-2597,515,-91,47,-5517,-5747,1724,2573,2844,-9326,173,6430,-2963,-4948,-1547,5478,9018,3786,-6723,2875,-4904,5947,5444,800,-83,-3056,4846,-2019,-9238,-1473,-3662,-4919,4653,-1216,1428,-999,2490,3867,-6450,1282,1448,-11250,4841,-3256,-214,8339,-3962,-5781,-3984,2646,4013,-6464,2452,-2648,2257,-4599,2375,6962,-4035,3903,-2086,-6572,4572,-1483,290,-822,-3815,1275,2626,-3640,-5317,-607};
    Wx[76]='{944,3081,-39,-1276,-4479,-3771,3623,-498,1793,-2543,-225,1026,844,-3015,1488,856,723,6479,3107,-2193,-3750,-4174,3627,-83,2008,1608,58,-226,-7207,-2159,2165,1499,-3825,5268,-5668,-4895,2292,1337,20,-1189,-1070,-1339,-764,2827,2670,1842,-273,2592,1140,-213,-1755,2373,-9,1373,-430,4565,-1284,-819,-1162,1634,1435,-1811,-527,2413,4069,-947,83,3754,-2474,1188,-1284,-448,-4831,-2386,-1104,2286,264,412,-116,-2509,-3300,14677,-1636,6865,895,4077,-5629,-1604,-375,-4626,1060,6430,173,-5166,2585,-2863,-1140,1984,3439,5346,5922,-213,1313,-2110,354,2205,-4699,-7646,-1645,-134,9956,-4746,1682,12402,-14990,-7045,5117,7373,-1599,-387,-3444,-6088,-1915,6152,3732,1835,-3503,-5371,-11093,-5957,-6547,2763,1084,6313,-4692,3889,1069,4089,15468,-16435,-7758,-16240,-9262,-7016,2373,-681,-481,-13789,-5131,289,17265,15117,265,-14208,6044,7739,3901,1335,1412,-1948,-7036,-2242,-1508,6298,4306,4077,-952,-8730,-3684,-433,11044,-10654,-2303,6552,1195,5268,9604,-11630,12070,-5585,-2651,-10390,6586,6577,-426,-5961,9243,11992,-2396,-428,2741,1346,-6518,5039,-8007,3291,4294,-4909,4011,-4838,2198,4370,823,-5009,-102,-128,-780,731,-1271,-1660,-5927,-5141,-774,-4094,8608,997,302,-294,3835,-5473,2770,4333,-2135,2116,-4675,1884,3603,-612,-7207,-1000,-1024,-1220,2812,-7509,2209,-2507,-133,538,-3466,-4660,2390,4592,4306,-5004,-1275,-2456,2249,861,4348,-1156,-720,-5673,2023,442,-371,11259,422,2220,130,-631,4311,3657,-1960,-3881,1926,-6372,-1506,3398,-175,4145,-955,-5024,-186,-3823,-1440,4545,2452,-8242,9125,-2895,333,-4213,-5375,-6562,2204,-3925,24,-3564,1292,-2504,3532,-1139,-141,2666,-7558,-2502,-7446,-6572,3347,-3078,-4089,4689,-1859,579,-2185,-3425,5366,9033,-1540,3146,-7167,-4790,-4675,-357,-488,-3093,-3024,5170,1029,-3642,174,1783,1218,2644,484,4062,4538,-3330,-9272,109,920,1211,-3520,2644,-5224,-2541,-4560,6738,4064,-6938,374,1227,5092,-1328,5732,-82,-7148,-7114,4738,3127,-3598,-7700,5063,4467,10693,-3061,1120,161,2196,-1430,7392,-1639,2453,80,4609,-455,-8554,4621,9799,1550,-859,1232,3022,-4384,-825,7709,-1480,-4775,1195,-4055,-718,-4926,-7998,-908,11435,932,-9643,-2269,-654,477,1414,-7407,3061,2727,-1445,-1611,3574,1945,4758,-756};
    Wx[77]='{-2631,-3928,-2156,-1724,-406,-1066,-1110,-2427,3356,-3173,9072,-225,2479,-4316,-6074,3867,3969,1252,-4560,893,3632,-623,-2912,-479,-2416,-3176,-1271,-1341,3764,1818,2712,-1188,-5346,1734,-3493,-801,2507,-5253,296,-2418,-4101,-5292,1128,-7944,2476,2268,1921,-1444,466,-1617,2770,1762,3032,1007,3164,-2832,-371,3132,-2181,-594,-3244,-7934,743,1464,2976,2326,-3725,4855,-4174,-1403,5146,-3120,-1071,-3405,4479,-3444,1958,-1298,-147,-1828,112,5439,-3549,4609,-1319,1905,-664,2687,-546,5219,-16,-9370,-8662,4333,-3708,-1959,1784,-470,-5043,-5229,1014,2497,936,-6694,-8881,1776,123,-6879,-2121,-2602,17294,-1978,-7724,-8652,7509,-4311,-6611,-318,4682,4946,-291,1273,-550,2495,-4248,-8945,-2401,-2770,7480,-3967,8676,2124,-10634,20273,2086,-1617,-6098,-4289,5371,14804,4863,-1931,-5883,4650,-8681,-9609,-3310,3317,5981,-5908,-19423,-8378,-7993,419,-2929,9926,13183,-927,-534,-5537,-2639,-11806,-822,-4587,4924,-487,-1768,8359,-2099,538,5297,5493,-1143,-9858,3942,-19902,-3879,4624,-1535,3354,-6235,1999,-1613,-10302,111,8608,-6826,6171,-492,1785,9487,24199,2912,-471,-5854,4438,-6362,-16162,-8808,-6367,5395,-988,-2258,264,5048,-657,-955,5053,1391,3793,3796,-341,2749,6274,2440,4309,1331,1380,-2890,7084,-3056,-180,2561,-1491,339,1116,7832,682,11914,3911,-531,-6333,4511,8481,-1884,-153,-3830,-145,-1507,-4543,1949,1123,5747,1155,9184,819,14882,9985,4584,-1336,-4040,2712,-3718,-13632,2802,-1,2053,-1149,3891,-6430,217,2551,-3044,-8403,-3222,677,-376,7026,-322,-309,-7812,2644,419,-435,3559,2136,-2125,2498,-2023,123,1021,-6044,-4089,6367,7241,-3037,4116,2369,184,108,-4304,174,817,3015,13623,1439,-349,19199,-3991,1217,1335,1420,-14980,-3806,2917,-2661,-1015,6982,-7309,-155,7216,-1711,4787,-2773,5937,-3808,1658,-4150,-1386,-6787,5913,3195,-1296,-1064,812,596,1018,-2863,8081,2196,-3027,-5092,2432,-3085,-3154,-1065,-2130,-56,4665,-2529,-6469,-4873,2172,5932,2225,520,1761,31,7094,-1645,-4909,-4550,-16103,-5351,4887,5932,2985,-8193,-7504,-8935,-3286,-1975,2384,-3337,-2692,490,-7910,2824,-10078,-5009,-1947,-2729,-1531,3356,4890,3576,2575,-4047,-403,-3791,-1451,-3022,-4719,7480,6669,-6240,1700,345,-1628,-8369,-514,2282,-3630,-3024,9965,246,-4914,2148,-2412,-4775};
    Wx[78]='{-2902,-3862,-4235,4418,-960,1879,-1754,-624,-2568,893,-3310,-1163,-2014,2470,-295,-1402,-6352,-752,-5791,-760,-2000,-552,-4287,-239,-4863,-3798,1392,-1132,-1882,-2770,-1090,-4611,6337,-561,56,-1932,-4738,1553,-3447,3056,-4018,-5029,-3364,-3847,-10029,-40,2484,574,4399,2885,3596,-2858,1523,-2761,-4978,-4375,-3723,-762,-1497,-1341,-7827,810,-1009,-5234,-3063,6137,-1892,-3859,447,191,-4128,-617,-3933,-953,645,-9301,1125,-213,4746,334,1335,7329,2144,3122,6044,-4421,-287,3554,96,917,-1076,3901,-7470,6533,-3725,-1398,-3708,-3608,-1492,-3344,-4533,-8496,-504,2683,-3789,-2324,-4030,14082,2932,-1060,-9111,-313,8129,-10224,-2071,-6059,7539,1397,5034,572,-908,-2468,4602,-10273,-10605,-6958,4038,-993,-32,127,-1768,-9980,5107,15839,389,-3608,-5595,-3122,5839,2905,2900,-4050,3354,-4611,-14472,12216,3205,4804,-2427,-2440,2399,-4140,-2309,4079,-1201,6040,-7768,-2211,-9223,-1320,-432,6860,457,1130,9252,-2978,-1187,-3937,2075,-2631,-4245,11982,4536,-1279,3364,972,-6743,10234,10947,9165,-127,7968,-4199,-5234,3430,2641,-4584,12568,7563,2100,-4475,8085,5136,817,-15664,877,524,-20332,-6206,-4055,1297,5454,-2391,1044,7080,-95,759,-7485,505,2319,4216,-4584,-8261,2985,1269,-874,3291,5498,-7871,-92,-689,-184,-4077,-914,-2174,-942,1335,75,5815,2152,6508,-5249,2083,8554,4396,-1676,12001,7211,-4060,-3803,10322,665,13750,1634,-1951,5019,-22226,-2392,-2248,6586,-4282,3083,-1778,-2478,2006,13925,-3515,5908,6176,-1816,2890,3459,6503,-2238,8789,3632,-226,-12509,1955,-932,-1918,2346,-1975,-9638,1343,-2246,6669,-618,1436,5195,941,-1827,281,-3840,3378,7827,-930,1591,-32,2309,4702,-2761,276,6430,841,252,952,10400,-3447,10048,6826,5751,4162,2722,8823,1221,-1287,-6899,-4196,-6909,906,-3725,-2631,6005,-502,-5844,1688,-3156,-2836,2917,3081,3029,-645,1922,-2384,-2082,3264,2308,7910,-2512,5874,-4729,1058,5122,-2504,3881,1669,5380,335,3442,235,-771,3569,8774,-2783,2213,-9350,-1513,14873,-4074,-5166,-823,1711,2319,2034,7939,-3483,3764,-492,-3605,-3349,-2199,3310,-1796,-371,3461,-912,761,-7241,-10302,-2410,-5024,-5361,-6303,582,-2517,7021,2187,-199,881,-2873,-3806,-1384,-1641,5058,7822,-696,-3085,-2670,4465,-3366,839,-2369,6801,5683,56,4604,1113,-12001,5307};
    Wx[79]='{1622,-254,-1959,1168,3474,-953,-7631,-462,16,-142,5390,2410,4411,-3315,2592,4172,-2131,4338,3051,-1019,791,2324,376,-2421,2766,1188,1187,-572,2639,-1076,-962,4089,-4228,339,3232,1611,5805,-5151,1141,1087,1833,2321,2626,3735,3488,-757,-1818,3649,4721,1993,1644,-6030,-285,1328,-1721,8901,-1239,-4592,6855,8457,3959,-1630,4758,3959,3564,2447,4504,-4885,4152,3425,5527,7480,1695,-4125,-117,877,2496,-2144,-884,1734,-2244,-1501,-1680,2998,2983,-1470,2668,-2934,6391,819,-2467,-6474,-2041,3576,2534,5361,442,-3791,-2143,3125,-1015,6284,2357,-973,11542,2341,2349,6132,760,3205,-16103,-3066,-5141,-17314,8369,-6708,-17119,-8666,2712,361,-1055,123,-2675,808,419,5766,-6020,-4179,5610,-3430,-11484,-13369,1242,-4257,1433,9326,3291,-3188,-9931,1911,-2413,1654,-5517,4636,-570,1312,-1612,-485,9692,-1778,-3271,5312,2006,9125,-1959,-4956,-750,3706,-4118,-209,-62,-16484,-2397,300,-10488,-1524,-3820,-10585,1020,745,679,-3281,-1262,517,162,4326,-2478,-3669,4868,-1618,-217,836,-2308,17373,-7358,-8471,-1204,-7724,-8886,-1085,-4118,9018,2163,-2880,12431,2507,3532,-6181,-274,6157,-2622,15205,-1568,-2595,262,-1807,3105,2006,2934,-75,-1391,-1754,-112,-270,8310,-457,-2595,-8735,136,826,328,7724,2629,2724,289,-4409,-2081,153,909,-1052,1650,-9194,-3447,-1254,1898,1354,-2985,-2966,-1306,2954,-1271,2949,5224,2248,6440,2398,-404,-3393,983,2150,-1137,-16220,-877,-440,-3330,-4191,2171,-895,-2624,-6435,3100,-677,-2954,-8134,4426,-2314,3415,3117,-2087,-118,922,-704,-608,-3947,861,3488,-7973,-81,1019,-5507,-1357,-13671,-2583,-4296,3503,11865,865,1072,1430,-3591,983,-3676,3532,-4072,-14042,3205,3928,-5087,3625,-6416,149,4426,-10429,-1937,3513,5292,-2197,-1361,3923,1225,-1450,3186,-5249,-9501,-4184,-2683,383,-5424,4816,-999,2617,4157,-1188,-4130,-2670,-3100,2680,1671,-3417,-4667,-4792,-3249,-1121,-708,-4218,2091,5288,580,127,4992,964,-9335,10644,-7377,1528,7509,7114,5766,4951,-3295,-4655,-8051,-4230,3408,6083,4301,5590,1973,1078,5756,5268,2841,-12187,1525,2495,3129,10429,-12792,-5556,2580,2512,-2658,624,1185,7255,-92,4226,-2292,-7871,-1622,-1833,-9091,-3259,-9687,-5327,-299,3273,4157,3920,-2751,5214,-5454,2379,4155,-4760,3576,1351,6176,5893,-6391};
    Wx[80]='{725,4389,-338,-2003,-1462,-491,-631,2861,-423,-1601,-2094,-956,2482,4260,-7973,7436,-1065,-1569,-4497,232,1081,809,-714,-2651,18,434,728,1789,-2287,3447,1683,8813,4812,-1901,-2368,-3186,1405,99,4360,3159,715,1157,-5200,2342,-2457,6865,-3469,3176,1209,-1569,-1690,347,3662,2924,2709,8505,-467,-372,717,3017,453,2871,1219,1260,-7714,864,-1818,1182,1450,1499,121,5205,1099,-3967,597,1174,714,-154,114,-2729,-4118,-2971,-841,4816,2177,1892,2578,-759,2885,1577,-6264,-4372,5639,4902,4162,1881,3603,1005,-3063,7514,1693,-583,5751,632,-4213,1190,391,-1809,-597,11123,-998,-6572,169,-7954,808,-6074,-3757,1328,1745,-852,1408,4936,-1350,-2338,-872,-8500,935,-984,-9184,-2406,3068,-8930,-3386,1258,-3503,-8583,-6821,5742,-2634,8676,-4357,-2827,-21386,-9521,-1336,-3293,-15234,-2773,2221,-492,969,-4379,491,426,-1976,502,1849,-2185,8779,-4384,2426,-10019,7050,-7729,14560,-4479,4077,-1573,-2644,1529,18896,-5937,4187,-28,-4606,-7133,-7636,5512,9453,-4123,-8305,-5854,-221,17646,2391,-2785,-2995,340,-5039,-639,5849,-5117,1588,1748,3000,7758,-5708,4819,-7387,-22050,-4333,-13730,-2639,-4294,-3818,-1231,6435,6513,7875,-3208,-8603,4316,2377,339,9609,5527,9160,1779,-4187,791,2758,427,-2922,-1800,-8027,-539,2430,567,187,-1752,294,-1231,-1807,-1964,3046,-3491,5043,-986,1395,2292,-4274,8437,3161,4287,-5312,-2066,20644,7236,-1357,-11142,-4431,-5625,2286,-3549,3808,-12070,-2966,-114,7578,993,-2397,-583,498,630,3300,-600,-2871,-3991,4284,1279,1855,8510,3210,-148,190,11630,-4611,579,-8149,471,5375,4431,-3884,266,1405,-76,345,3425,4042,-1152,31,1533,4094,5170,1357,2119,-1983,2565,313,-1174,-1496,-5151,955,3933,-6225,1657,7050,8940,2846,-2961,-2678,2829,-2924,-1461,2802,523,8867,-1961,-10683,-1894,3479,2301,-1011,-7333,-2861,-1228,-166,-1923,-2484,5224,-315,-654,7177,2663,-6787,-3918,-6547,410,-2440,-2292,456,828,-2426,2496,3295,-648,-3400,2954,2697,-760,1375,-4567,4338,4604,-2565,-14902,1586,-3989,3671,-1295,-2556,1855,5131,-7524,-4899,-1077,-6372,-6235,-2797,3481,727,774,-4497,-5146,-7382,-1700,-5312,3122,5449,-3249,187,614,-11103,1260,-938,-1610,-6992,6035,3857,-1021,-3588,2651,4487,5820,2071,5922,4592,1419,-3054,2325};
    Wx[81]='{819,-668,-3854,-614,213,1276,-2675,3793,-2186,-1649,-877,-2512,-498,-349,3325,3776,2824,-561,2539,2067,2225,-354,-569,-1164,594,2160,2590,774,1364,428,-507,-1658,-1671,-2814,3439,811,1607,173,3688,-3039,-296,-3500,-858,-8593,4667,-2521,3747,-518,-872,963,-3747,-4138,-1589,4995,-2487,-432,-1372,-1333,-3681,4099,-2822,-5375,3505,1715,-4514,2976,217,-3884,-1187,305,-2604,5083,-1940,2800,-2851,-2292,-900,-757,-2182,-795,-4543,-3259,-2150,459,-3989,-2435,106,-5166,-168,392,-673,-1242,2636,134,-5932,4167,1868,2114,2924,-3813,743,-3503,868,2822,2257,128,-6093,-6665,-1243,-53,-9833,2763,-4372,-4467,7270,561,-9335,2895,646,-5712,1591,-6333,7148,-2817,2958,6909,2534,-1887,-2641,-5195,2563,17949,8437,5791,3361,4082,2529,1594,3559,-9809,1562,5024,-8891,6840,-4682,7539,276,1367,2327,-4345,8334,-16767,-1022,-7192,2712,-2907,-6513,-4006,3757,-1805,-3215,1748,2578,1010,-1405,894,-2934,-14345,3784,-6015,-4470,7622,678,6049,-163,-3801,-6782,4035,3183,6352,3583,2075,-6093,-4802,-874,5312,439,-2403,4914,4631,-3864,4916,6562,-5351,6689,4602,-158,-11689,4580,5483,-989,-8437,-1039,98,-2954,2043,2486,-4445,-1716,787,-4692,1520,3884,-3339,-2386,3190,-7836,-5546,838,927,308,2629,-5043,1242,2073,-3017,2415,1452,-2478,-3430,6264,-5034,5771,-393,-6308,1705,63,2866,-4914,-449,5942,114,4621,7543,-3947,-2753,-11699,6176,-677,2242,-1961,802,-3684,-2496,2484,-4177,-4716,77,-6333,-2438,-1861,-12119,-6538,-2008,2868,-97,1289,283,-578,-2341,2214,-4443,-4343,-4143,-1182,-1028,10068,3806,-97,1069,-4265,-4577,3613,1466,2056,1821,-2988,-854,-4570,-309,-1254,3552,-904,-8662,7094,-6831,830,503,-536,-4545,2174,-4401,1198,2602,-974,3051,7602,-4309,-9418,3063,-7319,-569,160,3994,-1436,-4287,-5019,-3964,1658,-6333,3249,921,-2457,-702,-1016,-2529,1147,803,-5332,-4897,-2871,-9809,2156,-3447,-5151,-1110,-1684,808,4899,1899,-5595,-5112,2424,3974,192,-7412,-10029,5317,8159,-975,602,383,-1386,-4074,7866,-1864,-6489,517,-4284,747,1201,-5532,-1842,-721,-28,4880,-573,-1112,-4511,-2541,-3254,-6899,-1291,-3503,1124,-659,3872,1134,996,-6738,-6113,-1006,2009,5102,413,-3837,-2272,-2194,-132,7026,-2078,2692,-8344,-8745,-5405,2819,4729,1712,1768,-10683};
    Wx[82]='{2091,337,3483,2183,-3671,52,2448,2524,1359,-2469,-7475,5566,1947,5888,5952,1440,4257,-5864,1078,-1600,-328,868,3723,-338,-384,941,-2307,207,1534,-1705,-246,-8657,6044,1732,7944,4594,1986,2119,4248,-579,4465,-263,3967,-3237,4790,-8359,7626,2429,-1870,621,-266,-2301,5576,-465,3847,3195,-1972,-1308,2976,7163,3759,4677,3100,-3078,-5053,-3364,2905,-6416,1561,2807,1065,753,2301,1939,1721,7446,717,-1356,459,-1361,-120,2978,2106,7612,-1990,-2071,-3889,858,3911,655,-5942,80,5766,-1872,-2309,-525,1308,-407,4274,-538,1502,10937,-1864,-6093,-1645,607,12158,-877,2165,2780,-3659,3249,3852,5112,-4060,-817,9667,-8540,-2988,-3627,1110,3613,-6796,7602,5629,6000,570,787,2001,5083,-4846,18085,-693,-1457,3974,-6948,1937,2604,-214,9399,-9428,-6240,7504,2355,6757,8041,-13242,4167,-5263,-2495,-9497,-9418,4963,-493,-6376,1906,-1447,4418,14775,6328,1251,4606,14267,3574,1241,3713,-3178,13125,-905,4028,1607,14990,-2226,3767,-3913,7998,8916,4619,-9423,-11650,1064,-7612,8217,-701,1275,-712,4541,1973,3232,5375,9052,-2839,-2770,514,21269,2683,-3100,-2237,8930,5122,-2036,5800,1689,-967,-6547,-1855,327,2337,-1536,-3789,7368,433,-4804,5024,-2744,-6201,-2196,-1416,5092,585,2583,-89,-1348,-4479,550,-1193,-3989,-1602,-1539,-4057,-1329,422,-6503,-863,-11240,4645,-7280,-2005,-1279,348,-6474,-2169,-1083,-2200,-11357,1306,2019,-2218,-2257,-6401,629,8208,1861,-946,6411,-6020,4533,-2218,-1772,-43,-1405,-3637,-5498,7592,-2390,3679,-2719,-5942,-1932,403,3693,-2985,-2260,9580,520,626,-8427,2912,-4006,-3032,-655,-5166,725,-2432,-2204,3784,3642,1762,-2604,-1309,-3129,-1157,-2807,-4162,9892,6210,-7216,-635,-3325,-2929,-888,7163,9414,-2041,-3664,5986,-522,1590,1678,-3837,3251,6074,3728,-1811,529,763,1864,4165,-955,90,1394,-671,5000,1203,-8911,2565,-850,97,1197,7583,4682,5292,-1575,-941,3137,2211,3198,-2150,-7104,-2149,-3420,-4731,5053,-8212,-1993,1730,4821,3066,-7324,2521,2702,4438,7895,8457,1910,3281,4916,-8232,4516,6708,-9023,1790,5209,-952,2844,-7802,-1243,-1411,-3735,5722,3474,-3916,-8198,10546,-4560,3688,4680,10273,2182,-2756,-656,1950,4328,60,-14609,5771,-3959,4157,2687,-6401,1051,2276,1774,-25976,-7011,3432,-8798,-14257,534,-1916};
    Wx[83]='{-582,-1033,-401,-1933,2026,-577,-912,-972,223,-3911,-905,-5029,2587,-1739,1628,6660,3608,-1771,-1656,347,621,-2966,-1280,-131,2465,-3894,-2232,-1411,-1236,2583,1002,1259,-809,-999,-3876,1892,-3303,-1593,-786,-3964,-1370,-55,574,-5595,-1088,-2471,-4663,-6445,364,-948,-8164,-2512,-1979,4440,2719,-1582,3085,-5478,5122,-6108,861,-3525,-4113,2934,-301,913,-941,-5898,1672,-219,-2973,-1334,5781,-301,-1090,-1550,-4826,-3613,6899,-3422,-1053,-120,-759,6000,642,509,-234,-785,832,-698,1522,-701,-4401,4128,-5546,1606,2263,3854,1580,2517,5053,-2651,827,933,-1412,-1651,5327,-1815,-12812,-209,10634,-981,5473,-9262,-15214,-4467,-14873,-4526,-5034,-4250,-2863,-7963,-6035,-6967,2449,-11777,-2397,3886,3627,-6840,4108,629,-5942,4670,-4916,-3479,219,-533,-15253,6494,5761,12558,-5434,-18310,-14716,2274,-13798,-4846,1132,896,-6816,1259,-3129,-5058,9023,-949,8354,1516,-4382,-6503,887,11992,4243,-9760,-1523,277,-3364,1087,-1124,4985,7763,4606,803,-9042,451,-3732,-6464,15927,4838,5493,3425,-13662,-2303,5966,-3078,-1063,-505,744,173,-233,5766,9970,1649,847,2607,4904,2087,-6826,731,-15039,-2448,-441,-725,-284,-4636,710,2829,-3583,314,-3549,191,-1904,-5395,-5463,-8725,3425,3132,-1496,1596,844,-1851,-3317,-3176,-2185,-2556,-1783,-2519,-5454,5385,-2181,43,1724,9497,-442,-3723,-3054,1413,3166,-3024,9497,-3256,12617,-2482,969,-7558,1682,219,11923,-727,1809,2475,-2259,-2301,497,-2437,4992,5454,-6040,-4313,1252,1994,277,-3151,8168,-3452,330,3698,11953,2147,-554,1959,4086,2176,3742,-890,2812,6928,4465,5292,-794,2873,9755,-4296,8769,997,-1842,-1508,54,545,2517,-7890,780,262,4880,-1484,7666,-791,896,-6625,-8730,1109,-6660,-19511,3811,-3337,-1440,-1100,1915,-6298,-3317,-3957,-3586,7978,-3596,-5932,-4638,-3972,-5522,-3784,-5712,-825,955,-9287,-3222,4270,-572,-1655,-2022,8872,-969,-3254,1726,8417,-2092,9819,334,-4118,4965,-778,10585,-3710,1079,-679,-5620,1148,-3586,7309,3889,409,-336,-2836,1608,44,509,-8354,-1884,8110,-10302,-1156,-3596,-953,-1264,329,-1979,-2624,-8193,8349,7080,-1848,186,6542,-1215,-1683,6660,-6894,1354,3967,44,9365,2392,3210,-5488,-5781,2614,-603,-181,-1414,-448,3928,1954,-5346,733,-5400,2797,1901,2137,3906,-9921,3073,-6938};
    Wx[84]='{2491,1916,-1733,-1373,622,-1369,1494,-1162,1933,-1331,2215,653,33,4189,5297,84,2670,732,-223,969,-1589,-3686,-3789,-1995,3383,-5151,2027,-765,1516,21,-562,-486,3974,2368,802,547,-409,-74,1319,-5957,-662,2810,1601,-3457,265,1568,10830,3442,-1833,-280,-3757,3745,1379,-319,2597,-3798,-153,3815,1405,-6098,-1754,164,2271,-1965,2458,-1821,-2396,-3100,1580,1094,-149,3388,-2348,-1689,-2680,-1674,3112,-125,5688,252,1231,6201,1297,-598,4865,2276,-2354,5659,-4008,-1041,2731,-2578,5854,-3586,-5092,3381,2934,761,1115,4841,3657,9013,1309,-3874,-3613,-269,5122,-6962,-1163,5195,2280,-3164,2768,5341,423,-19980,5590,-5937,-4868,500,-465,-3452,-1844,3811,4768,22,-3745,3364,-5141,-6655,4433,-1300,3754,-2817,-6674,6938,2402,-1134,-4523,-6171,-5297,5615,-1408,-2114,-8417,1429,4104,4826,566,3828,9648,-358,1226,14736,4941,8940,8061,1414,-1296,-3110,-852,-11171,-8046,-6381,-7172,3627,-570,21660,-4106,120,9697,-6840,-98,-7749,-1441,4916,1369,1229,422,-8378,918,-8417,2022,9169,6733,-443,2548,8657,-5888,3034,-1658,3493,-2587,4213,-6464,3647,10136,1182,2707,-17998,-1466,-11074,-2229,806,-6313,894,-4931,-1051,-4672,-4812,612,-21,-5703,-11904,-209,-1313,-7548,-1663,3002,1588,1138,-897,908,-9907,-2924,244,1939,-1052,235,-1235,-6352,-8354,-5639,-6645,-4028,-1066,-4572,-1049,-1582,3872,-5502,7832,4213,-2741,-2082,375,-10361,2919,-1062,-1773,8989,-1320,-907,-894,-2093,7500,320,881,1707,8588,339,-3828,-6406,-2983,-3381,2614,274,12597,-911,3366,-6718,458,2614,-3208,-6523,-1057,5590,-5322,1682,-1922,-3266,-7353,-7119,-3686,-104,-6962,-578,-1429,4782,2768,-874,-2634,-3713,-738,477,-330,1296,-5102,-2834,-9736,-419,-6318,-5375,-1555,-6445,-1383,-3698,31,-1452,-3439,-2028,5654,-1156,-1674,3471,1943,1835,2070,-247,-1728,-1389,-3527,-6269,-1844,-2360,12158,-769,-2639,9809,-6767,92,-1630,-732,-1389,2060,21,-1495,-802,-1776,-2442,355,8364,2215,-1640,-11,1992,-4187,-869,-8417,5825,8339,-2335,-6333,1566,949,51,6777,-4392,-1998,-8037,-881,1168,-9428,-6826,-1990,2104,-5483,1629,6948,-2846,-417,1700,4394,-2456,-4667,-1644,121,-5092,6904,814,-2047,-7045,-4865,-5229,3823,-1549,-2944,3403,5776,-2849,8735,-6259,228,1278,5517,-6079,10751,-7275,-6020,-3190};
    Wx[85]='{1004,131,2238,-1044,1313,289,3151,2631,3447,414,4130,436,4050,3879,2055,4602,-154,2700,3266,-281,-673,-625,3596,-3535,826,3437,-663,4475,-162,1242,-464,-370,-4997,-29,7094,1867,5258,2193,-8496,3178,2366,-1922,1446,-1623,-535,4291,8041,3127,-392,2807,9648,3410,4616,-4565,515,13339,-212,-729,-281,5688,6484,3281,3247,7343,5366,-1716,-26,9375,1818,1109,5068,1668,2788,1101,2111,5883,1055,1768,1522,7231,1846,3149,-719,-2115,6396,1162,745,3208,3649,2404,4543,-6542,1079,4995,-4560,5527,9643,-470,-3286,-858,-1074,-21875,2286,-3601,-23,1358,-7485,153,1774,2741,9458,2917,-1988,-3562,-5517,10429,-2491,-7402,-1594,1403,-729,-5327,-8349,3183,-1326,-3361,574,-3286,-6030,370,-1420,-9951,4309,-14521,-52,841,-1861,7504,-7973,-7739,-7387,7724,2312,5395,-9833,-18945,-12509,-166,2286,-1457,-5786,14951,-3757,8364,-7983,1556,-5341,4,-11123,4296,-8120,-204,7592,4399,3991,-792,-77,10273,-2524,4086,-15410,-461,-59,4975,-1122,-9458,15781,-3623,6347,11044,-7412,-15322,-3632,17304,-445,3737,-5629,2658,-2047,-3398,8115,5825,7622,-675,10546,6401,-2573,-6279,-6923,11103,-494,-703,-319,3515,2600,-420,-4921,8354,5620,3232,6870,4868,-1406,18437,7319,-98,186,3469,1853,3142,1481,6479,-38,-3476,-2434,1702,4794,2252,9965,-1175,2995,12021,-4233,-1672,-5703,794,-4423,1258,2636,3527,941,2435,-3107,-1550,13789,607,-3149,6313,2719,2983,784,1027,759,2276,2408,-4416,-974,-2966,4504,-4252,-2015,4345,-4697,2807,1041,-2041,-4013,-494,1074,417,-438,4328,4731,2309,1018,-1160,-8315,6250,-5292,6181,1175,2126,8164,-6113,-933,-2785,2238,5634,-1815,316,-3430,4282,3740,-4252,7285,-7177,-1634,11044,3969,1141,-3781,8706,-549,6459,3884,7895,13300,-5200,2319,1429,15488,8696,-1247,13837,942,-2795,-2797,12744,1838,-3081,-7641,9145,629,-3159,-7407,621,-2154,90,-1905,606,996,4821,2812,-2775,-1730,1378,-4489,-2006,4833,8720,-3134,7954,2675,4470,4206,-2194,-4472,5410,9663,3317,-4516,7788,11884,14414,4094,-4443,4238,-13691,2100,-7241,-2335,4450,769,3305,-2008,-13691,-2949,433,10781,946,6630,6748,3305,10058,-129,8251,-3454,8271,-1965,-1950,-427,10400,9799,-7758,-12929,3010,3288,9189,-1560,-9545,2614,2617,9423,-13574,12275,2420,-6103,-8735,715,9355};
    Wx[86]='{-1188,3090,4682,125,-1761,2448,1728,2418,920,3261,-6420,-1583,-3864,5483,8383,-1411,7216,-354,-2083,2319,-488,1821,-128,1960,-195,-3500,-2377,-824,2878,1857,675,5249,4550,3596,-3217,1510,4780,-1683,1533,5805,-369,48,-3959,3459,-8334,1635,-3889,-3276,-4204,-337,-259,665,-1740,-466,-1734,-6215,-2731,-2117,-127,-4958,-3747,475,-2963,1387,-622,-1949,-966,-459,-3322,-4111,-1917,-2731,-3361,3271,-588,4226,1328,-483,175,-3803,512,-249,3156,4760,-4162,-3090,-3398,120,238,-213,-134,2391,1972,-3354,10478,-4326,-1048,-814,-1267,-4108,3476,-1425,-4428,-1604,-2785,-3461,-4633,-10029,-4426,-6528,6069,1162,6166,1904,-21757,3952,-4670,-4345,-860,-1293,3911,294,717,-223,1755,-1706,-641,-6640,-5874,1501,-5703,2274,-1474,623,-1502,-5751,2724,1713,-3479,3481,1612,-11708,-4973,2430,-8110,-2291,-679,-843,259,-635,-862,5375,-472,-5639,-8852,3132,-3371,1373,-8432,2062,-518,171,-1379,2519,-17128,1505,3024,3120,1771,-1845,-3637,10429,1734,8437,1060,-6259,10546,-2517,1893,2551,-9306,19003,1566,-2232,-2805,10117,-4416,4111,477,-58,-5610,2687,10292,-5444,-1655,-485,1477,-15302,-9174,299,-4074,3740,1192,2883,3383,527,-5156,-8896,-508,-362,3659,-35,-442,1155,-6367,-3767,-6166,3601,-1746,-4770,1165,-1745,-3715,2386,2409,968,19,-3125,-2902,-49,4135,3427,1431,-491,-1370,3813,-2963,634,7192,-3527,-463,-9536,-1352,-3881,-4111,1860,-4331,4235,4348,4130,-184,1362,-154,-1695,-2054,4086,4282,-5249,214,2888,-1492,-1062,-218,667,3859,127,-3820,5576,-1619,-4206,1236,5312,-2481,6743,-1881,-6621,-11748,-610,-2019,2352,-273,-4682,-1341,9912,3247,-8642,-4,-203,-1782,433,9189,7192,-3713,-811,2626,-831,-1856,-945,-7871,7182,2990,-929,1190,5019,5214,-3081,-2268,3300,2717,5698,-637,-4606,-715,-156,-7402,5415,2565,-3610,4570,-4638,9638,5234,2048,3852,5449,737,-2209,-3315,-10283,889,281,2393,-707,2875,1436,3659,1359,-813,2797,155,-1674,-5878,2209,1904,-3491,2459,2658,3986,4846,-1882,-442,3737,4311,-7944,-3420,4172,1071,-2995,1158,4321,-2517,-2327,7631,-772,-1582,-4475,-12197,1539,-3432,494,-2463,-480,-10458,-3559,545,-1002,-7514,-364,-4975,-4179,4711,773,770,8437,848,1018,230,2393,356,-5131,867,1032,-2568,-15761,10556,-1633,879,-3815,-5766,4960};
    Wx[87]='{3398,1440,1127,-91,650,-1536,-7763,-612,-370,-82,2163,887,4372,-2412,882,6162,-5322,-4355,1099,2712,1966,-3210,-4140,4291,-3220,3669,-568,3793,-2468,-3840,772,-2377,3083,1,7280,1588,243,2810,3959,-2917,-1202,2670,316,3808,3176,-4291,2409,1634,4650,4023,-2398,-531,-3981,3305,420,-2819,-1689,3483,-572,-5361,1206,1572,-1267,-850,851,-1303,-285,11406,3344,-2744,1395,-315,2734,-258,895,-2037,-1992,-4555,3703,358,-2459,3066,1357,5981,-3461,-1984,-747,-1108,-1300,-175,-4702,3991,-1181,170,1295,4926,-3527,496,-897,102,1427,-19052,-153,2453,3068,-249,24687,6508,289,4460,15791,385,1861,-11484,12021,-1557,-6708,-1206,3344,3,-510,2653,3745,5092,2944,-4177,-797,-5434,-6528,-2452,405,1278,-13476,4948,4707,-3964,7553,1462,1441,9643,-1562,-10830,-1588,-4235,115,11884,-7998,-101,-5854,-2585,19599,-867,-9106,4477,9902,1662,-2905,-5346,10175,1671,-5205,6308,-2768,3095,13994,839,312,-8193,-1651,-361,-108,-683,2976,1402,-4338,2680,1887,3972,9697,1956,-10761,-9326,685,-7197,-1491,9130,-687,1380,7475,-2481,12285,-10087,2456,3305,2358,3955,-8437,-8789,-2066,-2517,3740,-972,1181,3190,850,-855,4641,-3867,1966,-2854,-5639,56,-231,-2095,5151,3315,11503,5048,-1643,3613,2731,-2093,-3029,2044,-2230,-3669,-2902,2406,4343,3464,3437,593,9516,-4860,-414,2136,3234,-1535,1329,-873,5043,-646,-10292,-1678,-408,4558,-6289,-1213,-1259,1529,-9213,1704,-1601,539,551,-7578,-1423,614,5332,-632,-3059,556,-6645,4624,-1157,-2839,1791,-6772,4948,-3796,-9057,-3447,1682,2670,338,9135,8237,2844,-4997,6132,1809,-3518,1409,-650,-1485,1222,107,-1645,60,-2646,7387,-939,5756,-1632,3261,3022,7543,-6728,-4272,-3251,3623,-60,5292,-670,2471,4035,5078,-8012,2043,5771,-2565,-4284,12158,-8486,-1383,-3818,-494,-3234,-4638,7187,1849,-1998,-1453,293,1137,-535,-8745,-1150,7329,8056,2551,3649,2817,-5810,-8085,4274,-7656,1696,3022,343,2563,-7153,1849,1150,-4182,-7583,174,-2985,2303,932,7138,-4208,-3813,4709,-11230,-6440,-1719,9414,6977,-7294,3308,955,11240,-3054,-8085,345,-7250,-3752,9477,-1518,2873,-4641,1456,1606,-4245,3518,3906,16,-661,791,-2709,-13593,2083,8754,-4028,239,-5917,-438,3876,12441,-647,-1853,-5024,579,8950,6875,-2680,-4880,791,1501};
    Wx[88]='{2800,-3378,65,-1748,-2604,1669,1877,1329,-856,115,-3159,1519,-1369,-5419,-1586,-6533,2634,-1289,1287,678,-969,-739,3217,1794,-5073,281,-80,-2834,2749,-3383,-901,-8291,6416,1397,-3381,-5019,193,3400,-593,3059,561,-161,-2036,-11708,-3100,1947,2819,-3952,-1093,1956,-1568,4628,333,-654,-2858,-1564,-3610,-492,-723,2565,726,-2421,2073,-1668,-2954,4558,-4162,-7124,-1040,1212,-2243,-5170,1667,-5976,736,2292,-4487,-3505,-963,-1649,-808,4089,-3173,2680,-1660,2003,-1275,-1220,1676,544,-5908,-4099,3679,1982,1793,1130,-6914,6679,1854,-4138,-1292,-7451,-30,-2907,2785,-27,-2067,-11025,4033,6132,-905,-1552,2124,1707,-6699,2817,-9248,189,3937,1781,3940,4204,-2521,3496,654,-1026,2626,-2338,-7285,6411,-9296,-7495,-2524,670,-2624,-4431,-2790,-1744,3146,20546,-12480,-1154,-1853,1324,-10185,8403,-12089,4555,2352,-7939,-611,8496,-1677,1420,-2377,1385,2312,379,2458,-1604,1916,-7290,803,-2927,-2133,170,-1512,2666,2790,-2919,1798,-6450,3413,8100,-119,-8486,-1196,-8007,8300,411,4816,-7016,-2471,-1267,-1485,-1484,1450,655,3366,5541,-1159,-4587,-4267,-2475,-5000,8320,-12314,4296,2441,-9082,378,-3581,-3476,1102,35,-566,2719,-5375,1464,895,-1575,-3581,-431,-610,5527,8911,-4357,-3361,-4555,1051,-569,1229,-3872,-2148,-274,3486,-1236,2770,-1945,-2177,-2988,1330,-12724,4770,5390,4760,-4423,-645,3930,-1456,5458,3005,10058,6494,11875,-5400,-5473,-358,-4008,5288,-6074,-3508,-4406,-7036,-431,-216,-2016,597,579,-2371,6948,-1845,1072,707,4357,-2275,-373,-10927,1530,-2352,-10029,6401,5395,206,-860,1243,8393,1983,3916,-4338,795,-1727,-1044,167,3435,-29,938,-7978,3701,4343,6323,-689,1204,2644,18925,5429,-5468,4482,-2563,1915,-3154,-1085,-15400,-1735,1455,-13886,708,-4562,205,4116,-3286,-1368,1768,-7700,-3222,2539,3581,3542,2160,2792,-5786,1314,1381,-734,995,4558,-4,-434,-1719,-283,-1839,37,-7036,-1158,4147,-720,-245,6811,-1429,-5952,5395,-1172,-571,1324,-156,-4663,-6474,230,-6704,737,-2362,-7944,-11005,-1168,4521,2595,3457,-4555,195,11962,-3762,5107,2160,262,-4411,-8271,0,-10361,-2995,-1353,-3315,-2692,1766,-5014,4167,3972,3159,-1334,-4284,-6992,2592,791,1511,-3176,-9082,1202,-3403,-9516,-2425,-4645,3122,-1207,2229,6875,9799,2709,-4868,2824,1760,-3374};
    Wx[89]='{2014,-2607,-1076,5043,1578,1616,-1625,-6420,2028,1015,177,-2464,112,5214,-717,-4140,364,-3198,581,-845,3823,-2321,-1276,-1093,-916,2069,-1529,476,5976,-5913,2778,-3557,-1324,159,-5756,-2070,2839,-3925,-4719,3134,-2410,-2374,971,-3547,6459,-1722,3339,-5283,2244,1359,-4191,-3530,4746,-1666,-1564,-3520,464,-2015,-2827,-2902,2348,1119,-4873,1331,-274,-839,-313,4926,4050,66,362,1291,65,339,-2927,-1619,-552,-3413,3388,-3696,-1151,-2320,345,-4782,-4255,-811,3146,-1456,-2761,-1998,-355,-2460,442,1182,-1799,3535,-2941,3256,-215,-5654,-7221,-12666,1137,4462,-995,-635,-14121,13408,-2047,2856,-7006,-10146,7465,-2432,-444,834,1546,-4501,1234,-332,850,-6679,-3596,97,-1668,-746,-765,587,-2138,-6264,-1334,-2441,-9711,-9072,-7265,4038,-3747,-41,8559,167,-927,-15371,2922,-7167,15625,-16416,-8608,-666,-4355,14,18994,6508,-2196,-7124,2902,5336,-728,1301,8032,-2949,-498,13554,-14794,12138,1104,-2185,1422,-1566,-1042,-4,1905,-6381,1704,-2277,-289,-688,-14443,9028,-7666,-8862,-10937,3452,5849,-1503,-7651,-3378,82,-1763,6372,-4645,-6738,10888,1406,4111,3862,-817,-3212,3537,9218,-6640,831,3127,-4462,2526,3090,2988,8251,-3867,-7753,1743,-2504,5166,467,-4782,-2573,7348,6235,-2413,1782,-1998,2274,1282,-443,2452,-1307,4450,916,2851,-2580,4436,1667,2839,-8803,-4465,-1333,-5957,2551,-2178,245,-2915,-2636,4416,941,-1628,-516,1669,-5302,-8041,2673,-1002,112,2883,1227,-3024,4042,-197,-2191,-1505,626,1658,-5825,-13437,-4023,775,7343,-4865,-307,-3400,2463,1409,-4628,-2558,227,-2770,-1967,-1857,9033,-6665,-6923,1400,-5058,3437,4497,-2073,1400,187,946,-5991,4135,-2436,-466,7734,-2270,-3686,-18886,-7568,-220,-2260,-4025,-5952,-957,7568,-1067,-810,-1452,1898,5034,-6718,-4672,-2393,4863,4267,42,-429,-8417,-762,5747,3186,-1837,2873,-8002,564,2489,762,-4116,3642,-2470,-1374,-7485,-96,-699,1033,-14130,-5864,1278,-4204,-3024,-7539,-7636,-2775,-1477,-4731,-1343,-233,673,-4528,-16630,-3710,-2084,4230,-4301,-5649,-3105,1232,-321,-5551,-3999,5742,1076,-3444,1120,-2832,-5087,-5810,-4250,-722,-3071,-2182,6054,1395,-212,6215,1189,-5634,-4855,2988,-4882,-4284,366,-1051,-5922,204,458,-4941,-45,-5322,2739,-6152,-3122,319,-3095,7812,-2941,-1096,-8481,-302,1861,-1795,-984,-7988};
    Wx[90]='{-272,-3051,18,-451,-2687,-2575,1196,2626,3366,3132,-1827,603,2492,3571,3669,4409,-8549,863,2548,-672,-2432,1213,-1126,-34,-594,2578,2846,1715,6479,-2536,-2368,-6762,-5366,-1614,2619,-1053,577,1582,-3503,-2469,-112,-5117,5039,-5122,8300,661,-60,4653,2099,-1030,5288,-884,-2973,3793,439,-1871,-2248,-1427,-5312,2534,-500,2507,-834,-247,-3596,-3491,1387,-10615,556,-1060,158,-2448,2529,1531,778,-4272,3569,2388,-1940,-1824,-808,-6401,-115,-1411,-5429,-158,-1058,514,2430,-3989,-5498,-4108,2246,-629,-1770,3666,1501,-710,-2012,-1943,226,3041,1738,6513,5805,-1080,11835,1760,-1639,1361,-4233,-2910,-3005,-5073,-6147,16787,5502,12910,3193,383,-711,-3459,6669,-2792,1824,3896,-1507,-2509,-9599,5991,-3322,15136,5087,4157,1640,-1152,3999,13193,14033,-5576,745,-8120,2016,25664,14199,-14609,11132,-3647,-3972,-3049,12871,12021,-2093,35,-1417,-2049,-1845,935,-12890,5249,1690,4980,19853,-1062,-12802,-565,-5668,608,-870,-1785,321,5175,-126,-3427,5195,-2604,-7709,3068,-321,3916,1660,-2807,2929,270,-3400,-10634,6621,-76,-2349,-4689,3298,329,569,832,6816,3120,-6884,2492,160,-11142,62,8110,501,-682,-797,459,-3530,-7065,3522,1129,-4042,-900,275,-3312,-3737,1890,684,-3955,3222,-3696,103,-2016,-376,-1569,828,431,-4655,2834,-9433,290,663,153,986,1619,-4899,6777,-1302,1190,-6425,2636,-2348,-7104,343,-680,-2687,643,8222,-7597,-2568,-1384,1527,-3566,1625,401,-446,-1071,8925,3601,2435,503,-2924,-698,-4079,6904,-5747,-2980,-1244,-685,-455,-870,258,-1888,3857,4990,2634,-1334,930,-5874,-4670,7797,-1933,4958,-2388,-3466,-6142,1398,1301,3425,1186,-3044,-1429,-2631,-360,1001,6499,1260,-5595,3383,2609,-4645,273,3383,3618,668,-840,2690,-3925,-1251,3088,9819,-5561,1614,8217,2915,-3344,2756,-2398,4694,2404,958,-219,-961,-1876,-2092,-2292,-5908,-5439,4812,1647,-1480,-5449,2880,-5229,924,5053,-514,-1037,4020,-1988,-5854,632,-7885,-236,6625,6645,490,6914,-4455,6025,-1013,573,-1513,5820,-4724,-1528,-5576,-1072,6791,3659,7421,1701,4770,-1759,-416,-1416,-8120,5195,-8359,10253,3317,1287,-3586,5229,3425,8295,-1097,-8027,4584,-4519,2602,3879,2342,260,1695,-11259,5102,-2890,9072,-2290,4221,1336,2976,-145,-1121,-965,3244,-8984,-2156,-223,5390};
    Wx[91]='{-883,-6015,-10468,3513,36,1048,1828,-10185,-2139,1887,4829,4978,4924,-1612,5800,-3664,2128,4609,3520,3984,714,209,-7421,518,2010,1721,1389,1478,5556,1357,1839,1976,7612,-279,-2398,926,-2788,603,-478,3942,26,-1051,-5185,853,3249,914,-1973,1705,5107,-139,1082,-655,266,-200,-5825,-3325,-2868,1745,1063,-2663,2291,4191,-2291,-728,-1870,-957,1168,-3015,-1448,650,405,5346,129,3032,-1081,233,10390,899,165,574,3767,-2822,-3361,-2954,3134,10566,1959,-94,2359,-1782,2604,-3310,5034,-1343,-2397,4038,-1796,3708,-902,2849,-1628,7641,3613,311,-282,-1147,6484,12207,4614,-5214,-498,-2322,4189,-776,-11640,-20000,2890,2597,3139,2731,-5073,-3015,10380,-3786,-690,720,6079,-2934,-463,10439,-2453,884,-365,-2661,-1522,4309,2423,2687,2489,-9726,4626,-6611,-5234,9545,-12021,1944,18906,-2022,6098,-2326,10322,-11103,1512,-9213,3405,-794,5600,-510,1856,-3037,699,-13193,3854,-8251,2636,-2257,-2254,-11611,-1358,-2741,-2441,-4536,-1290,-2546,-3342,3923,3161,1666,5776,-2626,-3217,2954,-8769,-15781,-732,3571,-2885,-12480,240,-8271,-343,6791,-5664,1647,5708,2568,3125,5561,-4401,-1557,6601,-2104,-5361,134,3911,-179,1007,10605,-2087,-477,-3618,-2687,6264,-10947,-1022,2171,-12382,2844,-1907,1976,-3146,-1330,1300,3039,2944,-1472,1856,2479,646,2792,-1101,-5966,875,-3044,4389,-9116,-29,-1967,-3198,-7080,1638,-2231,-3876,-1724,6035,-603,-4421,-6948,-2534,841,-2585,69,-539,5498,1276,-1883,-5654,6538,6269,-1025,-3371,-4719,-3581,-1932,-2409,-1695,1923,-834,-2073,-1053,5190,-8305,-1602,-5400,-1492,304,5786,-1600,72,-4020,2609,680,-5571,6879,661,-3144,638,394,-4497,-1617,4633,-7041,-10917,-102,5107,167,2861,-10048,449,-3361,6206,-2619,-3117,-1207,2210,7021,-5375,-2807,-338,-5986,-6909,288,6440,-8247,-6411,-712,-81,1817,711,7094,4560,-3022,2456,7758,1999,-3708,960,7534,6235,2534,-3156,-4645,-6684,-1790,4331,-6660,3393,6137,-2482,-1597,6298,-3105,-4631,-14375,-4843,-5976,-900,-3449,351,-1192,354,-2393,-9208,-5937,4382,-3735,-8173,6215,-248,-7749,1973,1397,-9169,6093,-3085,9941,5258,-4912,5244,1992,-8310,-8247,12412,-2973,2775,-107,6489,-8051,-1014,385,755,-3889,-3063,-2141,13271,-10322,2661,-3298,2181,8203,4284,-8378,-8774,9243,-3962,-510,9428,1654,-2858,-262};
    Wx[92]='{881,-6499,830,966,-77,-1246,4479,366,4372,1365,3493,424,-3410,-5727,-2403,-1112,4680,2995,-2274,-2279,1512,2795,1439,1036,2198,-295,277,218,2115,-2927,2456,-6508,7563,2224,869,498,-870,3317,-5053,1330,-746,1375,-3391,-204,-1954,1317,-5083,-1918,568,-3894,-6875,-402,-1624,-1590,4211,4233,2026,-6640,-314,10351,-7548,-916,-1491,-1890,-2108,-870,-155,-6835,-5590,-1605,-786,-2453,-450,-1738,1425,-745,-2148,-3779,-1196,97,-1143,-11796,-663,3210,-1011,1390,1083,-247,3017,-3481,-3576,-3691,2416,-323,-717,-2089,-6357,-1205,-2305,-2001,-1073,432,-5693,6977,2878,-731,-8735,-5410,-3156,-4616,-1748,1612,-6420,-2656,-7202,-5874,1225,-540,2467,-5239,385,8872,3408,49,-1336,-5507,-1340,2260,6005,8618,-5253,-10927,-902,-14013,9497,6,5126,-2254,7470,8852,2795,-17675,690,3623,18183,-167,6201,-16894,429,-8779,-5107,9521,9462,-4487,1401,8071,1892,6835,1561,2783,11396,7153,-3444,-5795,541,3122,-2219,4365,4484,-667,-14833,219,436,-12304,-1949,6264,1422,2761,-10087,2370,-3657,21230,-1853,3874,-5673,5942,-2524,4951,-656,-5522,3232,-3920,3500,-3093,-19902,-2507,-4020,-4912,383,7651,4150,7456,4372,536,5781,-351,-1249,7407,1492,654,-642,-2207,2083,2792,-1268,-8173,-9863,-4736,-1555,-3342,879,951,98,-996,4462,3530,-3188,-2851,-3559,5961,-677,2274,996,-2717,-2010,-766,53,618,-674,-514,5268,11376,4331,-1550,10400,-2597,-1507,1759,3989,-310,10722,2048,184,-3847,-5375,841,2666,-4140,-2558,-10673,-3710,4685,3891,-412,5952,-1231,-111,11152,-7299,1150,9936,1378,4924,2680,2963,-300,-4216,1690,12695,2946,-4003,4619,5512,4216,3803,-3222,1126,-891,470,-3320,-2335,-2437,-1472,4489,1878,2471,-3981,-824,4970,5200,6533,5830,-1953,-767,3935,-1804,-7563,3408,43,-9326,-1027,-549,-4980,1622,3061,3149,261,-5761,-4772,-2122,3244,822,-3115,-2239,9355,-6469,851,789,2546,6010,-2639,-32,-6401,-5273,-3015,-1818,-3229,8266,2548,-1486,955,8046,-4165,-6308,-271,-6567,1307,2044,3469,-8056,-3059,-8041,-4921,-8164,-8081,1622,1658,-3149,-4584,1584,-1545,-1947,9370,794,-3505,11220,74,259,2712,7724,-2524,-590,-1304,1832,-2150,-3505,-6928,-4238,-2108,1394,-3547,-1920,-2915,1904,554,2902,-50,1577,1527,-4357,-7773,-13046,6640,-6479,758,-2983,-3103,10917,2773,-6728};
    Wx[93]='{-946,1133,-603,1163,2453,-1799,-270,2880,966,2324,-1215,494,-1297,-2124,-160,-3210,-6826,534,-3994,-4567,1483,2113,4565,4055,-1259,998,111,657,-1463,1912,363,-3405,-717,-3071,2500,1117,-765,874,2344,327,1074,-1430,3403,303,-3359,2216,-6855,4155,-12,-930,12275,1287,842,1741,5571,-2541,418,-1301,-166,-1614,832,-3959,3527,-2194,-3918,2573,1416,186,-3698,870,-360,-4091,-2276,-1588,1629,2548,3962,2734,3935,-3137,2570,1131,3840,3601,3830,2279,-263,-1881,2739,1488,-4028,-464,1785,-4934,5629,-3564,-2221,-6210,1876,757,143,711,1431,4904,-3386,2626,2393,1282,4221,-1689,-6323,-38,-3298,3332,-8310,-1165,1597,3991,4501,-2685,779,8208,-5449,-2445,-3530,-443,-700,773,2236,4997,-1729,-2727,1741,2073,3894,-23,-667,-184,-134,3398,6796,1000,5498,1287,-2966,5463,2976,-6840,-1258,3674,-3999,1359,16416,2907,-6435,5898,261,1694,1748,4052,1282,-7285,-12431,-1345,-5527,-1711,3366,-9604,4655,158,-13828,-5859,-798,676,3798,-2751,-7700,4602,-6577,5136,1490,14296,586,-8647,4636,2580,-2980,-6582,-4418,1815,1834,-5170,1199,-2514,3400,-2406,9916,3876,-3967,-2526,2174,5229,-267,-692,2961,-1092,4721,-3234,1545,-780,-4882,-3159,-1434,-7314,5498,3771,-5712,1837,-1745,-2205,-794,89,-1904,1113,4379,90,-5693,502,-1210,-2878,4006,-6391,505,3671,-6503,-1306,1630,-5097,3435,-2429,-5019,-1278,5288,-1662,1428,-4101,2519,-864,-4519,-1433,-7861,-9794,7250,2331,3374,-4514,602,-3979,349,1000,-2355,-2802,1730,-230,3186,-508,-567,9477,-3764,10,3835,2015,-3903,-40,-36,-1232,-6889,-1468,906,-849,1132,-5795,4895,-3630,-1959,-5219,-26,-772,-3918,-254,-3227,-8818,-518,-1237,8427,1875,-3308,-924,3027,-3181,7797,857,-49,2149,3491,-2617,-534,615,6240,-520,-2032,3803,-473,-9531,2541,4523,1373,-3125,-3847,-3078,-2114,-3569,2412,4653,3847,19,-82,2432,6093,2069,2993,-3847,-545,297,-1839,-2115,7988,-117,5834,-4260,-2551,1785,-4025,-6640,-1207,2464,805,4228,217,-3344,9189,-4670,695,487,5419,3789,-3112,-1313,-1019,-2883,1180,1345,664,-991,-1429,3698,91,1198,-7485,-6118,2949,-6157,614,238,2805,4677,155,3586,2727,-6499,2890,-4536,2290,-3112,3132,-9804,-1006,-1071,1066,532,-6630,-4819,2834,-7314,897,2912,-6542,3266,2937,-3950};
    Wx[94]='{1278,-1942,-554,-3161,2247,-1317,-3459,-257,4523,-1707,53,290,2734,1262,1688,-38,-210,2218,3183,-1376,603,-3034,-1348,20,3537,-789,-402,3537,-47,917,-1695,1552,2556,2216,3493,-2685,-449,-341,1828,98,792,32,4956,3322,3239,2700,-1190,-3005,755,1495,-3547,-6298,-257,3027,-3793,3896,2218,-2358,4189,8681,-214,-3745,-4965,1915,-1173,-2753,2130,1940,3312,-1597,-1844,-5380,-816,1743,-3994,1408,-4055,1503,1008,4018,433,4721,-1651,5737,-1200,2248,2397,2922,-297,-3989,3413,-4980,-3823,1297,1866,1730,1078,736,1713,-2617,4973,453,1364,8989,6445,1612,-969,5092,-5922,-9291,103,-2360,-3569,-6923,13505,-11572,408,-82,-3020,-3884,-4487,-9990,4094,-7744,144,7685,-1816,-4265,-2790,2905,-223,15332,-12841,12353,-692,8701,1850,4011,-1209,-6567,-4802,19033,-662,4726,17626,3452,2395,-2641,11064,-3154,1138,15078,-2189,-10781,5415,-2956,1614,-2770,-12968,-2471,-2812,-1461,-5839,-2237,17255,1453,-1450,1614,-827,-1997,236,709,-1233,8813,-3725,9628,5830,6367,-1514,-816,6186,-5864,5991,6982,-2617,-7524,3007,12080,-578,-2189,2663,16572,1363,-506,6953,4826,-4067,-1607,3447,7700,985,-2744,5078,-3874,3183,423,690,-1779,5000,4111,-7021,280,1402,2707,4316,2800,-2156,-6474,-936,-891,-1857,2624,-1557,-1411,-1977,-4519,4641,44,8,-438,-2385,-5405,-8754,918,-3405,2448,4362,2424,-2922,4165,-3090,1148,-3151,3540,-6850,-3417,8378,-241,-4323,-2318,5336,-3940,-1689,-5800,1884,618,-87,2717,1844,-7587,-7377,-586,-2281,-8422,109,-3581,-2441,1976,-3718,-820,-3295,-3225,1063,-5170,-770,2927,-567,-752,11660,-568,1939,985,3256,-3344,4055,-8,1651,-2509,910,-1806,845,712,-5683,-6611,-440,-426,-2167,-3405,2178,-232,5751,-6254,522,-2495,2077,76,1253,-5117,3264,14023,-3481,-2164,3020,-1354,2658,1301,-3076,4116,-324,-5600,1781,1573,-8471,-1589,4223,-7514,7495,-1718,-12285,-4584,-4162,-7880,-5830,-1463,-1781,1916,5131,3037,-9091,5400,778,-5297,3835,3093,-1342,-3950,341,3691,-1328,3144,-4970,-4313,-5024,-1060,296,328,-623,-5961,3669,-14560,-3767,-1231,-260,-8764,-1912,2331,-2812,-1763,11552,-9233,1008,-8500,-6181,4553,1287,2504,-11914,-4079,5,-896,6542,-6176,-529,-4272,10000,-6098,4975,1499,-60,-9023,1569,-2675,-7221,-5488,-323,893,2364,-3098,4536,573};
    Wx[95]='{1154,456,1268,1986,2487,484,2968,1955,-2700,-1417,5942,1501,2646,4343,4467,4575,2619,-2125,1177,4423,-652,2768,1036,4079,977,-720,557,-546,11582,-5864,-478,11894,5527,2731,3979,2132,-3937,1135,1611,-1981,2193,3090,-1610,4265,-4750,2071,5078,-11,3173,-126,-3273,-2187,-1752,2731,-1800,-3225,1014,76,-1761,222,3991,8037,2934,5991,-4020,620,-4101,4255,1254,-662,-2243,4118,-1354,-223,1119,817,5781,3427,3359,875,1040,14238,7490,-4243,3022,8159,2078,5053,3161,-2062,-793,6816,5131,6201,2573,2270,1687,2875,2388,-1205,-5039,-6816,1176,2352,1768,2443,3720,794,4851,-230,-5898,-2687,2387,8237,7563,-5498,2070,5146,2404,1857,31,834,1510,-1380,-4692,-2795,1093,667,-4152,-5,232,-11923,652,7690,-2181,11123,1075,4028,12089,-11777,-6538,1205,1843,-4987,7812,-6025,-4633,400,4868,5820,11865,7680,-6035,5678,4160,-4052,-3022,-1103,10859,-3542,-321,18486,-4760,6318,8110,-2941,-2093,8486,-3608,2021,-637,5336,-1804,2132,2968,-9047,3339,5073,-3857,-3127,-6035,-15634,4313,1633,1997,-5615,2199,3122,-3286,-1113,-3251,-1630,-2832,553,-873,8642,-3381,1968,6347,-911,-4160,-2836,941,5312,-1170,928,-3735,-2573,-1927,-1431,-322,-3059,-3093,3413,-3962,-3845,-1783,-1801,-1597,744,1585,1356,-2644,-2218,2059,-2283,5151,2958,857,8291,125,820,929,2210,5512,897,-526,2371,2196,1541,-2205,-5117,-472,9150,1571,-1976,3269,257,-1133,4060,-2424,1199,-2283,-4038,-1529,-1455,-6748,2130,5815,-4372,1136,3322,-513,-5629,6093,450,1395,10351,-1005,-263,4277,1734,2076,992,2443,2207,4978,-6430,7915,283,1978,8471,3937,-6538,4296,6547,-1485,657,2419,-5507,-961,681,3107,-504,-4191,-1273,5034,-3715,3405,-1072,-5644,2270,5107,-2993,174,-738,-567,1032,-3737,-3217,11269,1427,2250,10283,3520,-1223,3430,6186,-4709,7387,4960,-3178,-2261,3371,-4677,145,5502,3688,9169,1954,2536,4895,333,3625,1320,546,96,-1307,-3298,3654,-3442,75,596,3076,6230,-1224,-562,-737,-6411,-240,-3820,-1768,1884,-6220,-2277,-6142,-5449,9667,-386,-8999,637,5380,-4160,1087,-2167,4208,3793,5395,-5205,3554,-2301,1928,8789,-5039,6635,5742,1044,-89,-750,997,5634,230,2059,-6259,7695,1888,2207,1911,-2583,3122,260,1068,1282,13134,1628,93,6806,3405,2143,-907};
    Wx[96]='{-952,-673,2875,2812,1784,-1928,-3164,3093,2541,-178,-919,1201,237,-1749,100,7221,-299,1190,-5742,3669,-3493,1835,-2167,7651,2117,2215,3325,-940,980,-6914,95,274,-5454,2282,-88,1452,-3901,-2368,440,4672,-1342,1021,3740,-1611,-2064,-5385,-7294,2145,-4094,2227,-2800,-1674,-34,4602,-2026,-2143,1354,1133,-1345,-5600,2468,-3723,-2352,3112,5732,3400,543,4516,3481,-160,3125,-3127,-3134,-2122,877,7675,-1157,-2116,5078,-4199,1954,-7426,-672,-585,-6040,-6284,-1169,699,2109,-232,-3303,1785,-2675,-3132,-258,-1823,239,-708,-150,-2612,-4855,-2783,-4025,4802,-1381,-2149,6997,4462,-1533,-259,13955,6342,4863,2006,4658,3955,1677,5083,-2072,4768,-3916,7065,-7358,1079,-1782,11503,-2236,-2197,-2106,-2432,-4462,-2646,-15517,8378,-1400,5917,2863,-2919,-7211,-2724,-6083,-10605,-1018,-1524,-2380,2435,14140,6015,4301,4343,-5014,20761,7431,-4077,428,9838,-5493,-1475,-12158,1650,-4213,-610,-1582,4599,8310,-4287,1434,-4582,1127,-2526,1486,5893,-2014,3500,-7148,-255,-2430,-5664,15029,-1563,2354,29726,646,-8750,1502,-12910,-3974,1347,-4355,5551,-1859,13818,-3593,1463,3005,7446,5849,-9863,-1431,7734,3881,232,2746,93,5966,-1007,-465,-8115,-7026,-3742,-6308,-4558,-845,-950,1215,3647,-4536,-2519,-2133,-125,571,1535,-3483,1815,-1265,-5004,-4277,-1613,-3056,7016,2413,2263,1875,-4799,2423,-665,-2990,1916,-440,2846,997,-1549,-8330,-8315,-2644,1375,-5532,-1928,9067,-418,-762,4252,177,-4025,-2283,4267,-3449,-1171,-2437,-996,5751,-8935,-967,2661,6674,-1524,155,1079,1365,-3073,-1422,-994,-919,-1149,-4653,-8588,648,-6425,-6791,-386,669,-4560,-4453,-897,21,-7851,-1566,-4067,-2919,-1182,5205,-1682,-364,-664,823,-2858,5317,1901,-3815,-4597,3166,-9028,-563,-6704,6074,-6694,-725,3642,-2968,-2939,1733,-3186,3706,-8134,-3566,925,-8476,-1583,1102,671,-6230,95,4250,6240,-355,6186,-1440,-692,-1921,95,-106,-5791,-4548,-10781,-1888,-2675,-3056,-4313,-4799,4987,2646,914,5688,-15644,-8886,1531,-1452,1166,-1073,-930,-3337,-11572,-2255,-880,1967,7646,-1192,4311,-2160,1766,5449,-7714,-3320,-3735,2177,-7182,2666,-5312,-4904,-1866,-2307,-192,-839,-3225,-3041,-1793,-3732,-9995,-3684,2292,1303,-7265,6914,-3090,-2624,-1568,966,-3237,-625,1511,-2307,-7680,-4990,5429,2614,-8686,-2619,5493,1429,-5161};
    Wx[97]='{3718,5190,1887,-1628,-1796,-2110,1901,1026,-2890,841,4128,-605,1130,1325,2277,-1851,7124,136,-78,3039,-1431,-3261,-657,-370,2326,-1536,4650,1239,2276,-1745,87,7631,-1069,960,4973,1124,2709,4272,2814,2467,1699,-1773,-266,6386,-9995,-4685,-1133,-321,-3061,-605,-292,-4450,-4868,-2277,3103,3947,-1860,75,-1248,-1978,1095,2575,151,-3911,-5058,-3376,1370,1005,-2619,-2634,692,2805,5463,-3452,-1910,2736,3,-1606,-2066,1501,-1497,6894,-1549,-3320,-957,-6357,-2949,-674,-3339,524,-393,2822,-5952,-3671,-538,2150,1195,-2634,-2995,3208,4140,9384,-1408,-637,1227,2041,192,-4924,623,-5249,-6323,422,-2746,-3049,4414,-7568,5009,10400,-1330,1833,-4221,-879,4091,1870,199,3676,-745,1197,-16318,4521,5947,6630,21601,495,3103,2387,2749,11582,3247,-9091,-9936,65,3657,5434,9663,9604,3769,-11621,-8183,8305,11669,3093,-7021,10205,933,-8701,554,2624,6132,3916,-5122,-3374,1021,2180,-1942,3630,3027,6831,-2194,-877,12832,-4401,-1375,-7592,-961,7783,15859,-2819,5039,-3635,-7299,729,10078,5717,4741,-5917,5551,332,2318,-563,855,-1958,19619,-1345,-9091,7133,-6845,-15527,3125,-7021,-950,-1113,1445,3381,-2174,-2120,4340,-1114,1658,-3496,1674,4775,-5678,592,-4709,-3015,2817,4667,7709,1660,1403,2741,1303,428,-1092,-675,2066,-2077,5141,-3527,656,-733,4802,-10429,3483,2998,-1190,3010,-223,2695,-1231,-7148,-2347,-1947,2125,-1547,10410,1469,-2797,3894,7329,4919,-298,7631,-1363,-5737,4216,4853,-6801,-2360,479,3659,-3735,-3547,-473,-4770,-2976,-5478,-4111,-597,-1881,-1501,-277,-943,-843,4328,2200,1820,7329,4047,-1179,3017,1194,3530,-3352,-312,-847,3356,1629,903,-6679,6030,2319,2919,-3930,881,-9462,2204,-2988,314,-2127,1761,10478,4187,-1043,-8066,4238,917,-476,-1884,5502,-691,2639,5175,-3916,-1914,4807,7988,-5810,-574,2274,3569,-6098,-2021,-471,2841,5844,-1499,6157,-4196,617,-2213,1602,-7460,7529,2290,6835,844,1522,-1663,-644,-919,-4816,6992,3195,-4550,-2033,-6069,-500,-908,4108,6630,-279,3991,11552,516,2110,-5795,-2166,4230,4797,678,-4914,2198,2016,365,-5864,6069,-897,-8061,-7680,484,-3771,404,392,8896,-210,-974,-863,5131,-5136,-2198,2587,5527,5600,6494,-1436,4694,501,663,1492,599,-3112,2863,-57,4719,-7211,2556,-3859,3713};
    Wx[98]='{87,-5517,-1716,991,2712,2304,-54,-6552,-1965,334,1790,-1761,-1981,-1112,-4191,-6542,403,-3342,-1156,6225,1351,828,-242,3237,-2814,476,2322,-405,-718,-3129,-3833,-3212,-1466,-2536,-2027,-1280,-1595,1851,-1979,-2631,-1455,-2519,-2077,-6171,-5322,-6235,-1065,-5981,1170,-1447,-4301,481,1678,830,3159,-10576,656,4814,-809,-4069,1711,-662,-1097,-7905,-1110,4428,-1973,-2707,3654,2381,4482,-5751,-2524,2125,762,-902,-3874,-10996,2609,-1534,-5419,-3088,7133,-225,-7001,-6333,-1179,-1866,68,3728,-4130,212,-1236,21,1679,4707,-8662,-7377,-3708,-3693,-1976,5639,3339,2561,2470,-2546,2990,19121,-3598,3649,4804,-1625,1462,-6074,3376,-2678,883,800,6542,8056,-1604,656,-1689,4570,-9448,4304,-4638,817,70,6840,-4589,8334,-24941,326,-1522,4421,188,6708,-1127,23632,3388,4011,-2208,7895,6508,-914,9121,11953,3730,1381,10458,12949,2543,8876,-1719,10722,-2459,2020,-3071,-501,4296,-4409,-10224,10791,2668,-1726,-1244,-23261,-3439,2207,-9956,-3786,-1922,-902,1654,-12519,1743,-1026,3276,8369,79,4382,-4572,-15810,271,7827,-8427,661,-7421,2573,9833,22480,-9433,2093,-9501,-1096,-6210,-10166,-910,-17060,2294,112,-4633,2077,2384,-358,5424,2922,-2166,-4897,-5234,1822,3413,792,182,8510,-6171,-1605,276,2583,-2152,-218,1273,-2093,1536,5473,-3242,3483,-4763,-1567,3041,-5649,-2683,-10039,1751,9560,6811,-1248,4409,4238,-768,6328,3923,-6997,2683,3354,7148,-2338,3757,3940,-4733,1000,696,1850,-564,3996,-4807,3959,-709,3950,-1244,-6630,-404,-8125,-2291,-1904,1198,6069,4165,1901,6127,-3427,-4301,-2186,407,580,3432,532,3823,34,-614,-4208,1979,3740,-1876,-1634,-592,505,-1409,-1909,653,-2366,-1860,-2519,-8491,-7836,3432,-4887,5083,-10048,-4941,-12333,-950,-7036,2081,6772,2973,4147,-4123,-9873,-6762,-3330,8808,-1561,927,-1035,-3928,-9116,-2863,-1157,-1508,-3518,-5737,1082,102,-2993,2749,7412,-5561,-2414,-7373,-6020,-3925,-17978,1225,-75,-5566,4704,396,-3918,1835,19,-2985,-9267,-6879,56,3027,650,3208,-3254,-13212,-1862,-5312,-2668,8320,-2192,-7890,525,-2663,6206,8193,-7187,-1832,-9462,-6137,770,5673,-3840,21210,-1370,13,-5341,3552,-11289,8544,-2382,-1158,-10273,-5610,8300,-2915,-5717,7314,-11376,-2600,-6987,2485,-6445,-662,2088,567,-260,-6220,12910,-7202,-4785,-14873,7817,4604,-6708};
    Wx[99]='{0,-7602,-2697,-443,1141,1296,-1783,-1112,400,415,-2327,153,-563,1846,-5488,-5634,-360,14,-5288,-829,-4489,1727,125,1754,-3996,-1535,-1577,-1745,-149,290,-5390,-2209,-1810,-378,724,-507,1100,1977,-68,-388,-2863,-1740,586,-3640,-2493,-1866,-1348,-295,-3247,-264,-1042,491,-828,-3513,2568,-6806,-3579,1732,-603,-2067,-3486,-2042,126,-1699,1423,2056,-2634,-4362,2320,463,-1973,-8056,-6606,-2125,-747,-1213,-992,-591,251,1864,1700,4829,457,744,-277,-897,-3154,121,-2998,-1557,-43,2521,-366,57,-3884,-1716,-123,-1049,-1767,141,1118,5976,1807,-3088,-10214,-1951,-1481,-1502,2905,-853,-456,-341,4580,6254,-10507,4501,4860,-3969,1982,3044,-2575,-2949,-1315,-1212,-950,-5810,1614,4150,3237,-5200,1518,190,4799,-7358,-4174,-2883,1636,-5537,15019,-4580,195,2744,-3576,12802,-3481,3037,3337,3632,-3820,2687,8784,10517,2358,6650,-5273,-2252,-3146,-1790,2449,-5834,6606,-10595,-13613,1555,10302,-5322,8774,-6010,-5234,-1428,-3239,995,-6250,77,3566,-8178,-2827,-2778,4047,1341,5996,3017,4306,-13515,3991,-2734,-8481,-1158,1275,19,307,-808,-5356,7011,11845,-10185,-2497,1068,5053,2355,-3066,-10517,-876,986,-2038,2141,2956,835,3498,-779,-612,1542,6894,3828,-152,-5883,4260,-114,2690,842,-2568,-3811,2186,-1673,-1174,1539,2622,2656,2812,-710,-1730,-5629,-10605,11191,222,-6035,-10078,-8413,4143,4604,-329,6767,982,11025,527,-6005,17119,3742,3508,3149,2080,11279,1481,7041,2805,8227,-7939,4233,1612,9833,-3659,-1578,7182,-145,8867,-2746,-359,6616,5439,2563,-2414,1064,-7250,-577,-2252,722,2108,123,-1982,-1748,2237,-5493,-2810,3066,-7382,1713,3076,2722,784,802,-7412,-962,-3925,3596,419,1516,-756,6835,3281,3122,-8378,318,2261,-2646,-9848,-274,-2636,-1668,-1524,-2031,-7104,3527,1087,-1710,-661,1892,-1572,-6396,-6606,-958,-12998,-4206,-200,-1390,-4760,-81,1096,-100,8037,-3078,-4267,-1982,-12685,7553,-7758,-6738,-3234,-3127,3056,2286,3625,8627,5556,7514,126,-1710,8159,-2044,-45,-802,-2476,7124,-1854,-1022,7348,534,-8432,1979,4108,3161,999,695,8178,-570,6088,-847,2005,-2585,15849,4685,-6787,-2561,-1418,-2314,-3957,5546,2941,416,-6567,2266,2626,3610,7016,2968,-2287,4069,5957,1622,-2919,5771,-3891,5976,-4685,17724,-7036,4570,2709,3901,2949,4821};
Wh[0]='{-639,1331,3195,1979,-1818,-1262,-5014,-3674,-2246,218,110,-212,1027,939,9321,730,-2362,-1622,771,-3691,2604,1707,-1196,37,1533,-171,-3359,1143,-4443,-1948,-1206,582,-327,3024,-325,-653,4538,1918,146,1809,-4106,1563,-10683,2702,2073,1412,3740,6674,728,-625,-6787,948,3337,-2044,1254,4880,700,2514,-371,-1955,-5087,-2167,-2509,54,-125,-653,-1619,3762,1617,-1341,344,-66,886,1839,4003,-1707,-461,751,-1530,-1618,1468,5327,-2990,2753,-3623,1536,733,1706,-2362,-4777,-2553,-1270,-571,-2322,-2839,-2497,374,4614,-1005,2006,-1992,2205,-2565,3779,-372,1890,-2480,-2985,-557,628,3605,-329,3540,22,3305,-934,-2113,-9125,-1254,-4633,-3681,-1566,1905,1395,52,4841,2489,606,-4311,-3842,-1079,-1669,-3510,-150,-751,-2707,-1834,2174,2673,1483,-6191,965,-4064,-1433,-438,-1629,-1484,3874,-3515,2900,-590,2866,3879,2678,-5136,-4658,-1062,-397,-2015,183,-4951,-1062,3095,4150,-815,3662,4252,-13,-954,-2337,3945,3710,1706,1744,-4914,4248,593,-423,-1060,-219,-1979,-5371,3764,649,2342,660,2841,-1496,-7802,-4592,1066,-680,1334,-3076,-704,-2702,-72,329,-1895,-830,3037,1015,2607,-5849,2590,-666,-1535,5126,2030,990,7050,307,2261,-4904,-3491,-1177,-1842,2449,4504,-1452,2481,-1495,-2473,3972,-339,3876,3344,1536,-1584,3173,2061,-6132,1099,-938,2819,171,-1054,446,-1343,-2900,4309,-3391,1835,-3588,-1284,-4704,-1397,769,-806,5776,-2347,784,2941,-314,-1849,3149,4396,1118,-1662,-662,2832,-2054,563,3115,-2115,-942,1730,3576,2937,-990,1046,878,3962,-1666,549,3356,664,-470,527,-3188,1059,-3964,1763,-3452,-573,-1571,-2939,614,401,-3063,5126,-557,473,2362,-1123,3576,-245,9,4736,-3210,4929,1600,949,552,1483,3535,2949,-2902,-609,2790,2003,-261,-2287,2414,376,2091,-3349,-699,6455,299,5502,304,-3913,-907,5126,368,443,536,1265,-648,2347,-1766,-6059,230,-1511,6147,4980,4731,1163,-1485,2639,1617,-5385,-4829,-6738,-3688,-7099,159,-1740,-250,1582,1871,393,1245,1171,-3242,2595,4182,-251,-158,-3398,-2226,-1765,4042,-1365,-960,3183,4433,-855,2849,-1947,-2033,1954,5541,6259,132,-726,-2105,-1928,-2321,-1396,-1018,1026,-1156,-2254,1234,1253,1365,-817,2915,-1474,4438,906,-2489,-2368,2054,-2452,-1568,2687,223};
    Wh[1]='{-41,-439,-3120,-6069,139,5219,-13271,-5351,-320,581,-5214,6064,3962,-8251,-4792,-1395,-3481,-2030,3308,-2108,-94,1506,2390,-6733,275,-9199,-5810,859,672,-4895,1300,2141,-3911,-4631,922,3476,1683,-985,-1101,2496,-3486,-4750,1383,-9448,-2536,3354,-10781,-564,4035,-3315,1959,227,544,-2512,-7763,-14179,2646,-4597,-3898,8574,94,-3156,-5839,-25,1602,-3144,-3139,2465,-7128,-596,-3349,-5712,1331,6723,676,-1914,-1097,-6928,-4348,726,3425,-6191,-4062,5468,2978,4841,642,-2248,-7534,1535,-5146,385,2839,-3525,-720,3303,-3625,87,-1174,864,-671,-4992,-679,2670,5258,-526,-5380,1005,15136,-5473,-3076,4702,-2414,-3666,-2902,-839,-718,2142,1301,-4057,51,-2956,-876,147,-1152,-5205,-9106,3339,-741,4394,4035,-1785,-4167,1596,211,-11132,6235,-645,-4230,3049,19248,3752,5336,-4379,261,-9243,5009,-15976,-5292,-12,-7124,1700,-708,-1461,-1464,-6342,6630,3188,-1793,-17646,16953,-9169,-2661,-1024,-4172,736,3874,3789,2265,-5415,-271,52,10996,-1489,6118,-4487,4187,-886,-8105,880,-531,5234,695,2819,5205,2985,-2436,3837,16220,6787,6557,3264,-962,4799,-177,12,1116,-1546,-1894,-7167,5092,3232,-1683,5917,975,2919,7324,8745,-8940,5253,6430,-1875,2321,-2082,491,-2385,-4221,-6293,3957,1241,-3129,3393,538,-7656,2917,-636,3525,-2941,6313,7822,-806,4296,2534,2978,2188,-4189,6616,1001,3781,1379,4782,5986,1779,-2927,954,4528,6533,2661,2856,-657,-3632,-1510,-1618,6127,2900,6821,-19,2739,3,-4084,1043,40,23457,-2800,83,5874,4602,-2352,-3881,661,-1842,7954,2624,2744,-5268,125,135,-3308,2590,-2218,3708,2792,4802,7719,1507,2565,-6557,-2487,8183,6508,-1577,-3942,2597,-8164,7216,167,-299,-2875,-1396,5307,4458,2495,-6108,-3286,3435,-5141,-4389,-2539,323,6586,-2951,-1318,-518,-3952,152,-4870,-1253,-5556,4589,-5839,-1931,1701,1732,-4653,993,-4409,-7192,263,-2727,-215,-5766,-2032,-1238,-1876,3859,4970,-1845,-9047,-2763,3735,1286,-5483,-2143,-4978,-6669,4738,6259,4321,1745,3132,4431,-3256,2980,-1467,8808,3442,1693,9169,-14570,91,-5097,-227,7275,-1188,9135,-3168,-9291,3183,-1964,-1502,1194,5615,-210,-6723,-9790,4326,3071,-4775,-3547,-292,3447,7485,-3188,-5708,6333,-1362,-1214,939,3037,8046,-5073,-2226,8393,10068,-3522,4121,-4123,957,-3132,544};
    Wh[2]='{2076,-4062,574,400,-1826,-2153,-3430,3229,-3078,2000,-301,-2570,1149,-2069,-1693,-75,-2034,-3789,-3593,2054,780,230,1251,1750,-349,180,1948,2442,-1199,-327,286,-2749,583,916,-1315,1612,-4606,-3361,5244,3347,-958,-183,-3996,-523,-8886,7250,2122,-1889,-255,-5732,-1914,-814,-1252,-6938,-824,-3913,4694,1429,1293,-6748,3857,-4360,-1030,-5146,909,-971,-2858,3576,-2084,2993,-5605,-3002,-1196,2912,-1491,-2110,4294,-2106,-6835,-1128,1926,4265,-2122,4931,2587,3303,1518,-217,-2148,-3767,1611,2120,-2866,3210,2507,4069,-1414,-289,1771,-857,839,-5561,1128,447,-2194,-318,-4699,-3237,-15947,14072,-10771,4978,-10146,-1737,724,2775,-2751,-12998,7451,-2407,-3676,-2792,2958,410,-10195,670,-6977,331,8139,-2502,1380,-6552,4250,3225,-3413,-5288,-549,-3027,-2690,-111,5112,-1602,7119,4921,364,-2524,-12109,767,552,-2070,-3576,-6547,-2211,-7070,3571,1822,-2773,1423,1464,-1113,4265,-4721,2224,-9404,-1528,-693,2216,-95,6357,-5087,1243,-1619,-5405,2922,-4653,-3229,-3220,7734,-3020,1101,902,5937,3906,8461,5454,1088,-285,1107,9726,-4746,7514,12324,2087,3239,2344,-11220,-3640,-4648,-3347,-3081,870,6025,2318,2531,-1179,1473,2081,1776,-1034,-1654,5634,-116,259,2193,4267,-390,-5917,-4565,-207,2529,-2496,171,-3137,-1282,-2893,276,-1708,-1356,-1566,3278,2238,-1890,2932,2912,13623,-1008,1571,1143,4084,-2897,700,1455,-245,-4340,2504,-5615,-1632,5678,5229,1663,3422,-11,352,783,3110,809,2193,3000,-6015,12490,2200,-5595,1169,4660,-269,3725,638,-3120,1185,127,1519,-2194,371,-473,-107,-1036,1452,4123,2355,5678,-2929,-6528,3420,-2988,-1435,4411,3481,2810,-4611,-1964,-2839,-217,-526,-1396,-6313,3666,-1905,-1966,5205,-629,4143,-4628,-384,-326,2866,3996,827,-2907,-1705,4099,-1900,-85,3120,-3007,791,-5874,-4416,-246,-1850,4694,3618,2392,-2927,163,-1045,-3498,-3439,4504,2792,3457,432,-1372,1015,509,-2534,2119,-1789,-3806,-4213,6967,-185,1243,4226,6264,-391,3237,2384,1629,-339,-3801,-3576,-1269,7148,2054,-1111,-957,5375,9335,-5776,-1561,2673,-452,-1356,191,-1953,5273,-3400,-5458,-9116,5449,-303,-6323,-8808,-2103,-4726,-2429,-6635,-1296,-1213,-78,-2089,-10156,-937,2519,-1785,6210,7753,-2800,-1646,4680,-3210,2249,-550,-4150,3947,-1578,-5302,-3251,3100,479};
    Wh[3]='{-2863,4489,-1463,-1452,2243,1173,2413,2163,-5385,585,-919,1712,1478,3156,614,726,-1215,-935,3339,2264,729,371,-1062,-5429,-1192,-2210,-1134,1176,1079,-1776,2149,-4062,-5375,-960,3774,906,7285,-60,-3061,6054,249,3125,-3203,-3789,714,2492,2156,-20,-1174,-3066,-3591,4257,50,-2008,808,-3415,-315,-5488,2324,-274,-1921,-4309,1931,-1641,-10,-528,90,3686,2595,540,-1083,1810,1856,-6093,-3955,6025,-6010,2143,-466,1474,550,1217,-933,-3486,-3525,-5312,819,-2224,-6933,-197,-1782,-2641,1264,-1551,5200,2415,-3188,4074,3745,2489,1101,496,719,-7426,3837,-463,-1477,-2475,-3630,179,2526,-1182,-1809,172,660,-295,-657,6230,4934,-2697,-87,4833,-6894,-2060,-562,704,618,5585,501,-451,3208,-4138,302,2863,-6347,-4045,-1861,-2462,149,964,-5493,3374,4187,3950,-477,-3159,1309,-6967,4868,-4953,-306,1200,1843,-5444,-971,-2641,6064,4025,-1298,-3237,3327,-1413,-339,-9423,2753,1872,-755,2044,172,610,-1857,5766,4919,-5522,-1585,-3518,-5156,172,555,-3305,2602,-1820,3642,43,-6313,-4392,3908,-2685,-403,-494,1013,-5610,202,7231,1990,1262,2629,3227,-692,5864,2912,437,-3784,-5073,-315,1662,1982,997,1625,431,1120,-2509,1551,-2126,5263,1296,1029,11982,-913,-3388,2917,-3181,-3574,7709,-2893,-3725,3483,2473,-4133,4321,4243,2758,-455,3916,-2805,2768,-1027,-449,1864,393,-2409,-447,-985,-4550,-650,1583,3879,2415,-3891,2717,1172,2093,899,3137,-528,3601,511,-3750,-1177,-416,-2436,389,-753,-5937,1018,-1385,4658,39,-1734,-1122,2858,3796,-4626,5937,-4018,-1396,4594,-925,1752,-1870,-1494,-2841,-5991,2646,-1195,-777,-2780,-3586,6269,2022,2607,-102,-408,1806,1491,-558,5937,1042,3940,1462,1879,-4226,-3320,-4157,-1894,3161,814,3503,-4321,-1168,-3901,-2961,960,-3183,799,4343,-4645,2690,-1110,1885,2604,-2700,-2536,-3977,-7285,-2147,-805,1851,-2878,1910,-2583,-1851,1205,-1995,680,-2746,-1552,6040,-167,-1,-1101,2380,684,565,1539,3723,1718,3203,3779,-944,859,4316,-150,-2897,2435,913,-3552,-6660,2122,41,2065,-5805,451,-3188,981,-2108,2756,631,4787,-2731,-1066,1779,2878,2956,1614,-255,-2663,-628,1490,-618,-530,-1520,-3569,-6357,1520,-5585,2156,-469,-3886,-4216,5185,-2329,-5190,6298,1268,-1325,6601,2758,-2780,-509};
    Wh[4]='{-845,2348,-3120,-3098,-796,-265,1809,1276,32,-2117,-1944,1028,-1264,2109,-5312,-2032,-6132,-3283,-1325,410,1817,-1213,2203,989,-1770,299,1112,1821,158,-2263,-436,2177,-92,1652,3085,-1467,3349,-1282,2871,-1693,-2437,-2597,2199,-2751,1372,-2673,-2274,-1606,-2475,-202,1110,-2188,3227,2761,-152,-7446,80,-1469,2321,-3012,1362,-428,1070,-3327,-2990,508,2253,-1264,-301,-873,1805,-587,-148,1467,-1380,-2186,-1351,-33,2521,-277,-2264,4233,-1239,-1861,-1063,-1347,-1108,486,668,-1835,-2480,-5263,-1512,-2646,-931,-402,-503,270,1330,-1054,-2062,-853,-1899,5249,-1600,-1047,-91,25,-1984,2590,-564,-6337,-6459,1206,-3039,-2495,181,-693,-21,3161,169,-2878,-3220,-6440,881,2049,422,-1213,2418,5244,-4941,-2156,-390,-3598,957,1026,-1781,2006,-859,3071,4938,-2700,4851,1289,986,4711,1951,2437,-306,-1984,653,5556,197,472,-84,8959,-2534,-2731,-680,-3420,-3234,2368,1732,-3254,1086,-722,-560,-5024,-2161,-1401,-3186,-6718,845,2420,2347,564,-2209,3054,-1064,-873,2092,-1391,-3378,521,513,1663,1719,-569,-207,522,761,-3579,3420,4169,-1833,-5034,1523,-2094,3161,-2221,1920,5708,-25,5146,-1652,2851,856,1518,-3020,709,-2235,1893,-842,83,2868,-6245,-985,-1685,206,2043,-1682,-6030,-2122,-1823,-3481,-502,-4006,1047,2393,3225,-115,8789,-350,1033,-4069,2561,-897,2133,79,6118,-3698,3410,933,4748,-874,2027,-2556,544,-2237,487,1545,142,-191,-3081,-969,422,2004,-314,-168,-834,-533,-2213,-1940,1071,1452,-2121,-750,-1348,-1232,50,727,2578,-443,-1979,-128,-2027,676,593,-3493,-578,-1726,-221,-3186,4475,-1446,147,1227,126,-1480,-1556,-3657,-611,1278,-1196,-1282,2144,-1068,-5048,-2423,-1052,351,-65,161,3024,-578,-2519,-4182,3669,-567,-604,-1417,-1120,-4382,-2379,-1093,-783,-15,-1790,-2685,-1582,-4272,-6181,-962,2954,-1596,2022,-1578,280,-1006,1278,-4499,-823,4365,1953,-680,-1997,1378,-2941,665,-163,-3940,-1064,-223,1146,3068,2980,1453,-4685,-2188,1284,-2702,541,1656,-2556,379,-1463,-2231,-2186,-2377,-3161,-943,-2266,3811,356,2504,-5571,-2409,6459,-4858,-8115,2155,1982,-4650,-2307,-2160,-1146,-1757,-1091,1441,1867,-937,-34,-2836,1843,-2592,-2371,1280,272,-2437,-4091,-1890,1322,-1446,3029,1613,-333,1865,3823,-3237,-3271};
    Wh[5]='{-1496,6523,3295,-1099,-497,-552,-7524,-4521,-1317,671,-3007,-98,-4887,-3542,2086,-1333,1965,-511,-1333,-1536,629,79,-1770,-2854,-1033,-1541,-1412,-1400,-2486,1240,-1680,-5732,2287,1066,-506,762,517,2135,-2117,4611,-34,-426,-2205,-2685,-6367,458,-5869,-1269,2819,-2500,-2409,5122,-483,-1711,-3364,-3833,2312,-2189,2995,722,-2968,424,-3098,3181,585,-1759,-1159,-2661,-747,-2595,-3784,-2235,2807,-792,3723,-3471,-1575,-3789,-2238,547,2270,1563,-5175,6484,328,613,1616,3581,-1192,-3466,-7,-133,-322,-356,-5781,-2141,-530,3273,-2049,2570,-833,-557,363,-7373,-897,1776,-3041,-3908,-4865,2423,1387,384,-236,-1203,5014,3835,733,-2260,751,-122,-1301,-5302,6049,9233,-1252,-4294,2224,1323,-4956,-14326,3034,1016,436,-3383,-3212,1824,-1143,-396,2421,-968,1563,2612,3369,-1801,-225,2252,-5747,-5590,-3220,-3137,-5380,-6191,-3713,3627,231,-1185,-1701,2531,2213,8129,411,-5546,-1335,5268,-414,-1440,2207,2807,367,-3903,2279,13906,-361,4653,2880,-185,5639,-2744,1417,1033,-3378,-8159,499,-2215,-2988,3957,-1358,4829,7768,-346,2022,658,8613,-931,-3198,-9189,879,2103,-4885,-3247,-1286,-2067,-885,-1895,-4763,-258,-995,1149,3598,2121,3286,906,3752,5087,-1171,2661,-3085,294,2374,-6357,983,-411,2124,3198,1174,1928,3161,-3947,440,329,3051,-877,1337,2371,1975,643,3913,1394,9033,-480,4755,-7548,550,878,2648,991,3010,-300,1353,3225,6123,1262,-3400,1334,2517,-4531,892,592,38,50,2502,486,3464,1341,1708,-419,-877,2247,-736,1276,5571,-2780,4760,590,1748,-1916,4560,-2403,2575,1538,3901,-1569,-1845,1398,-2203,-796,-1944,697,770,3752,-369,7548,-199,-3679,559,2038,1604,-4272,6621,-2442,-1770,-366,1364,5102,-293,2783,1007,-4870,-567,2900,587,46,-1467,6640,1479,-6528,-2985,1148,3239,-2399,4797,1937,2797,-1700,-2059,1129,4582,-1779,-1627,-223,5068,1835,-361,713,-3828,5869,-1240,4448,-278,1262,5922,-4775,-808,-1004,-2147,-755,-6259,3864,9843,-1995,-4201,1453,2795,582,1201,-6372,3891,11113,3544,-2875,-3027,664,2227,4997,-2578,1035,-1115,-6596,-1480,2092,-1391,-3305,4985,3098,3320,-3154,-812,-1943,-592,671,-664,-1098,-4482,-1182,2271,916,-1605,360,2318,2454,-8388,-6059,4174,-6289,144,-481,-10595,-4045,1076,181};
    Wh[6]='{-2973,526,1638,1927,-1418,-1130,-357,-3164,511,-684,-1735,-3750,-610,-4489,-1026,-7114,657,9306,694,704,-1702,-433,2352,-2407,-1657,1783,5292,-159,643,6015,3244,6699,-6552,-1015,-9833,883,-7226,-3088,-4406,4794,-2744,-1961,1739,1693,-2985,-1250,3083,-2227,-2512,1108,-2573,1838,8715,366,5317,-5297,2464,-4855,-1472,-2622,-1916,2919,-1750,-2568,-1666,783,1088,1409,1278,2937,-3869,-320,4233,1367,-6904,993,822,1363,-7246,1126,-1406,-7500,-1363,10283,322,-3608,-558,3022,10,-5708,-1883,-1676,8232,3813,5092,-428,1054,2998,4438,-1947,-2341,2093,1610,15673,3349,828,2360,13623,2335,7294,4111,-6000,12080,-3637,-581,-5249,-2695,4973,2851,886,-3078,-11044,751,3146,3984,-2534,3071,6289,2844,-6665,269,467,-1798,-4865,-6049,5712,-2106,-7255,-2396,-1308,-429,9399,6215,-2351,-1004,-2493,-2131,-1787,1043,-1245,2399,-2495,2265,3715,-1148,-3249,-10507,2968,2365,-3266,-1622,3967,-4533,401,-1711,-3376,2915,-502,576,1019,-8828,-1192,353,3510,-11103,1051,-358,-2958,718,-2990,2937,-820,17031,2673,1748,2788,4213,4753,1604,-3264,4724,-1973,-789,-3605,3647,1557,-5332,-4892,9238,-3969,-1579,-1239,1425,2988,-1210,-220,55,5869,4689,-4047,1105,8378,1535,-516,-1845,7304,3847,-1804,1564,-1728,-2487,8950,8662,-3125,-426,3642,4836,-1107,-5366,-1650,-2137,2053,1602,214,6479,2358,1851,2014,8989,-3674,448,-4509,2651,4094,5947,-4138,-3342,-2949,10498,1827,2854,-2846,-1004,-1564,361,5498,2788,-4262,-3002,-3200,-3115,5009,-4240,7714,6284,1292,-3815,2017,-1571,-3098,724,2995,-100,-2849,-3808,-1231,5903,2561,-24,4423,4006,316,-6054,-1428,4738,22,1425,49,-584,2082,-4855,-4912,480,4799,5107,7856,4182,-696,5439,1032,1363,-8930,767,-341,-1790,5947,6738,4826,-953,-4108,2565,-453,10791,1965,-10371,-3371,6098,-5478,3339,2198,1385,8798,2396,-433,-905,6958,9311,3400,4843,3605,-2054,2106,756,-3608,3010,13593,1700,-1156,-6757,3359,-1246,6274,960,3100,-6069,-385,-616,-967,-1741,2946,2365,3789,-1735,4638,952,-4729,4497,-12167,-14443,1034,445,2432,-777,-3872,-7309,196,4252,1616,-3144,989,3940,3525,5444,-8442,3168,-272,903,-2595,-466,445,3435,-1287,6049,3532,-443,-2966,736,-2148,782,-5273,-8681,4619,-588,574,2622,-720,739,-1091,5747,-49};
    Wh[7]='{-858,49,-1000,2321,-608,2902,-1904,7509,-1369,3471,6845,-1602,-5854,4899,-8461,-5800,3203,-1925,-4484,-147,-831,4541,-242,-2177,-1552,2222,-1190,1053,1226,-1650,-3840,6313,-1467,-3017,-4306,2556,-7397,-4199,-233,8774,-2390,-3874,-2580,3845,-6181,-9399,-5590,744,2946,-4814,6347,-1979,3220,-4460,-4804,-835,-1627,7695,-1036,3786,3527,2434,-1862,-5512,-8881,2462,-2673,5825,563,2073,1407,7143,-2565,-1152,-8969,-2143,8833,-1593,-1644,-2302,-1076,2260,-6860,2995,2269,1507,-3002,1545,1840,2283,-3291,-4777,-578,9125,4277,-617,-6879,-1574,5434,1397,3916,-1004,3535,3974,-2467,-1879,-6743,-4826,5737,-2454,5800,774,9658,-2944,-3361,-473,-3898,20488,3137,-4655,-1315,-7602,-4245,2568,6088,-8525,3491,2009,2258,3459,13535,-2749,1303,1199,-8847,-2352,-1835,-720,1145,-1712,11777,5942,12353,-9863,2758,-3913,-6352,-2431,-2661,1188,2814,2636,-3786,-1710,8920,-585,-17412,1365,2324,-8852,21425,4692,2680,6469,-1462,-12636,3295,2014,2695,-3520,1721,-1667,-572,-2410,-5107,-3674,-3481,-4274,2800,3117,2185,2271,2714,-1556,5844,192,777,8266,4992,-5434,7182,1022,1162,1534,1195,386,835,3181,479,-1579,3046,8208,-1738,13281,4572,640,2225,12177,5058,-366,2888,3537,8779,9184,4997,8251,-473,-8251,-1154,8173,1237,-2687,7207,862,3366,3269,1441,1926,-2039,6235,2763,7675,-972,4104,1639,-1127,6582,-2639,6293,-591,344,202,-2478,5185,4042,-1361,-2443,1575,2460,-631,-2095,-2539,1866,778,382,4460,-2445,1403,-674,2641,3627,2895,240,-1741,6538,1367,2016,1062,-2277,1802,2915,10312,-2758,3195,1297,6606,3908,1688,1932,-1483,6054,-702,-2320,-2259,-2744,1292,519,3220,-1855,2758,-910,-1933,6049,93,-2153,-2072,-3723,2412,-348,-1139,-521,-1397,-3715,1314,-2612,4414,2139,3088,1478,-3911,671,4802,11601,-5942,-5917,-1514,1738,1412,-3283,-2924,-1406,3483,4375,2695,-982,3615,-3520,3798,2790,2968,-2756,2493,6782,7470,587,4055,587,-2707,-1901,10263,-4028,2380,-1851,-631,-1826,1843,-5664,3496,7680,7514,-114,-2042,2790,4206,-4223,-6123,482,2990,-5312,3168,4455,358,-1918,1784,1727,4,170,4384,2302,3276,-31,6645,1183,-469,-7524,20,-3535,-1358,-3352,7080,4736,-1160,-292,3530,2080,-2722,-1006,6591,-2636,-4243,-1617,2479,-1433,3308,-2553,-4763,-6372,-3696,-429,5722};
    Wh[8]='{-1418,-455,-2354,-2661,-2048,2297,-7587,-2739,2299,2812,2232,-1697,-3894,984,-852,3415,36,1875,-921,-218,-32,1889,4614,2407,-1918,2873,-3898,-1702,-2221,706,159,1336,-1063,527,-247,-2312,610,-397,3364,2590,625,-2861,-2692,501,-3676,530,156,-507,-919,3837,-2235,-6567,-3615,-4089,-1954,-4472,87,-1148,2971,-1502,-2744,269,-1849,-3337,-6108,-6098,-333,-1183,4577,-550,121,2756,759,-4428,-1925,4079,-4262,1348,-2197,-1614,160,962,-2663,1140,-1130,270,1188,-5063,-5830,-2829,-1012,5449,-939,216,616,-3222,1431,-2261,2474,-1829,2932,-2939,1682,-1541,5454,24,-1652,-2457,125,939,2321,-3979,-2395,-2644,-1494,204,3449,3896,2028,-2358,408,2084,-1252,-2578,-8676,-7744,1861,3203,-1717,1800,-4206,2910,-2192,-2675,481,1744,3513,-1403,2008,331,3925,-1203,4433,-2509,-5341,2083,914,246,1494,-3125,-1047,2661,-984,6938,-6113,7968,924,4162,-7011,-2695,-4624,-1268,-4733,1124,3198,-1394,-1771,3620,1450,547,-6127,-1146,-2084,169,-1094,-611,259,2678,1413,110,623,-2471,2303,-1123,90,1193,63,-1290,2227,-3244,-6967,1133,2585,2420,-6625,6484,2076,-3337,2246,4836,-615,-718,-2178,1768,-317,1038,-1315,1227,96,-578,-4516,120,3935,197,-1660,-3134,-3330,466,-5009,-6040,-1893,3842,-4726,-1776,-1246,-4516,706,-3461,2111,1358,-1959,139,-4768,4631,-329,-1732,852,-1418,3469,-4785,-3215,2089,2678,-3024,-1181,418,850,-1765,-2198,597,-3830,-2785,193,-3063,-4062,-1401,-2320,-3193,1546,653,-2729,-7705,-3554,-5180,-2917,-5307,1185,389,-414,800,-5698,5273,-4355,-248,1657,-523,3601,-1218,2268,267,-4514,2205,-2197,189,-520,2797,349,808,-356,5,3056,6020,691,3171,1207,-1745,2091,-3730,-4875,2685,-293,-3432,-2541,231,-2197,694,-4541,-1865,-427,-6689,6928,-1730,-3842,-4125,418,803,-708,2194,-4245,-5581,-1138,-3261,-967,640,-1174,-1397,-1428,-3330,-6630,1708,-1613,3342,4440,-1669,7485,186,-267,-3803,2187,3283,-3598,2116,2133,-1743,-2391,4716,3654,327,5170,200,3264,-1102,5102,968,2744,1723,-105,-6469,-3327,-3310,-4907,-1917,1789,-3342,-4362,3916,-3107,4060,-1208,701,-5590,5278,-5932,-4992,-5175,-228,-562,-2242,-2641,-2115,-5327,-4841,-4885,-2169,-117,-2457,2244,-913,-6542,655,-740,2241,-6010,-2727,-2687,-2233,-323,-2248,-1750,1829};
    Wh[9]='{-3085,4235,1091,-458,3920,-1107,249,-1989,3657,-1075,4736,216,710,2006,6938,1749,4296,3842,-834,-308,1551,864,-2213,2208,873,-1679,997,-379,3415,3054,1896,1511,2335,2174,1072,2631,-226,2447,1368,-3098,-68,-3161,-4321,3457,-2019,4218,3979,4753,-87,199,-761,-403,2612,3513,1284,5395,186,-108,1798,1026,-1724,4172,3925,-1024,1729,-1144,-1192,6826,1873,-2294,1861,1561,1015,705,2469,4033,3569,2749,-3059,-1238,-105,5966,-764,1397,-3725,888,524,3510,5937,-1826,-387,4733,3825,842,-1220,-447,3464,-1064,3432,5551,1110,-2346,-193,1661,4694,198,5449,3193,-5454,1342,273,-2885,2241,5351,1253,-370,4218,-5917,3469,1340,-1677,991,-3796,4204,-1062,-439,3093,290,-4855,-6367,4028,430,2416,2115,2054,-1190,-3666,2648,-396,-2629,-7495,-3781,640,-2851,-4846,3745,-2575,1594,2770,-1014,-4382,-665,-1280,296,-3112,-3940,469,627,-1510,5175,-670,3117,229,1192,4057,2778,4089,-4,-741,-1155,8203,5966,-2279,-2788,-3620,-1518,1267,137,4912,742,-463,1906,6391,-3596,-39,-2052,-339,-393,-7827,-2456,789,-560,413,3198,4357,91,1289,880,-1362,-3823,2342,-328,-3757,3127,1745,-772,-796,401,5771,4743,20,-1733,-6171,-4067,-4313,-3605,-1267,3176,-63,-659,-189,4675,1844,-233,81,1759,4599,-381,-2734,4140,828,786,4182,-336,5585,1223,3872,725,-1185,940,-1295,-6435,158,-508,-1398,-4663,-1495,-1684,-1997,4816,-1141,-968,1212,-2861,1938,2293,-5278,-3312,-925,-3894,-885,758,-5000,3332,-774,-1723,-1632,-5063,877,-2722,1712,-3110,4130,-4880,-722,-3476,-812,3410,1213,2917,1992,2893,-2839,-5107,-14,2019,-1273,-1041,-3383,-1407,7973,834,-235,56,-892,-1386,1062,-286,-58,2963,210,1228,-4672,406,451,5820,4392,-3632,1942,1082,2202,-2056,-1072,5664,-3034,-249,4609,1605,1545,910,7734,3503,956,-1256,3701,-721,2614,334,-2330,1397,6298,-2897,-4562,905,-3574,4111,2008,6684,3371,-5004,296,-1167,-491,620,-1914,3891,944,1993,10000,-1166,275,794,147,2587,3337,-5771,2788,1948,-2561,4775,-1273,2296,-346,11,1296,-4833,-2597,-5991,-1215,1889,917,-2451,6245,1204,5478,-162,-2215,127,1900,2003,5600,-1983,-1256,-3122,-1643,2142,495,564,-1824,2298,3161,-2000,914,3039,-1900,3974,7998,839,908,4624};
    Wh[10]='{-725,6064,1993,2310,1364,3750,-2352,3896,-299,-1916,-2211,2294,7377,-128,-1846,4465,3981,-236,2770,-3522,739,-4216,-5429,-1472,-181,-1613,-1315,-392,1546,3012,1533,-707,3205,1074,5693,463,-3845,829,-1055,7250,1285,-3427,-2490,4729,-2775,1599,3835,-493,-3166,30,-462,1308,-1807,-734,-5898,6904,3376,2985,-914,-2958,-1915,311,4594,-143,-2218,-3374,558,7236,5175,-3911,3803,6210,-831,105,-214,558,4704,8232,58,-3395,-972,10166,-906,-3208,-2539,4494,-1040,87,-3901,1123,5742,-2242,10937,-2666,7944,888,-3193,1903,3459,-2108,-855,4438,1207,8505,-382,1335,-1678,-6230,5366,-1188,5869,5029,4548,1568,4707,1011,-1480,6801,-2493,-12724,172,384,-4777,7500,3071,-8740,11591,-4082,-8793,-1104,-3854,-2246,-6064,5141,-2734,-2072,-3212,679,-5942,-2132,3945,2226,-4455,4733,-1513,706,4143,-2902,-1416,-2849,-448,3559,-4829,-2873,-686,620,-9726,2692,2502,-162,-13935,4353,1569,-7685,8120,6723,3273,3188,468,-1958,-2435,203,-1762,4401,1439,-6972,5854,-2072,3603,-3811,-1585,-10117,6933,491,-634,2131,1317,3681,-1539,5805,-10214,-4868,-864,4453,2204,1790,2220,-3579,7460,1613,-1021,1993,-2078,-7070,-1307,432,-1124,1035,7739,-2719,-3076,-456,-8784,2536,3720,-2095,2690,8388,-2834,-1832,-1223,354,-1522,-91,-2817,-11220,2915,-187,-4057,-4819,-4914,7856,-3486,-1235,554,-1265,-2751,2301,3737,447,-1064,2658,-1413,8867,2988,-919,-1263,-1026,-3967,-4599,-4370,539,-1801,-94,-5048,-5732,-4323,-1795,-282,-1767,2946,477,3840,-903,2644,-7397,44,-130,1823,-2470,1610,2016,346,-2294,-844,2340,5263,-6582,-785,2468,10849,-1717,-1986,-2629,37,6997,-1542,5224,3886,-116,10615,3535,-4584,2919,2080,-2279,570,-1715,2127,-1877,1132,2807,6879,1243,1928,12080,1833,4257,-1481,-2770,-811,5405,-1041,-3889,-2944,516,4816,1494,7368,-625,-304,-2236,3911,-1896,-1746,1630,2790,3493,5844,3005,-171,-147,3103,-1533,-980,-1867,-621,-94,5971,-3066,363,-279,2412,2915,3908,-2015,2438,-891,-3378,1121,6015,78,3310,-6005,-3369,3374,853,812,1185,-58,-3085,-3879,4670,-2148,6347,-7006,3439,6367,862,-3784,4184,7846,4047,-3312,5351,-159,1395,331,5908,236,4230,-1583,507,291,-2702,3530,-1915,7563,924,-3005,6748,-3876,4931,2883,2800,5180,1701,827,-5043,-5112};
    Wh[11]='{1755,3503,730,511,-2644,-1209,880,617,3742,1267,-1257,-1746,-1163,3225,-856,2250,3120,1384,-3686,-1940,-705,-502,429,-437,-1583,-35,614,-27,-297,-544,-2493,-122,3125,-569,-11,-2509,-2470,-2827,-1436,-597,6035,1373,-942,2009,-3688,-1165,-1093,266,-5288,-591,-177,3068,-3298,-3044,3754,-225,2788,-4020,-302,-247,-734,-75,-128,-167,6015,-2362,2976,-560,-2893,3149,-1944,-117,2687,1679,-1424,-2231,-152,-1820,1545,-3933,455,2563,820,2685,-797,2026,-1345,-1160,4509,-319,-4436,-1220,-196,-1268,769,-1069,182,-2741,-2257,1428,-2004,2171,1933,1510,3564,2482,2563,3747,6181,-3437,2247,-7978,4697,1604,-339,1572,-5390,-1044,-5185,-5146,-501,1796,-1368,-1683,742,-3239,-2374,2358,-410,-1953,-7988,-517,3215,-1468,-3071,-2274,-933,518,-1553,-1774,-1210,321,1956,2484,-3598,-4758,-4843,-252,-1956,748,-608,-1867,299,-6298,1970,5361,-2194,-2298,-464,4426,2062,2548,4118,883,-480,4846,4475,4514,2807,-1580,823,-331,558,-540,-1254,361,-3627,1276,1850,-434,-1740,4941,3159,-2966,6669,-2132,-3610,-6108,1790,2770,-5053,1370,-6660,-1224,-1600,-961,-913,2863,1474,-1478,-862,-616,1558,344,1092,-656,1904,-429,-640,3793,-4331,1546,-2164,-3930,995,-9501,-2348,-2438,-4201,-4758,-419,-3142,1312,-4274,-36,1126,132,-624,-3232,-44,3579,-1343,1331,-5717,-5449,-317,2729,545,-4543,48,1422,-2022,963,-1495,-2707,1549,-1220,594,-2871,-3486,1082,-1811,814,4248,4597,-710,-974,569,2420,-4125,3120,1948,-2468,-3034,-308,-2473,-222,2070,-1486,2080,-53,513,993,844,912,2150,-6333,-2727,1174,3168,8198,5585,2683,1995,-485,-793,-3742,2683,13,-1778,-1049,2556,1186,-736,-638,-238,-147,-5498,169,-1582,1560,1812,979,2690,-98,1632,76,820,-4921,2731,-94,971,-1978,1385,-1184,2380,-949,-1159,2491,4768,2331,4335,3117,938,-4367,-799,3786,823,-3491,2985,71,-76,1481,-2036,-4577,-1418,-4121,656,825,-7,3095,-4936,-455,-3298,-2137,-2739,-3671,-2980,7382,-1192,-2154,173,-957,-2436,1545,-3728,-2873,2231,-809,-48,3823,1728,-78,-837,1569,-2387,3457,4345,-217,484,-5581,-3120,-606,-4064,-852,-1448,2595,-3669,-4938,4311,5468,3698,1756,257,-3918,-4306,-4809,843,775,5356,-4882,-124,292,-1060,1258,-1601,3256,-313,-3723,-4531};
    Wh[12]='{4030,-146,189,2648,929,-1872,-4299,3754,4252,2736,-444,-1186,-3483,-88,-3034,853,-1051,8750,-4589,-3713,870,1102,-3000,2148,4985,-3779,-331,-1032,-14716,791,2797,-7294,3488,980,-3759,-2203,-597,-2336,-1284,3791,3188,3439,3764,2012,-9365,629,-928,203,-1458,3151,-6904,-745,-1650,2807,652,4729,2912,546,1452,5610,3603,1257,3405,-17,1688,-3347,3378,-605,-2435,-814,-8759,-9975,-3579,6293,2105,5205,-690,-384,-3366,1258,-871,-1500,6225,371,3837,1065,2220,-2697,-2023,-4221,822,-1352,7788,921,-2437,-1177,5781,2954,-6093,452,-2880,-814,1816,-8056,-1442,2824,-3220,4750,4829,-5771,3879,11943,-1008,-674,1264,3085,-840,2370,-741,-2646,-2116,2932,-8369,-2949,2629,4511,-3439,-1721,-311,1824,-12343,4208,1878,-373,-112,1707,5039,582,5380,-6362,-396,-3312,-92,488,-2990,372,-4238,-7055,-468,332,-3518,-729,-2678,4372,-4125,2861,-5864,-819,1982,-2521,10537,-2075,-3449,5927,-2500,2127,-1752,2917,643,-1101,4125,3041,10605,-132,-3410,-4768,-874,1503,4558,1105,-4035,-622,4113,-2963,6220,-3022,-3010,-826,-5327,656,-1640,1373,-3735,-913,2376,-1594,-880,1146,220,1014,7,-6489,-2,-38,1168,-1489,-5683,27,-1655,-1871,3046,-1546,887,2314,-2800,-2344,-3984,1235,-4179,-1446,1027,-3088,-8354,3039,3613,3459,-2868,-4479,4572,3847,-3642,-2631,-13857,-494,998,4575,-4787,-5664,524,1002,-245,1787,-459,-419,-509,427,3308,-1623,-7324,-2105,70,2580,11,341,-1165,-1101,-2333,6113,1539,-6347,-2133,6118,4763,-2235,-921,-771,1799,-3288,-142,297,3269,-3967,4509,-2368,3918,-180,5117,-3134,-2536,-2056,6767,-6542,-5483,3327,161,844,547,-12763,2481,499,223,1021,-3457,5043,-1962,-8559,-767,-105,1467,1029,-850,26,6005,3950,56,-1436,-6806,-507,1883,-1832,4433,-5126,-247,624,-3549,7548,-3283,5966,-2127,-2473,7299,-2529,-510,321,3808,1667,-2421,-1209,-4235,-115,628,-4252,3996,5361,-3854,1997,-4663,-3630,4804,709,-2319,-4672,6318,1182,925,1278,-5810,-535,-2250,3676,-4323,744,5014,5732,-3483,-413,-298,278,4648,156,-2498,2644,4204,-817,-5029,5468,5659,-2352,1127,2900,-742,-5117,810,3576,-546,-1407,-2836,5097,-2834,-3945,4975,-6093,-3107,-1766,4514,-2406,2312,-8496,-7075,5883,4223,451,6049,698,-4382,-7646,4011,-1723,-6547,-137};
    Wh[13]='{1318,-2736,2849,3657,798,1824,1989,-4602,-1994,978,-247,-5498,1223,1021,-3222,-7114,4125,1633,-1746,2127,129,5488,-2197,1645,-884,-2239,-3540,-502,-2414,1193,-853,4821,5092,583,1475,1105,-1662,-6459,-2354,6025,6430,6562,-3720,1341,2088,5966,-7036,4489,-288,-1296,3356,1312,3083,-3356,-4018,2266,2822,2519,3388,1905,-372,-6064,1436,-2749,-2995,3859,619,1166,5415,-4335,219,3046,-7036,-989,-28,-949,8540,-811,-3098,4228,67,-65,-3984,8496,231,-1345,-1629,1166,-2907,1046,1807,4196,-1756,-3264,2666,2014,-2183,-499,4116,2224,-7163,2213,422,-7285,1231,1849,-1857,600,5444,-4624,-4709,-2827,2561,1593,2193,-239,3708,5800,2384,145,2507,3398,-2668,8330,5371,-12255,10439,86,-6557,-2351,2502,-569,-71,13,611,-1937,1253,-7373,-2014,1147,-390,779,-3793,-7495,3105,-3864,120,-5195,1944,-199,412,-1334,8032,-59,4147,-1,5898,2460,2111,-6020,525,3183,-3024,-7202,5092,-2770,-3601,-765,-614,1469,-3894,6176,-8515,4692,1324,-867,-3493,-4641,-2622,2309,5961,-3933,-5908,-5249,-1008,563,-217,2980,-5771,-256,-3574,-3723,-7031,-2641,-1616,2099,8012,-4423,6513,-1706,1101,1416,-1083,-10097,-3220,-1420,-4155,1971,5156,2983,-2724,1291,1236,1785,-660,-294,3642,242,-1186,-906,-288,8432,3405,1448,1199,-4255,-4069,-411,1202,-2340,-577,1956,-2161,1954,1446,-2897,5693,855,2976,4536,-5151,800,1583,-994,2386,-445,4973,-3898,-1550,-3000,-3093,560,-2810,1024,444,-160,-3344,-661,2019,1237,4187,-2565,1165,-1955,-726,2419,-1425,1144,870,-30,-3225,1739,1898,-1027,1545,-956,-2458,-2347,-4592,-3298,-7226,1947,-410,-2829,-863,-1617,32,-7,-643,2019,-726,-5043,-964,1362,-809,-4772,1330,-5541,-2381,-3029,185,-2426,-4313,-647,-1618,690,2832,-7470,-4020,1883,203,-8193,-983,-7109,-2536,7651,6596,-3264,-4545,1257,-881,10380,3315,998,507,-1812,-1036,844,5312,232,-2078,-806,-1026,701,-5747,5922,2695,-3557,1928,-2968,3430,583,613,3425,2746,2045,262,1643,480,-2548,4821,207,701,1423,3217,-443,1473,2188,-194,-1021,1734,-6875,-1651,1704,6787,5317,8857,-2534,1958,1859,1178,2519,-3896,-7553,-2517,-6665,5957,-4887,988,-1685,-2474,1667,-4841,1883,69,1318,-8032,2110,-5410,4570,2958,581,592,-1066,-572,-160,-3857,31,3659,789};
    Wh[14]='{2225,-6958,-1249,2617,1492,2277,-519,2041,-2614,2968,-5209,89,5507,2071,5053,-8706,4592,2008,4799,5366,1312,2717,3493,48,2844,4707,3918,-520,3041,3188,-1232,3076,-476,-80,-4572,-750,-3911,1906,890,-4062,7861,-19,596,4714,2546,6064,8183,-2473,-4208,-1194,-1162,626,-2056,1340,1066,-4694,1888,2404,-2396,1017,-1610,3847,3222,2504,2656,891,-2924,1017,3005,4291,-619,-1855,2851,8291,776,5776,-2368,1274,-3085,617,-950,4853,-1936,6103,2675,166,-4311,638,3129,-1093,-1289,3937,700,-1572,1054,70,3720,-743,2261,4536,-1600,334,2399,-25,5483,-76,3173,8774,1676,2529,3125,910,-14199,-4072,-1970,-717,1628,-1392,3686,7998,-294,-835,-6508,-2261,-2905,4042,-3225,1628,786,6123,2565,-3850,384,914,502,4101,1414,-4284,679,-2541,1569,686,-292,3742,-3933,-3107,2017,-2846,737,-3962,-285,592,130,-982,812,-6811,5751,-1445,-3676,-11269,684,-4995,-4216,-6005,272,2597,2141,-3835,2895,-2546,-1110,527,7978,-3676,-1427,-98,-3747,-1549,3425,-1213,-699,2548,3581,-5253,-1949,-2176,-192,1453,3417,-1530,-1137,-791,-3088,-1928,-3491,1445,-2277,877,7729,4030,-584,676,-1446,-1022,-2517,52,-1313,4565,1097,-2749,-215,1054,851,-918,1467,-3493,-408,-6982,1365,-856,-2534,1713,3344,-4616,-3395,9082,-3132,-1855,-4016,2509,-653,-83,5996,3215,-642,8959,1491,-1474,-2448,5590,-5434,-3332,-1604,-1676,1324,3447,-2993,-1150,1311,-839,-1452,-851,-6118,-3054,-4897,445,-4423,-8715,1448,-61,3352,-2073,-1348,-876,2873,-911,-7431,-1008,269,-1107,1137,3991,-1097,-125,-6538,7573,-6499,-1733,-4338,-1218,-3088,-1770,-980,1971,-926,262,-700,3825,-220,-1029,4604,-5869,4377,5688,4067,5092,-987,-1805,3215,2790,-414,-2031,-5708,4831,-4313,4196,2834,2500,-1192,-5581,-95,1280,-1322,-4240,3784,-2624,9204,1401,2351,50,-2229,-1247,-2069,4421,1585,1536,6621,-97,6591,4091,588,2209,2402,-2347,-1035,-405,2250,4348,-795,2191,-1348,5166,-2175,-6547,-2163,-1152,5742,-7592,9238,-846,1193,998,-2556,-6064,-996,3146,-1422,-1171,-6269,849,7109,753,-2512,-1048,-5429,-90,86,3413,-3649,6782,-2213,-989,7045,-6186,8154,684,1181,-1573,151,-1816,-5219,5092,9560,-3161,-5307,1793,2722,1226,688,4892,4733,-2519,-3417,4467,-451,5380,3752,1165,6635,1414};
    Wh[15]='{4309,3547,-3256,-3666,832,548,-4868,-1104,2303,4172,547,-2004,700,-4577,672,-9145,-657,4169,761,1593,781,599,-2052,1594,5830,809,1374,2797,4655,139,-3325,6259,3708,-1407,-5126,3840,-3618,-1646,1213,6933,3872,3569,7973,-3056,5556,262,-11201,-2125,-6293,383,2426,-503,-6645,5927,5742,-599,-3332,6362,-6572,9335,-5502,3679,-3381,12070,4958,1593,-1817,-3615,-4477,-630,-3298,-484,-2275,252,2218,-1029,477,75,-1712,469,-330,-659,-2502,5136,-6186,475,-458,1898,-2695,2600,1572,5981,-3496,-3171,-6000,136,-5366,9594,-4504,9121,-8408,2156,1729,-10380,-8291,-2110,-3747,-1064,5732,-5336,599,1300,5815,-2105,2546,-6772,2336,1704,2661,84,-1591,-2717,5791,-2905,5463,3127,-5395,-7006,3103,-2885,7631,-2631,3991,3776,13818,3010,11220,1735,1099,769,4323,-4086,8012,-1100,-673,-378,6367,-8754,997,4562,168,-2890,-2641,-2416,-5468,12187,503,-5488,1654,21816,2368,2490,7802,3061,-2644,-1248,-564,1075,1794,-2272,-1452,-519,-2854,-4245,1927,4628,-1544,559,-3654,1340,1966,-1179,-4187,1209,1964,1690,-2086,-180,7734,3242,1706,2585,257,-3874,-6372,5361,3820,2135,-3410,-2426,2924,-4287,-3972,-2463,-2907,1472,-3671,-7231,5136,3332,-9326,-2379,10507,-878,-3674,-7045,-121,-3640,7163,2604,1679,1878,4616,3911,2824,-58,3002,1295,2634,-2346,9951,-2164,-2398,2203,-2266,-1608,4555,3337,-2961,-1591,878,674,-44,-3356,836,189,3269,-2495,578,-1954,-1997,2749,993,643,734,-6958,2309,5351,576,-7597,-4223,-2558,11816,-3676,-6372,-6479,2697,-611,1503,-328,-5727,-2602,4084,-2281,2374,6894,-4052,427,-2,-3017,5454,-4912,-173,9033,-765,-59,-1962,-10576,249,3063,5800,3725,-61,-2104,-2619,-5830,-9,543,-4287,4294,-2531,6835,-4133,3039,-5991,-5043,111,1704,-517,2027,-597,-3364,-1800,3798,-1740,-8330,-2347,284,6977,-3176,1925,1043,2624,-3100,3964,4592,-1112,-1813,-4196,366,2006,3591,1735,-1391,414,-402,-6679,-4106,6372,-1684,-2578,-1763,-3527,-2592,-1850,1022,2312,6674,-3461,-80,-3095,4641,-1335,2700,7670,11972,5830,-5585,2313,-5390,-6665,-5092,8437,3308,4350,4060,-8212,-464,3308,-7451,-1143,4567,-2060,-2814,-26,-1525,7089,-1284,-4199,-5380,834,14111,-5122,2714,-93,-707,-7270,-2946,-2083,-4846,-509,-3205,-1385,636,1910,-1177,-3220,-2446,-1134,1187};
    Wh[16]='{2117,1224,-2548,3327,1593,-1968,694,7031,1459,-1108,-1901,2066,3347,-3466,-3774,5478,2239,575,4030,1287,-6411,4602,-4707,1260,848,1904,6787,-3315,6533,-4519,5307,1702,-418,2077,706,1254,1607,34,-3735,4233,3149,4902,1800,2332,2032,-1690,3325,-3630,-1851,1920,1138,-5400,5527,1710,5419,-5649,73,-1270,2047,2739,-5151,3603,5131,-1822,3679,2770,-1248,-3598,3745,-4541,2966,219,756,184,-1165,6284,3232,1807,2507,-998,1395,6679,9819,-551,3544,-874,1883,5556,-1823,-641,4040,2541,3449,776,-1403,-1927,-544,2871,5585,1193,-5527,306,589,3330,793,4208,6738,1851,18750,-5283,3828,-9765,3557,1669,2071,791,4846,9770,-748,1614,167,16269,7324,7480,-7021,-546,211,1279,-4519,2829,103,726,-2597,4868,6845,8515,16728,-2215,2028,1094,8203,1560,-5771,240,169,2917,9101,-11718,346,-1854,6748,1458,653,3989,-4594,3918,8813,1048,-5659,2122,932,717,-204,735,1711,-5419,-312,4814,-5961,2178,-1833,-6337,-297,1724,3088,2978,455,-5283,-875,-3703,5615,3620,-2188,-4580,-5747,4970,-2717,4545,-692,-1396,-4956,-2144,5961,-6127,-4858,10224,4089,-5087,11357,1981,-3505,123,73,-8930,4414,-1185,-4282,-3212,977,2357,-9350,-240,2124,703,-428,-2307,1456,7963,-1628,-1130,-3212,-4702,712,-4150,3183,-4792,-5385,2404,-7861,661,-141,304,-3508,923,1593,-4548,-817,-927,1,58,956,1495,-4042,3640,2612,1152,-3388,392,-6113,-963,-5449,-4902,2269,2766,186,-341,-379,-3659,4235,-2338,-2622,-1065,2839,-5375,-9326,-5883,795,-1074,-917,-3544,865,428,-4462,-181,-5712,-3554,-3405,-11767,-2210,-4196,-928,2534,-1641,-321,-2612,-3623,-2941,-7177,-761,-2293,15937,-2744,-2408,-5717,2416,1351,-3654,-7758,-2080,-3471,-2998,-335,3063,-2924,2119,-1185,300,297,-2697,-3371,5253,-5029,-3007,-5571,-2177,1162,-2563,3947,-576,4528,5737,265,-3183,-8061,-2114,-1259,2995,5234,-1795,2795,-745,-769,-1573,-3679,4875,-2222,-91,2587,2041,-2966,3269,-981,-206,1508,-1138,-468,1209,1596,-793,3305,-433,3330,2498,-3852,6127,-248,1601,-5493,2403,4602,-2141,7,-1280,-3928,1505,4357,-3850,2324,2875,-8627,-896,-2932,2180,-6748,809,-212,7651,-231,-806,4287,949,6108,-2053,-3117,8173,-6713,-6225,2646,1223,4350,2070,195,3984,400,-5463,-4006,-3093,-154,4042,-5336};
    Wh[17]='{2614,1950,188,4067,76,2514,-6132,960,5883,2138,4638,5039,-2008,993,4313,-1335,3933,8251,2434,212,1370,2773,1927,856,867,1562,2363,-1771,739,-4343,-1693,-2983,-1418,-3269,2619,170,-214,1640,523,602,-631,-1494,3457,-3806,-355,-4052,-2727,4689,6171,2456,1584,2546,-3032,-6909,-2856,2673,1658,968,2092,-684,4350,-2670,-4702,-32,1130,3195,-1209,3635,1870,391,378,-856,947,1656,-1088,-218,-4140,-274,-33,-1311,-475,-870,-4855,-461,3154,2941,2512,68,-61,-3942,1933,-1732,533,-5283,-2066,429,-2858,673,-3542,2203,-7905,5097,1157,1593,-2934,-1464,-3642,2145,-1433,-9384,8632,2802,3486,-51,3864,-1993,7250,13554,-8437,-3281,1424,6533,11660,1938,2044,-13574,-475,-1124,-1329,4775,3146,3310,244,1828,-1074,5415,-2810,5859,1575,-422,6484,662,659,-3747,-4694,3232,10029,-3964,-2556,149,6630,2009,-922,149,3310,-1624,741,-2204,5170,7480,2425,-1290,-3493,5400,-1955,1213,-1169,3198,-1510,662,2247,5166,2236,98,1148,-1005,1705,-961,-6625,-3117,2751,-5883,273,1907,-7358,-336,-71,4870,-2749,-5600,260,-1650,-344,-646,-587,2910,4697,1630,4814,4099,4738,125,-2497,-1706,4421,376,1429,-295,6884,4143,4328,193,10000,5932,-601,-995,1325,740,5952,1145,240,-5117,-4184,235,-1014,-2380,1701,2302,2320,2368,1630,5717,-1726,4199,-1197,1806,-3557,-776,620,-125,1746,-3771,-457,1585,1801,4431,-4833,-1981,-4138,1954,-4060,-72,2127,4538,363,224,2020,1704,540,989,4089,1309,3825,-4738,640,1374,-153,2199,-2452,764,3574,-634,-374,-2951,-1375,-383,7705,-1124,2205,3708,807,1905,2517,-590,1579,-319,-1361,4428,-3312,-2347,4743,-5195,-2683,-5805,-5532,2467,-2866,-1525,-4108,-1130,6762,3605,-2180,6181,-260,527,70,2362,983,-5068,1091,2293,-3068,-3793,1373,6005,-1220,3881,7094,-3952,-1936,-41,-932,-2968,-1040,1398,659,6855,-4201,3496,499,-1927,1551,-1588,-5009,-4770,1772,4594,1737,3598,-1229,-2280,2507,1729,1323,-3063,-867,-425,-3583,-1127,-1550,3527,1524,858,3903,-4169,3342,-6923,1765,1148,7568,5126,343,-4418,3378,5800,-2668,2321,4116,708,492,-3869,2619,-1777,4616,344,1856,6967,2268,4748,4492,-8989,-1392,-4250,4130,-4919,137,1005,-1978,1639,2265,-2624,7978,-6591,249,-1867,-3449,4570,-1190,1394};
    Wh[18]='{183,-7089,-76,-3771,-880,-2636,-9,-1289,-4899,-223,4978,-1962,-4587,-617,-2553,-881,5410,-4694,-48,3103,-302,377,1414,-3710,-931,-2592,378,-723,-1231,-294,-1267,2480,-5561,2436,2622,1873,-1733,64,-1427,2724,-1589,1020,-1645,1409,576,-1281,-1284,599,5566,-4423,-1116,3066,-236,-538,-628,-1105,1929,-1834,-283,-3808,1226,-2072,2387,-1473,-2142,1435,-299,2851,-2707,-1617,-4877,4113,-2491,5747,572,-2263,-895,-3479,562,2298,-1398,1181,-5947,1317,141,-1047,-534,1851,-3288,-12,-775,-611,-1513,-1067,-471,1834,484,11054,4709,931,-2541,-2021,1738,1849,-6083,429,-237,2470,-6113,5434,-8154,5439,-2836,-2225,3652,-1527,-186,-4587,-2773,3081,-2126,2626,1600,3227,-5390,-822,4428,-2814,-2285,2597,1489,-2905,-3269,-1197,-5410,-2614,-5957,323,4052,3666,1856,-965,1348,-2666,-3996,3681,-3732,4245,-1216,-2717,2410,1923,-3430,2413,3579,-731,-6806,958,-4614,6728,-1901,528,2076,161,-2220,4572,12,1030,2263,-1059,2053,-4821,-6625,4809,-1370,-3913,-2861,-2556,-4685,-759,710,2824,6337,-1799,7133,1990,-2056,2849,-3100,3476,3471,2143,-4040,-4133,-1488,-8950,-4443,3125,-1374,264,1589,1514,1779,-293,-2519,-1251,2130,1021,7905,-284,1787,-4328,308,670,1658,5058,107,-2447,3566,2797,118,-469,-3845,367,-3027,681,-1591,-365,3210,7138,4079,3569,1644,-326,-8,-4326,1270,-1315,2089,-9760,5439,-3378,10126,-2202,96,550,-2846,316,5166,437,-3354,-174,432,-3996,2897,1784,1497,-1026,-2541,7050,2270,3193,1121,3356,5268,3603,348,-2668,1525,-517,2464,-3146,3115,-3894,542,-1155,-2670,-1124,2282,4990,-3029,-149,4768,62,-1893,3974,1853,2343,-3247,2152,-491,-550,-849,-2512,-2376,-1579,3857,-2058,-57,-1789,1663,-1610,214,-1490,-1943,7114,4343,2224,878,522,1278,-3933,1820,-3081,1184,1212,-920,121,2458,2260,-1579,5004,1064,1478,-786,1766,4279,744,-289,1903,2132,285,-7114,2653,46,2536,-4665,238,-7519,-2105,1340,-5224,6157,2524,-6748,-751,-2822,1683,-1403,-344,2753,1572,-3813,1986,820,-3464,-604,-1437,-2496,2858,-2432,-4216,2224,-3728,-461,784,5000,-3845,-1072,2700,3723,5053,-1583,-1064,941,-1712,-3186,-3466,388,599,-2248,156,1687,-2956,-146,-1021,2037,-1649,-711,3095,-6030,1953,-7377,4460,2150,2807,2105,1992,3117,761};
    Wh[19]='{-1257,-6694,81,5019,-1503,116,2597,-728,-83,-44,3078,3115,539,-4023,7460,-6928,-1152,4453,276,1459,-842,-2004,1170,-378,-4475,546,3784,2097,2741,3041,-2308,5102,-5458,-2524,-4304,-359,-6181,736,-411,735,-1859,-6235,-1115,1804,10527,-613,-1767,2391,3574,2268,2470,-3454,7612,1473,1488,-718,-1568,934,48,-1984,1203,4072,260,-697,-2336,7524,-1439,-1467,774,-575,609,3564,-2810,-2946,-2841,-783,-1960,-955,2910,1629,-414,-3718,-3872,1705,701,-3537,-3308,1214,-34,-2768,-3969,-4226,-1030,-2014,-8779,-41,-1571,-446,3728,-1818,-2336,1802,-4157,10195,1800,-1545,7714,10693,-291,-424,1500,-12275,-1555,3278,5317,3344,4594,7846,190,-47,-33,-3200,3557,1669,-2773,3415,-3442,-3498,7963,-17890,6206,-776,-3640,-606,4501,1413,-1976,-3515,1502,1165,2482,3493,8134,-2180,1635,-3483,3190,6030,2539,-3081,1673,4394,3491,1129,-4108,8183,-5937,-4340,3208,5371,6528,3784,-113,-699,-167,-6176,2382,-866,-3486,-895,-3117,-1295,-2344,2026,-875,2807,3269,-5034,-1156,1865,3881,-563,6757,9638,5786,5751,2218,10107,36,-5434,1226,-2100,586,-590,-2388,4973,-476,-4711,-5942,1226,2663,1490,3188,3305,650,327,1834,6245,-3657,-2927,-2163,2700,4038,-1257,580,5649,6684,-3942,65,-1534,1646,4184,5639,227,-127,1729,6508,-159,-1022,-2351,894,4807,3715,3234,2500,4045,1287,1937,8857,-6557,-2836,8090,5244,-3049,-2802,-1517,1864,789,4658,-2011,-618,182,2102,-1549,-281,-404,2337,-776,-2490,185,-2421,-4470,1890,4282,491,3020,-1547,-1319,1287,-1466,-7724,5263,-1315,-424,-1009,-2066,-609,1109,-253,1949,-2279,1679,2421,-210,3425,-2158,1247,1386,-4626,1234,-8129,-542,2622,-940,3283,1376,-219,1593,6855,-1519,-3847,-3867,-5048,-815,-644,-6323,6215,2083,5742,-1015,7749,-1364,1972,-1809,-232,-2098,1718,2227,1032,-159,-3076,5356,3515,-755,769,4328,8383,-2597,2617,591,-3911,6372,-1336,-1181,-827,7939,-154,-160,-682,2629,-4709,6899,-242,4863,-331,-5039,3093,3229,-1385,-839,-620,757,-5683,-2978,-5156,3425,-1,-13076,-12929,601,-1192,1128,1469,-3352,-2225,1158,4206,1044,-973,424,7983,2098,-5351,-6411,-3239,1860,1899,661,4174,4206,-435,5317,5927,110,-95,-7773,-4245,-5620,-402,-1579,-9389,6513,-1066,2275,2841,-4052,-4082,-898,8388,-1330};
    Wh[20]='{-498,-6962,-2366,-1527,-14,1022,3635,2658,1043,-2495,-2297,2177,-621,3083,-210,-1916,-911,1638,-1871,1039,-2941,-2004,1859,-1906,-311,-690,620,-2192,1304,-1672,-544,26,-5737,378,-2971,-2849,-4797,-1130,617,-539,856,-1726,3156,-2414,4482,2517,4372,1226,-4248,2092,1975,-1813,1353,34,4826,1254,251,-1361,-3977,4519,3298,-3112,3288,1004,3530,-326,3964,-2595,-1224,1879,2907,2895,-1861,2561,-2639,1635,-1456,-1459,4057,578,-2963,-5385,1721,-3908,4035,-1804,-112,1282,1998,1220,-2285,-5366,1638,-939,-3913,-414,444,-3537,-1945,-1520,-2998,-3911,-3779,-2761,2285,-1602,40,-2056,-1049,2182,-1380,5258,-253,-3681,-1893,-1665,1270,5517,-756,2832,983,-2104,-1936,-3105,-1290,246,-1455,-12,2222,13486,-3842,-1629,-2431,2822,2091,-2379,1397,364,-1533,1564,352,484,-1160,2312,4038,2003,-3073,5639,1813,-1439,1027,341,5512,-5229,-3493,-1423,-35,-2083,2587,-6152,-3999,-384,1060,-2963,-2526,-3554,-6494,1705,-2685,-6,-3400,-8193,-3720,7670,1562,-1877,-3269,1627,1799,2187,1766,-2824,-3215,2678,2244,2326,872,1560,-3159,3947,-2963,127,-6708,1835,-656,916,176,-1396,-363,-2454,-930,2751,349,1652,-1374,65,1356,2585,-840,242,-9794,-2583,-2368,-300,687,1993,5864,2053,-6181,-1199,-317,2054,-4331,2077,-177,-3100,-5786,742,660,-2034,-1483,6625,2871,-1070,2277,1614,2993,-505,-1876,-2271,357,6723,-4309,469,4636,1828,-3293,2293,-1113,-4487,-1860,-242,-332,-3859,681,4121,-3847,-743,306,-2778,-1106,-4470,1783,-370,3535,1818,2464,-983,245,900,3029,-2543,-4130,1492,39,3190,1029,-1342,-7192,-1240,-3452,-6289,1163,5537,2307,6059,1191,1323,4125,-2622,-3459,-2015,-1888,390,5737,99,-4504,2553,-2690,-3845,-643,-3383,411,-3166,-2041,-4174,1129,7421,1611,-2644,-2739,-131,1335,3134,-299,3071,-4829,1763,-6391,3203,-6459,268,-1588,-445,-2641,-604,-562,-3200,3242,640,-4104,-1391,5976,-1854,-3715,-2038,3051,62,-1829,1010,-3347,404,-484,2924,1050,1773,-1329,-1660,-5786,919,2368,3059,-825,289,-765,120,-6733,-10175,-1818,-4008,-2573,-5258,3747,-362,855,-3103,744,597,-327,-3725,-560,-1779,-6484,-2290,-7651,-823,3032,1571,5483,-2536,15,-2052,-1683,5541,-1485,1194,174,2590,-924,-1008,1781,2519,1336,2561,6796,-8198,-1058,3278,-6162,764};
    Wh[21]='{-440,-3913,5195,-854,-2685,-252,-528,-2573,2376,266,2270,-2502,-295,1602,-6494,2104,1832,-731,-1517,-603,-2410,-5268,-278,-3986,-1395,-36,-3676,-844,809,1220,1915,7431,-2022,-2191,-3024,-2043,-1380,1926,1706,1981,-1165,-1008,-740,-785,2425,-2553,-4289,1888,-2143,793,7729,1719,12578,896,1059,-1716,1295,2144,-2985,710,-2607,2893,-1436,-3383,-583,1243,-2489,751,1436,269,-2578,-644,653,-1083,215,1594,-5444,1336,2160,1069,2103,-1958,-535,634,3176,-5820,-84,-2519,-1705,-2646,3198,935,-2093,-675,-3325,1,-922,-5146,-2202,-2487,855,2468,-2106,5561,1420,1600,-485,1425,-2761,4467,383,-3640,-5458,1800,1488,174,805,2875,2646,-2749,-1578,-4399,6469,-2351,3371,-3354,-2186,488,3349,-2558,1705,-1262,401,-2326,-3066,-1495,-2269,-396,680,1166,297,1787,-3540,318,-4096,-556,-1334,1967,3522,406,-49,1796,-2697,-3310,-2255,4218,1715,-1712,-2490,8100,5502,3977,-790,5039,659,7016,-1032,-3381,1202,228,-5410,-3701,7187,3845,4953,587,2103,938,2102,764,214,-3002,1774,92,5830,514,886,-653,-10703,4848,-1315,-129,-731,538,-2302,-7631,-2890,-936,3081,-292,237,1867,1160,-633,-5712,885,338,5507,1256,-2312,847,-3432,4960,1068,5292,-7099,1589,1977,192,149,-266,3322,-1960,-624,-1811,-1365,514,1499,1239,453,351,2690,2634,-566,-1669,-2919,6787,1571,1883,2131,-3666,4782,2727,-944,-568,1809,1271,3178,-2048,1597,382,-4013,2714,-1395,-1591,-3361,-4624,3742,1341,-2442,-536,-4384,4123,-5698,3833,848,-2047,-3662,-586,318,486,510,2420,-1080,428,-4624,-778,-2296,-1702,2442,1352,-1871,598,-3642,-1323,-1542,1358,-7558,-2038,-1533,1926,-2416,-7104,-1466,-2393,-2070,-73,5390,1572,-4064,-3105,5654,576,2010,-4357,1052,1627,357,-178,-833,3237,-238,-5185,-3620,4375,-869,6542,96,946,-3764,-6230,-2810,2705,-1367,-5405,2895,1138,-1300,-2526,1546,5034,-753,1256,2081,-2354,-9272,-4367,4301,-2854,2153,889,3947,-1016,4904,-1268,298,10029,-1811,724,2570,4714,4291,-1013,-546,-2575,-1057,-4875,-838,-6240,-869,2042,-3193,-1645,-4382,2521,-33,-30,-1966,3830,-1602,5898,-6625,-4912,-3481,-3098,-678,1846,4072,-1696,-7299,-933,315,3232,-2607,-3723,-1019,556,-6923,2210,-3283,729,-2016,4182,-415,2653,-4235,-233,-6,1230,-757};
    Wh[22]='{1689,550,-933,4160,-120,-799,5444,2768,270,-171,1372,7592,737,1856,-3129,-2054,1534,-187,2761,1884,-1009,2661,-694,-1347,-924,-390,-1595,44,2602,-540,509,10302,-2792,1997,1552,-4089,-1678,5375,2225,-731,4326,910,-5112,-572,3317,4162,5825,8427,1557,-1732,2558,2233,-2634,-957,-1608,-2399,-5605,2286,2597,189,3122,1960,206,-1589,-1502,158,-2026,-551,-803,-559,-2797,3986,1330,2398,-3618,6958,1076,1066,-3684,6889,-802,-2839,-2086,5087,-6391,559,913,-293,3012,-965,-1022,-1301,4345,-688,4206,-999,-2056,327,2949,-17,2639,-1612,1611,6645,-1297,-2800,1607,-599,136,-142,484,-2548,-6401,2083,59,-1021,-2156,2459,1416,-905,-1462,-2048,-6040,7392,881,-2127,-1252,841,1334,1453,4633,-754,-166,-802,-4455,-1629,-9760,2249,-2568,-62,895,-51,4165,-1011,-1350,-388,-1927,90,770,-1325,-957,123,-1511,2047,3232,-1154,-282,2210,-1036,-195,-7456,-1356,1833,-2294,-4716,4035,2456,-532,-223,-726,6518,-2858,729,4306,-2731,120,-3735,-1669,1333,-1405,-734,702,4340,-1616,-2362,-7241,5083,963,-3369,-1174,1076,-2486,1233,-2382,-1343,-5458,-4228,538,-298,-1386,831,-2121,-862,4680,-1614,-1275,996,-1435,165,2753,3879,2858,-269,-1024,2519,1054,1623,-1109,3742,1683,-2109,5502,2017,-2766,3100,2059,2719,-2298,1676,2629,3886,-558,5966,-941,916,-929,-695,222,4194,-283,489,-1481,643,-6171,-562,1613,2358,-4396,1489,842,1413,-1578,-531,-1593,1949,2264,960,-509,-725,6342,-3449,-2431,-5639,2456,2067,-1896,2082,2343,-1412,-3293,4787,-3422,932,4309,-398,-9267,-1235,-4443,2059,4594,-2008,1341,4277,2663,246,1119,-384,4992,1491,-366,10,-994,1146,-2337,515,6250,708,-878,-347,-597,-1314,-8085,150,2651,-560,-295,4477,3937,-1052,3664,-4169,-2910,-2434,-2489,-3479,1256,-5063,1132,1412,3830,6723,5429,-2700,-3215,334,1407,1850,-1517,-1398,-1048,355,-228,3012,-2443,-2539,-2863,6577,7890,-1481,5239,20,4470,1517,5478,86,-679,-1540,-30,2128,1409,2766,445,1678,-5146,-2373,3544,-140,3205,373,1320,2707,4384,503,133,-6118,4194,1246,3549,1773,1868,1722,-2834,-2841,2858,-2106,3403,-1220,-3178,2287,311,3466,3393,7807,-1773,-6059,2514,6250,2137,2185,-3298,-241,2729,1687,-3579,1052,4221,-76,-892,8149,-1372};
    Wh[23]='{2824,1776,1765,-4050,414,-2800,5068,-4,1783,-1641,1015,3476,-1402,-525,4211,-2060,5732,4553,2196,741,-70,2159,-5385,-3122,980,-4023,-2077,-721,-1679,3498,2156,2171,1766,2541,-1459,-4809,662,-1934,2922,6894,4057,1557,-1015,3417,469,-1047,48,-816,2524,-2722,-2531,2583,-5732,-1124,431,4040,2700,1669,4091,6367,2440,-166,6821,515,-770,2878,-4865,1813,2954,2590,373,2670,3833,4377,-1196,927,2343,1793,354,-3808,1047,-4138,-1069,2712,1909,1530,-492,-1265,252,478,2731,-1221,725,2717,1329,-3327,2310,-1762,339,2751,-2241,4538,1624,3054,569,91,6005,7,6738,-225,-3969,-1586,-140,7900,527,143,-2445,619,3933,-4814,-605,-1706,-5532,-1975,-656,-8911,5063,803,1378,-11093,-1324,2366,-1993,-3303,-3979,-4050,3881,-78,383,1633,-4904,2551,1000,-804,3261,-4396,1021,-3513,2585,1867,-1340,2474,624,-92,1420,425,7153,2298,1190,-5922,1992,-4614,459,-8007,6196,1816,1032,-493,352,1939,-651,2078,-352,1666,2043,-3505,-1958,2861,-4477,1772,-1695,-5366,5214,-3273,3220,-709,-136,-1232,-3334,2465,-4807,-1146,-4528,2795,-3479,-2164,-2985,-291,5527,239,-3774,1564,1433,-2215,-928,-1568,444,2219,1217,666,-3815,1656,523,-1300,-791,4174,-2780,3168,970,-787,2077,2954,6679,6381,532,1738,3176,312,-3486,3669,-1051,-4421,1892,-527,6123,4416,905,-2448,828,1944,7622,-2790,722,325,-1254,1026,4272,-847,1370,-42,-1118,2954,-2244,-1206,-488,1119,5502,-110,5590,715,1385,3037,623,-4291,-6484,2337,-2069,-62,872,1221,-2500,1336,4165,893,-5468,-6889,3615,1859,-1101,1168,2529,308,-6376,2290,68,1354,-1856,5400,-3164,693,6542,233,74,2612,2770,3935,6508,5844,-2946,-3041,-438,-397,5224,-3129,3198,7309,196,-1812,1396,669,4106,1484,2502,2454,-1326,5180,1420,3054,-81,3166,3833,1411,2790,4047,1176,-369,8989,-1116,-92,509,4960,1545,1705,-1903,6298,8417,-2231,1660,-4042,-4997,2235,972,-3872,1243,4025,3403,-10781,-1882,-148,-957,-493,952,-2250,573,1762,-2829,6791,2968,4772,-907,-2600,2739,1459,-2714,-4987,12314,-3415,-5048,411,2937,-1162,-51,2202,4729,-5561,2066,-4150,1832,2408,5278,6987,-386,-2873,85,2364,1156,-96,6738,3103,61,698,-4770,6723,-2042,1497,-3522,6479,2810,9570,346};
    Wh[24]='{-942,2512,771,-1721,2481,-1436,2556,-4997,7177,3352,-415,188,1139,-3745,4541,3935,224,1478,-1524,407,-1323,983,-1829,1766,1508,-247,-2824,2517,-1163,-1950,-2042,-781,478,-707,892,3276,2937,2219,-5688,88,-1253,-1484,-10205,4255,-4533,-2380,-2458,1291,-1055,-3493,1987,-3183,-3022,-6542,3095,-2081,7226,-3024,650,7729,-1437,1612,-1940,4489,5439,-1248,-2807,181,855,1333,-2915,975,-4519,413,1842,-403,667,786,420,-217,3708,512,-3300,1718,-612,350,112,419,1341,-318,2778,3481,490,-1281,-2380,1300,377,1002,2458,-354,-344,29,2135,-537,-3923,149,-2390,-4379,2440,-900,-211,1634,2354,-3859,2011,-1386,-679,3215,8720,3457,-3740,809,2514,3937,-2121,-2629,1339,-1551,3952,-1629,652,3046,-1317,4326,-1920,4853,7861,-1429,-3342,-2308,386,-731,-1211,-188,390,-1572,-2832,-8139,-409,3999,2332,-1503,6909,3557,158,-566,-5708,958,-6806,-1652,-1386,-1423,-2741,7070,-1590,-1156,4172,3527,3007,-523,5312,-2315,-1099,-2502,-1003,52,2130,-264,-2753,489,-4189,-406,835,2072,-1385,-2551,-3481,-461,1784,-1027,-1077,-3161,-2282,1406,-534,4978,5097,4218,-144,-2436,-2272,-969,2539,1619,2130,-1055,1567,2578,-2663,2172,2836,7768,-438,1418,558,-2492,-1964,3254,-996,-1947,-375,1004,1900,700,-147,-1856,4033,-483,3876,-1474,1328,-10009,1213,677,5844,-392,-4208,-955,2336,5859,2841,-3491,-2185,3371,1785,1270,2025,0,3857,-5429,-3947,3698,-4831,4829,8403,5361,1865,-4780,2802,-1418,187,2104,2172,2673,-7407,4340,561,2614,1376,107,-1932,3894,-2207,1914,-1097,-2993,8754,-561,1345,1075,5175,-501,3784,-3796,1920,4091,2016,3547,-5654,5927,4204,237,-268,-881,-3059,2685,-1715,167,144,2224,-1531,-1801,5004,139,3134,100,4489,-1739,947,2832,789,-334,295,-187,147,-784,419,2558,-1385,988,4042,-1269,-2247,-375,4931,1295,1506,663,-2180,-499,569,-308,266,53,-2912,205,506,-3251,4458,1806,3986,1068,-927,209,-3425,1392,4025,4184,-3461,-556,2639,-2352,-191,2419,652,2929,2125,1436,-155,-3698,437,-343,1295,6791,3706,4152,-7080,3710,1632,2185,-6254,302,4204,647,-1142,-1270,-477,-1106,2595,3078,5532,-1469,2283,-1542,5698,-3015,2102,2849,1039,1727,3520,-2292,3566,-10507,-7470,3896,-83,1595,6743,-632};
    Wh[25]='{-64,-494,-1726,38,-1181,473,187,1046,-3044,798,-3015,4372,3845,-3063,2727,2573,-3476,415,-4309,825,1301,-2856,1649,1132,3466,3032,-5825,-3330,393,-1430,3356,-4860,-991,1209,-2814,186,123,2683,-785,-3051,-6538,-1080,1017,-4638,-1623,-5048,-54,-2739,-1297,4562,-2341,2895,5185,5327,-1823,-6079,3054,-388,1873,1135,-365,-4418,-180,330,-376,-2509,3193,1082,-1667,-6562,-6000,-2705,-5952,1652,1810,5458,2047,2298,-2130,-1129,-1083,1222,-1938,1270,3754,2158,574,-5541,-47,4125,-2839,-6782,4301,-4643,-1804,2001,-296,-967,-2291,-2810,-1067,-5268,822,-8100,-1027,-196,2583,-698,13164,-4858,250,4228,4338,-2692,-2264,-2634,-1879,3618,-1481,-235,574,502,2668,-2053,-1556,-6088,5185,-1572,6206,2286,960,-348,-2128,-2651,1066,-433,5712,-5917,-1966,170,6079,-333,-2100,-1260,830,1625,-1002,-121,3488,2612,-303,-3447,-3439,5776,-4240,-3972,-2103,723,-3481,1542,2399,758,715,902,-3715,-4777,-377,-3176,-3212,779,1376,776,-4633,1005,1992,4704,1441,238,853,-562,-2670,-1802,-1395,2526,-3110,2137,-4726,3017,2474,-4379,-2322,-823,7773,2092,1923,4396,317,387,-3906,3237,-392,-805,328,-139,4960,-396,-2919,-3818,-4267,-6186,44,-839,-1024,-1636,225,2482,-3767,-3356,-1138,-1691,-2966,23,-3359,-1577,-1580,-2697,-2272,470,2939,626,3554,451,-1190,-1297,-3925,3081,911,-5327,2729,-1781,-229,240,-47,947,2587,311,-4367,-4768,-361,-1025,1756,-2349,563,-4353,-1143,-132,-1149,-2773,-1402,-2347,949,3747,-2464,4023,-552,376,3229,-2866,308,2558,4365,-1094,-795,-543,2014,7050,-3215,2927,-55,-2521,-3967,-969,-1293,1229,-1054,-5239,-1635,-5756,424,2357,-2614,-1529,-37,15,-2492,1291,1131,137,-2744,4523,-1734,631,-745,-1273,3769,-3061,-2158,-447,-1551,-5771,-504,-1015,1340,2958,-3891,374,-8652,-232,-2033,5493,-209,-203,-3479,-1459,-5668,-948,-2310,-3205,4567,-4057,2432,591,1586,1883,-6318,-193,887,-2373,4072,4470,-988,-2314,3850,-6933,-1627,-1302,-63,3610,3359,1102,-2749,5517,-1740,374,-4555,3325,764,2010,1374,2315,-405,-4497,2102,3564,1573,2878,631,-191,1430,-4440,-2197,-5561,-1112,1489,2661,-2441,5043,1472,-3793,-1768,-4160,-1679,-1995,-1711,-3894,-2291,-2849,-4963,-3581,-3452,1140,1776,-786,-823,4094,1077,1337,-911,91,143};
    Wh[26]='{-913,6176,2734,-1777,2149,-1712,-430,-1312,-1325,-939,2014,-730,2034,1665,-3662,-473,905,3312,2144,-788,-242,3920,-1934,807,-487,-23,3347,-2304,5634,-8261,-1876,-2966,-2071,3833,4130,-1138,2128,328,137,1096,37,3122,-2158,1148,533,-68,2318,1274,-3239,2000,1840,-1406,-3200,-2861,-1800,2539,3144,-5937,-4272,4211,241,-6733,852,-384,3330,-18,-375,-602,2639,1293,2148,-1291,-2846,-2084,2673,-1827,2746,1750,1713,-1225,-156,-1510,3078,1078,-1727,-2834,940,-2239,-252,-326,2905,-120,-1237,-3149,-1183,2196,-467,-595,1060,-1507,-1892,462,1479,-1850,2985,-244,3164,-3859,4577,-2602,-1038,3371,-7797,-3820,4797,-1611,6303,8852,4055,-1950,716,5302,-4797,1340,1516,-91,-7905,2966,-3896,-2352,-1183,3730,-1246,493,38,1470,4855,1102,-337,-5185,-1748,1069,-3823,2595,-29,-13,2061,322,-2288,1879,4602,-693,-3957,-1230,986,-7231,-3898,3081,-3205,-2442,-9184,-1419,-3955,3547,2644,3012,-2419,-1706,687,-2719,-1319,5048,-4687,1036,3723,1900,5195,-2362,368,-3183,130,3107,-2758,521,-3579,-320,-4006,-3566,-3920,2448,789,-3732,2536,-2749,872,3835,-541,-2318,7324,-386,-1556,2907,-1851,263,772,-849,239,-1889,440,239,-5268,-1112,-1478,939,925,1205,-611,-905,-5908,-5893,1394,1354,2175,1871,-4699,-2398,-3039,645,1357,2247,-314,1414,-4423,-1203,-492,2778,2106,-1483,-1582,130,-4191,2410,-6577,-2890,65,281,-7451,-2412,-3681,-4299,-1240,-2692,1663,-4865,-3454,-5400,-605,1013,1156,542,372,2486,-1447,-2492,-3010,-628,1148,517,880,-2561,-3767,179,-2100,3435,-5776,-1682,859,-559,1181,212,3430,-4472,-2836,-3115,581,-1890,-2113,1959,-656,-5371,3759,600,-6284,-2130,62,-709,-3999,-2083,-9741,-2834,2044,326,-4101,1672,1437,809,881,-1595,3496,2009,-1212,-473,-556,-2088,-2834,-3420,902,-328,-1354,7451,20,-4702,-2604,475,-374,565,9008,466,-6015,-834,-807,2753,-3132,-2587,334,3515,-1373,-5629,-1030,1928,2036,-5708,1549,1362,-917,1367,3752,-4841,-969,-3664,-1428,-3361,1427,535,-1842,-3774,-3249,5810,833,-2208,1614,-1865,-3798,1101,1247,-3862,-560,9057,2270,2110,-177,-494,-2788,498,985,-1364,2534,1781,2220,-3188,-1333,2153,-2717,2264,1807,-3505,-1115,4587,1933,-2008,3459,5434,-5688,3662,-191,816,6455,-3041,8374,-1425};
    Wh[27]='{-648,2390,1024,-643,1619,-969,-5517,-4270,42,2335,-497,-321,1280,387,4313,-4350,-817,-3317,-1868,-1706,1350,-3798,-876,1176,2578,551,-508,-1008,-1871,3007,2,-947,-851,-1545,4416,1884,1944,825,-1625,-3020,2531,4409,-1726,3833,3750,880,-5234,612,-304,-2885,-350,4567,-3068,-2163,-3125,-586,2666,-578,-1085,-2185,-2995,1650,832,1671,-425,-3293,-233,1711,1180,-359,-1942,918,-907,-776,2849,3229,-1222,-6059,-497,-4050,-2058,2761,-1215,3505,446,1772,1555,-2553,-2746,-1412,1477,1119,-888,781,-3996,-17,-1469,-2435,2001,757,-1594,-2196,-775,-1058,-614,494,783,-5629,1616,750,237,621,231,1551,-1728,-1707,-2009,-4130,4313,-25,-837,-444,-1066,2924,-376,-1888,4328,-1716,-95,-6489,-345,2495,-615,232,-4956,-1657,2587,-1202,4509,1146,2814,1837,-1755,-4079,218,1739,-2340,564,2238,-3225,3242,594,-2297,-2993,1368,3017,2003,-513,2006,-2800,1936,45,-2497,-599,-1918,154,699,1756,899,-665,67,2214,-2054,-4382,138,1105,2189,1016,-2641,669,-2487,-3625,-1024,4978,62,3312,3212,3286,1783,-3288,2695,1813,3630,-5522,-3645,-2202,-3601,626,-5537,2016,3513,-4741,156,-1967,1172,394,3278,-3125,-3632,1370,5068,1031,2239,-2440,2384,-254,-2253,2172,2856,-4711,1627,699,1983,453,-1177,3710,1614,182,1520,4062,1273,-5590,1540,-993,-9599,-3205,-313,81,-2429,-203,1098,-7187,2052,-4890,-3063,1083,-2810,-1071,4104,3977,3315,4152,-1282,3823,-5732,-2478,993,1446,3059,3276,1017,2749,1291,-1942,-1209,2463,1228,-2141,-921,-546,3701,4321,410,-673,596,53,2797,3730,6088,-1480,-158,-4133,-907,-881,-87,3090,614,314,6191,3259,2995,1599,2364,-1600,-3376,-3256,-2553,1918,1527,1224,2,1490,2834,1536,957,2739,2015,-4184,-2487,5317,-819,-476,4001,821,2292,2194,-579,-4687,1716,721,996,-999,54,-1447,-1683,-2230,362,5288,809,-321,2895,4453,1171,4301,655,3483,-2497,291,2871,5375,3430,2917,-3686,-8120,238,5004,-1084,1447,5747,-265,-2512,1610,637,1538,-668,-603,523,9589,2617,377,189,4838,1702,1296,97,-2414,4387,4042,4821,4343,-6489,4340,4250,2093,2910,704,1201,-648,2291,1083,-155,-100,593,3615,2680,149,566,-339,3190,-1503,650,2199,783,-7475,-883,1459,-1734,1684,2191,1264};
    Wh[28]='{-1152,1925,-1087,3854,-2073,1480,10009,-2333,4963,-2003,6044,-4870,2692,2680,3623,5429,-2192,-2426,4055,4040,3835,455,805,-186,2993,3156,6694,-731,9360,1702,2595,-69,1406,173,-3125,3664,-5585,1501,-3186,-2048,7182,3469,1773,-330,-1093,-429,5170,-2602,4406,-3994,7192,-2512,-1242,-5727,2059,1098,-4062,1237,2543,-3508,-5595,-4130,3310,277,1333,4895,-2479,-1624,-3237,-1403,3662,4499,-1340,1704,597,-2043,-1326,5312,3847,1896,1778,4001,3298,382,380,-1843,2135,4111,2973,287,-935,-5009,-4399,-4572,4826,2609,4274,-483,5678,-1445,-17,3691,1108,-3349,2531,-800,2053,3286,-7734,-3535,-6196,-2561,-2961,-894,-2651,-837,748,5073,-2597,2839,650,-164,7651,4826,-7202,-6157,1144,-948,-11074,1531,10917,2514,-1514,-2327,2048,-3725,-722,-3325,-5073,1302,-3911,557,4592,-580,979,-4301,5278,-9511,-3476,-5156,498,3813,-2712,-3156,6909,1633,-3171,-1303,-2145,6704,-2597,3081,1166,8730,-3386,-5356,3403,2126,432,-1089,-573,-1098,-6899,1796,2120,-2343,-1499,2160,-2446,2985,726,196,529,7509,-1318,3300,2473,2249,-9345,114,-974,-287,10849,-2272,1243,3400,1468,20,1940,4038,-852,3820,1405,-6,3525,2680,304,3520,-1771,1948,-2646,379,2014,1613,5024,3503,6367,2468,5048,3598,2133,-1374,4426,-2222,1528,-494,1466,1987,-7851,-369,4187,2580,3608,2644,3227,-1890,-4645,2418,685,-1934,-5893,4204,-296,147,-4340,918,-2215,-4606,5307,-3476,2531,-1922,3024,-3503,-2272,527,5449,-5771,1842,3239,1883,1997,273,1586,2687,6645,-212,2052,791,-2797,2072,-6669,947,-392,-5053,3188,-3977,2846,4570,3107,-430,-1384,4902,-2377,5957,-1008,3403,722,-1857,-2673,567,-3740,-1881,-1665,2067,9516,-7817,-2308,2409,4404,-4301,6284,-1849,459,-299,-3181,11298,449,3464,-13,-1433,-1057,11191,-3947,578,-6313,-1578,-1602,11640,14677,-2016,-166,-2722,1453,3342,89,-4470,-3588,1375,3015,3181,-3122,1293,-3718,-6367,3249,1169,-728,8784,-1022,1694,-7651,-4882,-3554,1290,3354,6347,3666,1403,-3520,-143,2401,-2629,-3156,-1691,4821,-1135,-1444,4123,1506,2792,6293,232,512,2375,-4372,-5732,1950,657,-6289,-3881,2807,-2580,-1340,816,5913,2995,929,-1336,2163,-1112,2176,4838,-7661,-3615,-3659,1666,2128,921,-1632,-1523,2425,755,-3020,3535,1214,-440,1475,2814,-277};
    Wh[29]='{-936,5561,1749,2658,-318,-3571,-1483,-21,528,401,8593,2302,7368,2370,-2320,4426,3981,802,400,-2983,-1540,-6689,4160,7089,90,-1341,2504,-3120,245,-3771,-3913,-1202,3696,811,-2587,-1114,-4719,1524,-2741,1445,-3508,-5986,1759,-1795,-2683,-1302,8676,-3649,-2248,4367,-5146,2812,-2249,-1560,-591,-690,3930,-13007,2978,-1798,-1875,-5234,3481,-1280,4462,-1878,2902,1085,-2954,-154,-6596,-5781,-411,-2580,-888,5097,-855,-1627,-5952,1907,552,-8364,5644,2152,348,-436,-589,-563,-3122,-15263,-117,-217,-154,-2990,123,1900,398,3691,777,316,-3317,338,1912,15712,-2279,-2482,2392,3872,772,576,2880,-7636,6420,-620,3012,1043,-4140,257,2512,225,-2934,-9189,-3598,-2502,681,16250,-3037,-1903,878,-6005,-12724,605,-9086,-69,3732,10068,-5639,-4331,4938,1467,-4533,785,723,-1093,2922,2272,-717,4582,4804,-6611,-1171,3103,-2922,3063,-2993,1333,-195,3662,-4118,2320,1557,-484,1696,4921,3312,-28,3498,2639,3610,316,-4218,-2790,616,-121,-8403,-654,968,6567,5498,2451,1811,5361,-1461,-3107,3134,3466,5371,1975,1132,-5698,806,-285,-5854,-539,6484,-5004,-64,499,5205,-603,-814,1337,-867,-6562,-1844,-2763,408,4851,-1252,-1633,-1257,-372,-10605,975,3000,850,-961,-73,-2480,-2902,1668,3410,-5834,-1595,2407,-3659,-4926,-820,-3059,-5966,-9018,-1045,4414,-5014,-3015,1352,-1302,1932,1218,723,-292,1770,-527,-5883,1132,38,4599,-3400,831,1848,-1765,-3105,1518,-5297,-6733,671,1835,-9775,1945,-3325,-9746,11,847,-2294,3476,714,-473,-2137,1342,-4421,-4362,-3520,-357,-609,1185,-7202,265,-3476,1240,-1776,618,3977,6132,-5683,-2575,-10556,-739,-1527,-3937,1697,-6899,-4138,231,626,-158,1168,1708,-9658,559,271,-1979,-10996,2282,-791,-760,-2578,3618,-2963,-3371,-2293,-3234,-3444,-4355,2028,-7768,-1414,11337,-909,4582,6396,-69,5585,-5195,-1795,237,1878,1462,-1427,-1748,-933,-5634,2325,-4926,-9360,-359,4003,-635,-4934,-1319,204,1295,2362,4069,1853,6254,-2634,1403,-7495,-1752,3125,6586,-2279,-6,3769,-1095,1953,2932,-5458,-1120,5366,-3515,4301,-2424,-3562,-6049,-6757,-732,-4226,-2932,1362,985,58,-4567,1823,-2673,-51,-1711,-358,-600,-1911,-3652,1271,2082,-2391,2419,2078,948,-513,-1027,3327,-7060,4814,-5991,963,-8666,3535,2587,241,2150,-5634};
    Wh[30]='{2841,-913,228,2937,2810,-2393,1484,-4790,-1542,-287,1950,2257,-2170,1286,4855,-682,-2958,-429,1789,1782,1739,-2401,-6767,-574,2001,1456,3376,-748,1100,-2047,-2271,6118,36,1350,-1784,1456,905,-1291,1049,3598,-147,-713,-3068,877,-3581,1004,2795,-1290,745,-4479,-3249,2941,-4335,-2963,-935,4978,-1428,2736,-3745,-555,2736,551,-2321,1907,5698,1071,245,1166,-1976,357,3498,-229,3442,-1578,2111,-830,3796,1617,-4294,-551,456,-530,-2064,-1234,-4533,854,3513,779,3920,1832,1086,-282,4228,-97,-1099,514,-710,3937,-1523,2169,-1960,1330,-1529,13427,4011,336,-1412,-1855,3129,5151,-4423,-1693,-1868,5615,948,4343,-2717,1556,-1820,-3566,-1959,-287,1909,-5976,746,-2541,-4396,1439,-3015,3989,-7382,764,-1398,-3928,-5302,-6708,-2360,3569,-3776,375,-2546,1306,-3925,2327,7207,-4365,2539,-3674,-234,2968,-1790,-3674,-751,1658,6523,5537,-3762,-411,-1027,-637,886,2183,-12,-7822,-1782,5400,-1640,-3547,1851,-981,43,-1434,7905,1000,-527,1149,-5571,47,1296,-2714,-814,3630,-1431,-2509,-953,949,1861,5937,-4882,-1215,-1116,2705,1669,-3457,-2286,-2546,2308,-2666,-1402,-7075,1066,493,1333,-1597,-637,-39,-561,5922,-2005,2836,4401,3442,2371,-2370,2147,884,579,1500,2775,2292,2194,5146,3281,-2003,3225,-1077,736,497,2675,442,-485,2406,3132,2376,-470,1111,-1181,462,-123,3789,3166,2600,3942,18,-2751,957,3823,-5332,646,439,-777,1074,822,5786,-2678,613,-431,1876,1804,5937,5776,-4277,-4489,-616,-1400,2476,25,3552,-914,-1085,2492,2783,-419,819,1627,223,-442,2093,-31,3789,1489,616,-2152,-3425,2484,3381,800,2966,-137,-1691,2692,-6450,4028,1419,-665,5058,-393,692,-14,-2363,3305,690,4604,4716,2373,4482,-141,-487,505,-914,-1623,1914,75,-4421,316,4514,6616,-1314,-152,-2617,3825,632,-3950,-1711,4660,2829,-1722,1392,465,127,-2272,1423,-180,4050,-135,2587,4035,-22,-250,2326,2434,2314,-2403,-755,1729,2062,2531,-797,2200,-717,7495,753,1761,-978,-1702,731,475,1822,-1704,3352,8505,2130,-1146,-1695,-2180,-524,1562,-162,-1835,-1057,4975,1342,-55,421,4914,2773,-218,-1157,-653,1326,2946,359,-733,3876,-2670,-2636,5952,3693,1235,-2670,233,-3603,807,3793,-1730,4838,-4177,1403,406,-1301};
    Wh[31]='{539,-75,-380,-2418,94,-226,149,9624,-2604,-4133,2220,542,1148,-1866,-2122,-1556,1905,11,655,3796,-242,-1456,-1267,-4123,-1196,1150,4909,3117,93,1767,722,-7895,701,309,2277,1662,-2387,852,1315,2592,5664,405,-2766,2983,199,725,-2739,3825,-888,1553,1135,3803,2734,3376,1651,4868,1328,-208,-1611,5419,1617,-345,2254,3903,3037,2137,-6826,-4020,2231,2320,-5200,8481,-1021,4260,-5039,7714,841,3264,-608,2324,-247,2561,8789,-5869,-5122,5092,-3283,-2213,-1152,2573,-244,5991,4157,664,3317,3117,-1005,-2047,164,-3576,-2431,-6250,791,-154,-2807,555,-3784,-3991,-1447,-3808,-2968,10253,-5815,-2895,-946,-3764,616,5595,8925,-2447,3112,7343,-2382,6757,7939,-7807,7705,-26,-6293,-2269,1713,6206,-5263,3793,306,-4538,474,2517,-4821,4157,-1004,404,-3449,-4189,-3732,1241,252,993,4648,-2807,-1966,-4953,-3557,-866,-4108,-6074,4367,-415,67,-11083,-4162,1357,-2770,717,715,10224,3845,6025,-1813,1673,-1859,2456,-258,2266,-4638,-3166,-1790,-3176,-4353,1656,3793,-6918,1166,-1413,-5136,-1862,5283,329,3051,3859,-1761,-5537,-5395,-2663,-1348,4804,-1705,-4211,909,206,18,-3239,1761,-3022,-5517,957,484,408,2225,-3828,-4770,-3950,-651,6411,-1239,-885,-1308,3881,-92,-339,5068,5839,-4411,-1771,-1988,2282,-4780,4453,3232,-2351,-2304,-1182,-5478,-1646,3955,1176,-2307,-1748,-3103,-1113,833,115,-3698,1639,-1759,1691,-1566,-5297,-3818,-1087,-4042,2690,1840,-4025,-1428,941,602,-2368,-2658,-3537,1169,-353,7070,-3640,3220,-2976,-1072,1212,-730,1264,10,-1883,-747,-4047,1211,3149,1202,-7895,2023,2010,3234,-1424,1793,4665,-4265,-3559,3320,254,58,1018,4902,-812,3251,-2673,-230,-5102,3222,4226,-2453,-761,1401,4172,1336,4741,878,6845,2858,4885,1451,116,-1259,-4438,-3071,-2427,1503,-296,-489,-4003,6694,3935,3095,-806,-138,-5942,1375,-5405,-1636,2104,1159,597,-7207,4643,2958,-1050,78,-2132,-3413,5214,-5366,-3688,-960,-3249,1188,5253,1555,4497,-2917,-3239,-4323,-21,5000,3825,-781,-5341,-2563,1392,-7001,-2307,7148,-3750,1323,761,3129,412,-2136,-2464,-3515,-634,3911,-3930,-497,-4030,4909,681,-2185,-3020,6669,-2614,4704,4362,6518,-5546,5307,2460,3061,5146,38,5883,-280,10322,3283,1042,-6440,-482,3806,529,-2069,-54,-2362,-1672};
    Wh[32]='{-2254,-9633,-1667,-3422,1873,-1373,772,-6318,5107,40,-3620,-3527,-7890,3659,434,4008,2807,-574,-3225,-1120,935,1166,-222,1320,-506,-3088,-112,-657,-10244,-802,-2875,-5727,-2880,-1596,3681,-2277,605,-1353,-4235,963,-10537,-1495,-9594,-5488,-4587,6010,-2998,-2573,2717,555,7290,-793,-4399,-2783,-958,-3395,-2602,-787,-6240,2749,-414,-5419,-313,-3188,-2702,1743,-2373,-3342,-4692,-5024,1510,-1442,-5966,1379,-3598,-5766,4606,-4914,4348,1857,-218,-2200,-1267,480,-407,-839,-2702,3515,-3828,1984,-2775,-1990,-10175,1496,-2609,-1243,-1251,1708,206,-7617,2474,5585,303,2880,1403,3049,5092,5146,2727,-1483,-4064,5820,13310,-3818,-4580,1973,1450,10849,5068,12,3256,3173,-72,4289,5639,-8432,6953,-677,5771,-2756,-2729,-1000,-6044,5673,4230,-6176,-316,3137,2377,3281,123,-1625,-687,132,-1165,-3847,3654,2283,-4809,3347,-2048,-1017,2255,-5258,1938,-16103,3049,-603,6440,-25097,12089,2846,232,3676,2469,-13076,-4694,-552,3784,-482,-659,1279,-8217,2072,1518,1342,-507,889,498,-2147,5786,-2546,-1247,20,2626,-253,-2893,7065,11572,2687,3093,-764,8750,329,1049,-935,2553,145,-45,-150,3786,575,1138,4191,-2631,-253,3969,-2512,674,6977,-3945,1201,5668,2822,7182,5483,5922,2844,-1198,3681,682,221,-1412,1563,2489,2736,-5854,1065,3166,772,-2846,2812,4704,979,-708,6757,-1744,-314,-6660,1228,6142,-257,-744,-9023,9125,4558,629,3417,-6567,-1077,-669,1571,3906,4714,3750,2580,996,2435,-4038,-8564,-1237,5249,1058,569,867,-553,1953,-2463,-2420,678,357,9047,-2580,-41,-1489,-276,4125,1845,3168,-368,1757,1390,-446,6250,-1334,2556,-4504,583,2998,3312,-1839,4145,-2286,2827,1491,-796,-6333,1661,-3615,3891,5649,2849,-2678,7866,1418,-10898,-2299,-2126,-701,-2056,-6264,-4736,4516,9746,-6191,2541,3525,-2410,-9897,3190,-2858,2636,-2954,947,1251,2434,-5053,-2250,-4477,-1943,-734,-629,1171,3754,3710,13935,980,-7895,-2453,5458,-3554,868,1004,-3527,-676,4602,495,3874,-16113,-148,5117,-1025,-1614,-1337,3666,-900,-3803,2556,-6748,-857,6733,-2044,3291,1890,3095,-196,-4516,1468,111,-1268,-350,2150,-10048,3732,5034,-3095,1995,1052,-86,1473,668,7548,-4035,3657,-3251,-253,-5117,-2369,1844,-2846,2164,-4,-7500,798,-6113,-2102,-5195,9028,3627,3188};
    Wh[33]='{717,-8090,-857,-1063,2651,-261,6816,3991,-2824,-1931,-1209,-4699,-3244,-1467,-2910,3208,-4694,3498,-317,-2573,926,3002,-1690,-2056,-1042,-2902,-2152,1023,-7866,3967,391,-1594,1396,-3605,-4741,-687,-248,101,-4523,5058,-303,1402,-5263,-521,4323,3562,3752,7099,-3000,-2714,2199,5952,-64,-5947,963,3173,115,3232,-247,-12832,1756,-155,-2330,-1015,-1097,2115,1628,-3627,4501,-3757,1959,306,2292,-1171,703,3405,-5000,-1387,4343,-1749,-1340,2344,3952,-637,5180,1926,-4541,819,2998,245,-462,-2475,2181,-12539,-2315,1483,-3168,-2384,2429,1661,1007,1270,-809,-5351,2990,2242,-59,5244,-8657,5581,3132,8847,-2003,2575,3657,3078,-3139,-5092,2386,-3295,2880,626,-5156,-5180,-3146,-2471,650,231,-6108,1970,1857,3757,2426,-9028,2641,-1727,-1601,1527,-3967,-2045,-4899,1606,-5024,8198,5205,-1159,-1751,-689,-1008,-4433,-1026,190,-4433,-3786,-1009,-1657,-2756,-3105,-5126,-1525,-12988,-221,-885,-2751,42,6997,769,-5917,-431,1195,2150,2161,1837,-536,1027,-3122,-3969,-160,1962,-883,3942,-2381,-2614,540,585,-2551,-4887,5048,-6982,2475,-1109,157,-483,-3605,5424,-13427,-622,5708,5781,4384,1339,1503,-2077,-5488,-6044,492,-61,-257,1384,-1718,-97,-1756,-6762,8017,-486,448,2143,2531,-613,1264,855,2489,-7680,1560,-2065,-6440,-2526,-2844,-6835,133,247,5034,1373,93,1386,347,2922,-2071,-3400,3435,-2912,1290,-1671,6601,1260,962,1732,5522,-3095,1567,-2849,-2239,-4226,2578,-428,6093,-6806,1345,-4877,8427,1992,-506,-2561,-771,5825,-2443,-640,-3701,-372,-1462,6953,-3669,733,-5952,1536,-2078,-4523,2524,-4340,130,-4138,-1607,-1900,-3789,-4760,3532,-3251,-496,-1994,-2454,-1921,1198,-6171,-2268,-2663,4294,268,2429,5488,129,5751,-3708,-4890,-661,-746,-6445,7299,916,435,-421,-3879,-1779,-5073,5712,-4660,-250,450,1525,-1569,1220,-8325,3562,562,921,5053,-1805,-1662,-2719,-1258,4873,5068,2424,6586,-428,-2182,-8295,1154,720,2022,1039,1938,-5664,18,7,179,-6064,9467,108,1960,-223,4252,2156,3544,-4699,4458,-505,-3383,-424,8178,-245,-2539,-5947,-324,577,4904,-5092,4938,-4821,-3000,406,-1849,-2788,2893,-3586,-53,-6279,5615,-7436,3242,2419,-1455,-5996,11816,517,-6323,4179,-2407,1278,1646,4445,2956,4992,2910,-88,1030,4433,-3989,6596,-1168,1612};
    Wh[34]='{-3029,339,415,178,717,-122,1199,2863,1738,2692,1136,1916,-4658,1738,2170,-2829,4169,2624,470,2617,3244,-1595,-1428,-445,-3376,67,-173,-3193,2368,-5668,2449,1622,1115,-2995,7207,317,-12773,3664,232,5063,792,-1094,9,-516,-4055,2675,-6762,1462,-1763,587,4833,2492,4450,58,6435,-5693,2067,4187,-1448,1955,2783,-2309,3730,1069,1623,3669,-3901,4218,-3298,-3837,6816,1990,1729,-2272,-1778,8598,-1005,4238,6586,2683,5688,2651,-1335,5878,565,6806,-3149,1530,-2927,4116,-833,7651,3447,4218,42,-191,-1295,4372,1403,2133,-1236,1422,5239,1029,-4677,1762,737,6660,-10712,2086,-1312,2192,1154,4621,-2026,-2211,923,687,3405,-109,717,-2709,-574,1232,-1320,-7675,1114,-5566,146,-2233,-1519,-74,3354,897,22675,2147,-9228,6464,-2785,-43,6406,1959,7465,61,-4279,-5737,-568,-5087,-2247,2468,-1586,2558,-2132,4318,-7182,1776,2023,-1024,1372,5288,-3205,477,3769,5263,714,-5869,2355,-3806,4267,-2370,9853,16,-6430,-1235,805,360,6684,-3942,2958,-5229,1392,-1857,963,-1699,267,-1975,1010,-515,-6708,1571,3073,3603,172,539,-476,8002,5341,1470,-1719,-4868,-3981,-1450,-412,870,787,-1044,-1229,1796,-1602,4121,-5756,1101,-4504,-1821,-2851,3466,2108,-4199,1427,5014,1226,5219,5219,1054,2153,2479,4792,-596,-4128,1800,507,1892,1578,2624,15458,16767,-865,1450,-273,-2861,-6259,-118,-2951,2861,1354,3232,3347,-745,-4333,-2868,-122,797,-3571,-1851,1611,-11064,-2271,4636,-1412,-8256,340,-1796,1379,-1431,4230,8666,-6152,-2604,808,-2333,-4077,3107,262,1130,-2369,-1508,394,-2360,-10742,1100,7011,-5322,-5502,-1069,-676,-2683,-4169,-340,3681,2178,938,1718,3803,-2105,-5141,905,393,-728,2529,-4877,-7749,3864,3901,1658,551,-578,422,1531,7319,-2420,-3469,-1939,4311,3000,237,-10605,9780,4724,6997,1979,-1367,4689,4304,282,1198,1256,3430,-1275,2145,-2570,-3139,-4780,2827,-7480,-5922,5292,1006,994,1610,-3872,-6782,740,-6127,-6752,-4455,6723,5258,-778,733,-5830,11064,-245,1234,-3481,-2526,9072,2082,-2188,-9091,-1218,-4750,-402,7705,2436,195,-511,3786,2004,781,-3588,2580,-3598,-692,-4208,3613,-1578,6918,-2427,-3305,546,56,7871,2324,1336,-3151,4431,-8212,6826,968,4777,-1539,-4028,4199,-2364,-10771,6826,-896,-100,-2174,-1105};
    Wh[35]='{-3591,-3715,-1462,-1607,-1612,659,-1298,4685,-3417,-2731,4160,352,-991,-795,-112,953,-4291,767,-2381,4997,-599,3791,346,-768,546,-2034,1171,1133,-2070,152,664,1756,-3620,-550,-1790,-979,-2434,-1721,-2341,1445,-4458,1102,1369,1612,4433,-3505,-2191,98,1402,4294,-3745,-3630,2226,1155,-498,-3769,-2841,252,101,-8549,-2946,-2391,292,-1887,1165,377,567,-3803,1296,-2734,4274,3054,-2283,-2932,-1034,2819,340,-1809,1466,-1973,-2661,671,1593,1206,638,1619,1950,-2985,-4033,3908,-5180,-6459,-2890,1373,-509,4775,-971,4050,1757,-938,3903,-1667,-2912,-7763,3745,-186,-4545,-3974,-4655,-355,1225,3696,5268,2587,-2073,-4079,2,2144,-3852,-1373,-2561,4938,7656,177,-5546,-5957,6757,4035,2866,-1435,8486,-3103,-1831,-3833,-2152,2644,7177,-3249,-286,3176,-1068,2188,-1420,-1389,1606,1955,8032,0,-204,-1904,5107,1925,5747,-1289,-3977,2993,-4233,287,-526,-3085,-4787,2049,502,-141,2790,-6083,-2105,602,-383,1185,-1417,1137,-8242,-10,-162,-880,803,641,982,3981,5976,-1851,-4211,1997,-566,3872,-2229,1778,807,2071,-5585,-1348,-693,3679,528,3176,148,-9282,7924,5800,3376,-601,1259,5415,-3771,1472,-1003,-4455,-9599,-1496,-2167,-3764,-2340,3264,-1025,-5253,3344,-1489,-1481,-2897,1951,-1135,-601,4865,-1091,-2055,1550,189,-3293,1250,255,-2536,-7500,3886,-3583,881,-429,-97,2536,-1209,-2568,3203,-6127,-393,-4323,2634,-5717,-1572,-544,1687,-4150,1970,-1838,1063,1953,-2493,973,-2805,-3288,3391,-713,-2722,-2458,1739,-4843,-3027,-944,529,-900,-357,-113,-55,-2524,4384,-2824,217,-1572,-2069,85,-725,1079,-946,-914,2824,-1124,-3212,4167,-1547,4660,1546,9741,-1978,-471,1812,2421,-2573,-4965,-12,3898,-359,1439,-1195,2086,-2454,-2338,-3193,339,-9672,-1019,-3459,4206,-2941,-3640,858,1183,-3933,3632,508,-4333,511,-18,-1033,-2670,5195,1569,1700,-500,3010,-648,809,-1875,749,-8,-1178,1106,1882,-960,1090,434,2497,-332,-5576,1594,2440,1078,-3618,4465,-2298,158,3488,-707,-4057,5166,-3300,1001,2995,-935,1903,803,3649,-803,-938,-2568,-1522,449,-4538,4504,-540,2856,-955,-3588,-1822,-7568,5708,-1311,-7451,3869,-1445,5087,-1661,322,827,-900,-916,-3974,4350,-1479,-1239,-3137,-1799,1683,2690,-1745,-465,9501,-3354,-2377,-2995,737,-4853};
    Wh[36]='{-516,-556,-1314,-4350,129,1223,5541,-522,-768,-2680,-4250,-4724,1738,-1331,-2418,-866,-2824,241,-4145,-693,-608,291,-4887,-502,-3801,-1185,422,-2155,-9296,-3034,4143,-2568,-2978,2678,-12958,-919,4218,1364,-5458,-1328,3969,-1746,239,-5253,635,-2868,-9741,377,-1341,3596,-2636,-3398,2426,-1199,2661,1159,1265,2673,-509,8583,261,-3449,-3354,3464,1611,-3647,3918,-2463,-1217,-869,651,-858,1190,2116,-5571,3269,630,-2193,2478,-2496,-394,2158,2827,2770,-574,-1055,-855,1859,1206,2097,3300,-4008,2851,-933,-5527,-1474,-2902,-2890,2023,-5390,354,-1269,-95,3088,2553,-2065,2766,1306,7954,2558,4074,4160,975,1101,117,4077,6713,3188,65,-1657,1171,-877,-4907,1933,-4848,-6308,1865,-1779,-178,-1400,-2462,1296,-2629,3371,11474,386,4660,4462,-603,3364,-707,3457,-1071,-160,-354,1766,773,4265,1673,5805,240,764,-1097,4460,-6723,2088,1145,-1910,-1051,-1185,-10722,-2203,4831,-4016,5625,-561,3974,-671,-2805,-3857,-5229,-3015,2453,1053,-252,2592,-4938,-613,3305,-7753,-2988,2910,-1662,-1021,372,-1567,-4050,3798,-2800,6665,-3964,-14,578,3842,-5097,6699,3107,2792,2230,879,-4150,2446,1076,2517,-980,-1518,2044,3156,-1477,-274,-4052,-1337,-1403,2675,-1491,-3955,275,4414,-2956,-7089,-131,-1633,-8305,-3471,-1629,351,387,-1198,-1483,970,848,-92,-1187,-1219,3654,597,-2084,-4257,-3044,-6376,-2127,3286,-7373,5009,-197,-3330,-226,-3525,-259,-1750,-7358,-4707,1058,-2766,-4902,-2011,99,368,-34,-4985,-4833,-4494,-2758,-9521,-5517,-4345,-1505,187,-3247,-953,-5800,2122,-2410,-1782,-3183,-548,-2468,-3293,-1308,-3984,4553,200,-2296,1951,140,6528,466,-3183,-3403,-4372,-98,8520,3366,-582,1776,560,-528,-2253,1224,1347,-3557,-2746,-130,-4433,2196,-5068,3427,-1656,-1940,-8559,2958,-1949,822,2893,-2656,-5815,-2773,2187,44,-6333,-5024,-3928,-4736,-3652,-825,-1301,2880,-1691,-1078,-3842,-3337,-3232,-2675,-8876,-6508,-7412,617,-6289,-1217,-3854,7451,68,-4721,6293,-285,-4387,3803,1431,364,-1947,-2993,-4641,355,-2521,-1937,791,-865,1857,-2381,-5415,-4265,-1734,397,-2690,1907,-6826,3750,3503,1020,-7924,-1788,6083,-5317,-7343,-2995,-5756,4621,-2792,-5795,-4589,4550,7016,1373,4174,-5180,-1992,643,-287,-2052,508,-323,2071,-2081,441,-1688,789,662,-4541,-1185,-4638};
    Wh[37]='{-1599,117,-391,-3774,1353,-654,-1260,1148,3220,897,722,263,467,-2312,-2209,-1433,-7011,-843,1945,2448,1173,-297,-6660,466,-341,2619,946,2442,1334,-2761,874,493,-4628,-4638,776,-2729,-797,-3828,-147,-2944,-4536,-2495,6284,1791,364,46,-6875,-1890,-853,1251,2556,-3476,3056,2832,4941,-548,-2266,369,-5175,-2663,779,888,-5825,-216,-276,1812,-1628,-5620,912,-649,3466,-999,-1632,223,-2756,3828,-3098,-57,2519,-426,-3002,-5410,-358,-5668,1326,-3012,1745,2261,-523,4147,-2451,-7065,-208,-608,4855,3676,-1856,33,-1149,-2103,591,780,2631,256,-98,-2519,3049,-1939,4548,-2388,-2805,202,-1239,-3393,3303,-3803,-785,2115,-2910,550,3264,2110,-1883,-628,2705,-932,-4030,-2241,-1541,10488,-2617,-3059,1263,-2459,3476,3095,1200,1605,-3845,-1899,-441,-2919,2475,-188,4086,-1584,549,1777,-139,2027,3066,4028,255,3283,-8022,-1446,1254,-2763,3100,-1248,-4548,-4560,2293,-4189,3696,3974,1242,1297,-2536,375,-2978,-3273,3911,856,3852,3144,1597,-3059,1311,-2153,1325,-4353,-96,-2325,3630,-2932,-2036,-4851,-1008,2421,-3781,3569,-2775,1440,2374,2445,596,-1101,2812,4201,429,2135,-993,-733,564,74,655,-2163,539,77,-2788,-3476,-2326,837,3933,-5727,1752,1516,-2548,662,-1467,3005,-2379,2198,-80,-3774,-4326,-1204,-208,242,-611,5253,-3505,1362,-3940,1067,-7299,814,-1402,-190,718,5136,-4606,3222,1185,-3059,-3852,-624,-346,-3293,-123,-3190,-572,-3098,3369,-1784,-3359,468,-3618,1151,-6406,-637,1314,-2316,-2144,-1757,-3034,4724,477,-41,-3576,-114,-1433,-283,-84,-2910,-442,-2038,-2265,-3540,-460,1511,-2685,2376,-694,5019,-1959,-464,2379,-1820,-3330,-1301,1501,1196,3024,521,2263,4431,-3027,-2348,-739,-2219,-6049,-3669,1695,-6308,847,1677,1262,122,936,-2213,2521,-5170,-2427,98,505,1411,739,-1943,-3903,-3354,-4121,-2169,1657,1228,-1555,-3969,-5488,-1166,-3493,-2919,1599,-2192,1552,-4282,-2773,2312,5439,868,-2983,2265,3281,7465,-1121,-5839,2614,-3671,-4729,370,-709,1257,14,859,416,-975,-5332,-6025,-2243,-247,-1423,1092,-3027,-3740,3332,-817,-4458,4919,-803,-9169,9853,-5576,-4548,-2932,-6748,1846,-853,3366,5498,-2075,301,1047,-1242,-2443,-6455,-1586,345,-1325,1796,-1021,2529,-3168,2646,413,4338,-4836,35,5014,-3564,-1566};
    Wh[38]='{1875,-481,2773,1027,-3027,486,-249,-3732,-2369,419,-3813,1235,1894,1466,-4584,-1103,-560,4489,-6738,2500,1034,634,2291,181,33,-2773,-125,-3010,3012,1606,1756,3183,-1246,1113,173,-2137,245,-2495,614,2218,2539,450,5625,2626,3215,2211,-4633,603,-2683,1035,-5761,2182,3183,1054,-2829,-159,3273,-190,-3925,2362,-2062,1574,-1057,-2316,12,390,4057,-5375,-833,-3247,-1080,-2785,603,1490,1627,2966,-1978,-1510,-875,-6386,2127,-8896,2110,12,-1682,-2325,1295,-808,-4187,-2238,2775,-812,1978,-5336,5483,938,-5800,936,-3972,-336,-2307,145,713,5615,-5454,4138,-453,2670,1079,1300,-781,-1500,2753,-5161,3144,5136,4631,-531,-4450,4523,3171,2160,2910,2302,-533,642,593,-3791,812,3361,-3786,-1862,-2600,1342,-2604,-898,6684,127,-3454,-1699,5395,-1495,12167,-1092,-1192,335,-2048,-1411,4460,878,-3459,5820,-1510,3107,3061,1867,2059,-2326,3605,1535,-4870,-8007,1384,-1287,-1566,2658,-2895,2895,-1100,3166,-2413,4904,-5219,-690,-964,-1141,-1005,-1798,6689,717,-4350,-6250,560,-1024,408,-1496,8100,-3874,1822,-9624,773,2056,790,2734,-897,-3078,-1429,-2531,-90,61,-2287,-1524,-2819,-2539,-2612,167,756,458,-3715,3581,-785,404,-2121,-166,1204,1634,2104,307,2220,-5048,-2019,-5102,441,-5122,-1864,-3361,-4645,587,4252,-6186,416,-1158,-4223,-2155,-2856,-6508,-522,-1540,-5014,1512,-2075,1611,-2119,-9052,-665,-1877,7192,-6787,-404,1995,-144,1607,2050,-3283,-1361,-5239,375,729,667,-115,-3818,1402,4645,-3830,-709,-1473,-61,1010,-3386,-2675,773,5249,-1955,741,-1702,-802,3110,-2683,1790,-353,-1080,-3383,1042,937,-2203,-2880,2149,-716,8,2890,-1702,-5136,-2497,3054,3320,550,-2164,-3017,1741,1308,-1234,226,5517,-626,-839,-5986,-2161,2363,-272,-1610,-631,-2302,2705,695,-5146,-468,3269,-2429,3256,-3410,-1198,369,1384,-5483,2313,896,382,-2690,-1101,1505,196,222,3457,-6469,-5019,371,-1881,-1365,1612,-1875,4326,-1928,-1100,547,-406,-2148,-2486,4196,5146,3676,-315,-6220,3645,-2844,-2288,-1384,6049,3891,-2622,-1697,-1300,4531,1556,-4758,712,-1545,1684,-4516,2919,-7602,-2073,2666,-2622,-11220,-122,377,-1293,1323,-3833,2509,1280,2739,3449,966,-2797,5751,2384,750,-2822,4296,-226,5053,4631,1877,-1171,4370,-2362,5083,4121,1915};
    Wh[39]='{2780,217,-290,-1810,-843,-810,3095,1645,-4274,2252,3767,91,-5761,928,-1567,-1006,4770,-1829,1606,755,4221,-878,1145,-3178,-1385,-1076,-285,1801,-2819,2413,1876,4213,5458,5991,995,-4213,-1518,1060,72,2778,2117,-931,-1328,-373,4599,1933,-2095,-2551,331,-531,1971,502,4855,-8471,1793,3398,3454,2261,3486,-1166,819,2015,-1450,-1904,7910,2817,1228,7290,-3659,5161,-639,2390,6523,448,5341,-386,-1898,39,-3073,-3557,-70,-76,4228,-6289,6064,-4411,2592,3637,-3640,2198,2,5029,2961,5878,1196,283,1870,-834,-2454,-443,-6489,2346,2214,-4440,-5390,-545,4079,1613,-1672,5771,2836,-1429,-8735,1932,3635,-2474,1247,-8554,792,4648,1652,-7465,-3020,-807,-110,-659,-4028,-2423,7524,-349,-9711,-4777,1054,-3874,-3173,-3576,-2408,2148,4709,-2829,-5361,1887,975,-1352,1051,-2844,-3933,-1665,-277,-1901,9116,-2012,5297,114,3425,-344,1457,-4353,-2403,-1281,-5688,310,-2061,4284,5136,2482,113,-709,4304,367,-4692,-1384,8188,-4411,-3715,2048,-2973,105,-6982,3093,-3786,15175,-903,-5483,-1065,-6220,-1075,-60,-5786,5180,3356,2873,533,5747,3571,-11220,-3288,7182,2399,794,-1771,3210,482,-1961,880,194,-1684,2459,2541,6152,8671,2773,481,-453,8686,18,-2719,966,-709,4025,936,2115,4707,5141,6059,-3156,3813,-1783,-1772,320,2397,-4150,-1461,-88,-509,-2183,-303,553,4526,2293,2092,-2553,5068,4223,56,172,851,4343,3588,-1679,2381,-300,1252,-1016,-2211,-1046,-3320,113,-897,5605,2474,2590,258,5546,2878,304,2132,-2019,-1472,1529,1284,-2553,-3708,-213,3776,-327,-4609,-44,3215,-1157,-4128,-4,1865,-601,3039,1949,43,-3400,-1834,983,-3632,7309,-650,975,-3486,11083,530,3723,2117,-5991,-158,-3093,-8056,3613,-1859,6577,-5498,1424,2446,-820,3950,3908,-1892,3188,-3862,2854,-4025,-4184,4301,5014,5351,2248,-167,562,709,-1671,122,-741,234,242,3564,-4467,-3784,481,615,2261,-7221,5581,-1398,-732,85,3876,2349,-3198,-4934,1793,-748,4440,7304,-3486,-1183,8779,-4306,3164,-3222,-3364,3630,-1668,-4135,5410,1497,-6855,1794,572,-6083,-1809,-495,-7929,512,938,-581,-6210,1492,891,-1159,472,-5415,-2268,1467,407,-4121,-6376,985,-4301,-3342,-3190,1143,-3691,-2895,-2436,-1909,-1577,9062,3249,2756,-3198,-24,2330,3647,913};
    Wh[40]='{914,4023,2384,-2541,-3142,2746,1883,6098,1859,-1303,3374,2017,799,138,6386,-513,-1429,-150,402,-2561,25,965,2402,-32,-343,-3654,701,480,-2305,-982,-1611,-3085,4880,-421,-2216,6835,206,-1119,-4672,2297,532,3896,-2277,-1596,4680,1420,1767,3730,4052,747,-2761,2486,1003,-3640,-3818,5664,180,3071,-1741,1030,1099,2966,3881,-1641,-1945,-3022,-383,5854,-2148,755,-7290,-2414,1909,5722,4213,2851,-1577,1839,-4167,2171,2707,-126,3093,4638,-1273,476,3391,-1362,5429,-1884,2254,-1267,-4147,-243,1470,-1761,-1411,-1351,707,2126,-3417,482,-3107,1539,-2856,-1021,-2114,748,-4780,455,-3613,2277,4829,4287,3483,127,-3715,-1300,-3588,-5126,-601,-1242,2705,3818,-1248,2856,1076,-1636,-568,2746,209,2303,-2412,1346,820,-1516,4025,-4282,2330,-1389,-4218,-2575,2595,-1158,3203,-2661,-1370,-935,-2980,-1805,-3454,764,4016,-2915,-687,8496,-4182,1011,-238,12773,1759,2145,1233,-3837,-2968,178,1163,4699,-1643,18,-134,1114,3090,1933,-919,-1314,-649,-3073,1778,737,-4272,-994,-1716,6235,-3830,983,449,6,-4592,-886,972,1949,1193,-397,-3583,-838,-1817,-1811,-1939,5131,1309,-5576,1041,-1081,-1959,1562,-3898,-3288,5146,-1547,-1331,3959,150,-4526,-852,602,-981,4042,5380,2514,694,-1851,-360,1194,-520,-4404,2053,-169,4594,-597,-605,-2225,-3588,591,-4028,-2309,-1210,-2609,-585,-2519,-1290,-4016,-783,-1437,-1129,240,7080,-2092,389,-48,2000,-73,-598,-1038,-2839,-1939,3400,-3195,2541,-1014,3164,207,-3027,508,-1423,-2739,1737,1333,766,-313,-1959,-4499,1181,-539,3676,-1644,-1778,1301,1117,2313,7211,623,-1940,1813,1124,827,2297,-89,2025,-2646,715,-259,871,-2243,-2731,4838,-831,1285,-845,-2568,759,-4392,10253,-88,-5117,4614,591,2524,7939,-2158,110,-2318,5849,-3876,-2585,2281,-3911,2312,1218,1853,-954,4050,-2663,457,-615,-6210,-1268,3156,-5102,-626,-4379,-2230,21,-600,853,13,1688,2656,-466,1047,3903,2548,-3994,4846,7177,-181,-9316,2407,0,-2856,-540,-1933,312,826,1055,4526,7319,-3554,603,-2397,-3745,-2619,4479,-6718,1251,1827,8276,-7504,6049,1268,-360,4018,-1506,5317,1542,2242,-4216,2022,-2648,238,8037,1209,5854,4162,2305,2717,2731,600,2027,4775,-76,2563,-3605,-379,11972,-466,1926,1861,-31,-985};
    Wh[41]='{2856,-838,-584,591,2692,1584,552,-7509,2844,2137,-2320,2235,1314,1677,1763,588,-7045,1612,-2443,-1882,1872,2653,-465,-2471,-1315,-3789,-2084,-432,-4265,-482,2288,-4155,-7578,1223,2746,-2436,-69,-1199,1958,-1950,-2373,-2792,2114,-8012,-561,3361,-1690,1942,-1892,17,119,7011,-454,-870,4365,-5195,-1383,-1280,-2785,6562,-3798,-1840,823,1483,-400,-831,1933,-172,3735,157,2810,-2381,-852,-3867,-1234,3403,476,-4843,2775,2000,1535,2687,-2076,-4379,-1868,-3911,-3002,-4345,1311,8198,1422,2512,-3181,637,1514,1478,4624,70,-2902,-2155,-6533,2462,936,-9301,11591,-378,-2058,4624,-2724,-2993,-3515,4331,9570,-3830,-134,960,-2161,220,1737,-4797,-1495,-4848,-11650,-3259,975,-3278,3479,2683,434,-1437,1214,-5234,-55,-6684,-3706,-5253,1904,-2600,-1539,1148,-623,126,2366,-723,2363,-4445,1909,-11201,-4953,2973,4604,-650,1517,-996,104,-1931,-3776,-3662,858,-12988,9311,273,-1224,1303,-1506,-397,-3156,-777,1926,4584,-2056,-2176,-4831,-6391,-6547,-191,-2565,9033,2492,-3476,8007,5615,-381,-2612,1232,-2246,3813,3073,3171,2727,1856,942,2998,-2203,-1961,-545,-147,3041,413,-1193,1777,-2727,1745,7290,741,2431,-1865,2375,-3295,4208,3146,-6323,5122,7509,4819,2739,1474,573,-3305,3579,-174,228,2429,2130,1735,2727,-256,-1315,2600,-1093,1205,874,2130,6835,-102,-3352,-1216,4692,5517,5463,-600,-2824,4990,2673,-1689,678,-7719,-5058,3215,1966,4172,1573,1551,9,-2397,-884,-4079,4692,-3518,-3107,-2556,2445,-7436,1956,-1375,3041,1704,1056,615,1691,-6093,894,-790,3886,-5776,382,-1502,3305,-3054,-716,-762,-5571,2976,3029,2634,6250,-4797,5161,877,-17,-30,8901,4372,-781,2121,3452,150,638,-8940,709,80,-1564,-1593,5839,-2050,5551,-2373,6337,-1956,-4204,-3291,-3217,2403,1441,-1759,-1861,-8959,4606,262,2988,1787,-3642,-4106,1643,1386,133,-2290,9267,4719,-2313,4633,-2998,-1241,1627,-2995,3449,3315,612,-2863,2678,-3312,2800,1740,-1298,370,197,3686,5693,-9931,-3747,2481,8989,-1667,-218,3894,-2331,-1802,2182,4538,-2159,2536,-2078,-396,1789,2253,-4902,3037,1029,1821,-232,721,99,119,9296,3679,290,-2043,-2442,-830,-3662,-3583,-2355,-3471,-2106,3190,1722,-6333,994,-2639,-867,2460,-788,-4882,-4069,-2420,-1651,-3364,930,-2266,1895};
    Wh[42]='{9575,1096,1463,-2120,-3376,3620,6357,-5239,4128,622,-215,-3688,1580,875,157,5317,-1440,-970,-4316,-2880,2274,2543,635,419,1921,5800,-173,1295,4162,-2313,1810,1844,-668,-1450,312,-1618,2242,3293,1616,-2445,-1300,190,-6752,516,-2302,1163,2064,-1233,231,-2476,811,-3215,-4782,1173,-3869,1815,2951,468,1173,1459,-1763,-319,-4931,309,3613,3808,1425,-899,66,-384,-516,1423,-3747,-2807,3876,-3554,5776,-2198,-2475,3010,-2863,2409,48,2152,266,440,-433,941,-247,5395,-374,-2395,3793,4467,-2475,-4125,-2368,-1934,1170,2229,-3630,1759,-961,6621,-3288,-496,-3615,4697,415,-4799,-3190,3212,5854,-2462,-623,1586,-3122,-3774,-1744,-721,-1904,1625,7602,2597,-3715,470,7539,2504,1828,-4719,-1649,-1148,3977,-1330,-2639,1774,9897,-1121,4394,555,4106,-882,-15263,634,-4826,333,1914,-3789,-26,2768,-2429,2084,-6376,5771,8281,-1341,-221,-1953,1101,5356,6718,-2829,414,-807,-6215,-10498,-807,1511,1174,1270,-6645,-599,-4416,-4020,1654,-1864,-1849,289,727,6445,692,-1896,-1336,1234,-3640,3803,4160,-710,-2127,8159,5419,2061,3388,-1331,86,-1466,-4221,-6230,2536,1805,-1922,-2237,-9589,851,-529,-2163,4941,-238,389,4750,789,3076,-1292,1613,4709,2059,2648,-1430,5908,-5063,535,870,4377,1589,1474,4597,3066,1485,3703,209,-2717,1756,2543,4150,3366,548,4182,-1217,6191,2509,-5820,1458,5561,-975,4055,-3491,7138,-4360,1542,720,4064,1845,3098,-2504,-6313,-4106,4882,-4494,-549,5947,-969,872,2156,-1888,3952,1026,1704,595,3471,-169,503,6118,1511,2327,4025,1181,-874,6445,3532,-1934,1524,-420,2810,1816,671,808,-1040,-1724,-1045,-1801,-1362,3564,46,2580,-3576,2006,-3564,-430,1584,5976,4077,2194,-2149,-3305,-905,1148,1583,6250,3662,3559,1113,-993,-451,2800,-2017,3674,5996,3828,2800,38,-2161,1370,1376,2341,-4670,59,-3576,-3767,1132,-3540,3376,6093,3032,3615,3935,2661,3281,-8774,-1345,6337,880,1809,-7680,5366,-2844,-2375,880,1956,-774,2073,-4108,1339,-3618,2795,-7939,172,7773,3183,1021,3862,3442,1306,6108,596,1055,381,-440,2673,1345,-3972,2012,3266,1386,4189,-1165,5991,-303,3461,-2719,2303,-1928,1170,-894,-123,-756,4560,5063,2514,4436,-4975,2587,3723,6210,-4155,3430,1690,-6723,5014,4604,6738};
    Wh[43]='{-415,1292,-1525,2315,-2136,1420,4206,2268,2641,1623,6967,-944,1684,-5053,-117,-3937,-3503,5019,4721,-447,-218,-349,-1012,-1846,2460,1021,-364,-1663,3933,-2773,-2454,-3881,5405,4443,448,7866,1188,489,3696,-462,1040,-4299,-595,1469,-878,5136,-2624,69,1915,-1776,-5053,-88,5683,-985,2001,3574,2207,-3164,5727,-630,280,8056,1090,-3146,-3369,712,1245,-1053,-2934,464,1084,149,-2313,-3742,-1209,1385,-2093,-2609,483,2687,-3242,-10673,-1056,8295,-381,-4523,-789,11933,397,-7094,1909,-3825,138,-5039,588,1712,3195,297,3571,-896,7236,6000,717,-12500,5073,-238,-6489,3708,7983,1369,5917,-6132,-3444,2281,1124,-1892,454,-3889,-1601,-2375,282,-2435,-14335,-8906,-6943,-3544,1910,-2041,4379,-4213,-1045,-2861,3200,-2316,1328,-1258,-3735,-4685,1313,3408,-440,2265,1118,1475,1123,985,3994,1998,4782,2873,802,-235,-4321,-1610,2,-6274,2983,1802,5336,-5527,2489,-2200,-840,-2301,2418,-4614,440,-2541,-4113,-7304,-496,-2875,4689,-3037,-15,3090,474,130,-1687,-1970,249,-1295,2427,-5883,1547,1209,386,343,7133,-3515,-254,1058,-5722,19,8110,-5898,205,-4943,850,2839,-1168,-249,-2092,-9277,-4084,-1228,4270,1815,-4162,-1950,-4736,1756,-972,-2922,165,1884,1174,-9194,2910,-1326,-635,5253,2218,-1674,-2183,177,-5908,-1256,1546,-3684,-4565,670,-2425,690,-7812,-1574,3269,681,3713,-2775,-8305,-3532,-2290,-46,-5698,-961,2824,-520,-5532,429,-1350,-1528,-3947,-5698,-1005,-5273,-2612,6264,-737,-2675,-4257,-5673,1680,-1314,-991,-2775,-5458,781,-3117,964,-2573,3115,1083,-3908,-2135,1236,1446,5317,4523,3032,1132,5415,-7739,-2690,879,-1575,-2531,761,-2729,1949,-1168,2249,-3342,-3012,3088,13,-3806,-3842,-3786,424,-1357,-703,-3237,-4465,-6865,-7978,3266,5019,3591,866,1951,-2432,2846,6870,-1628,-1815,8979,-1827,-1402,3986,-7080,921,5668,-642,-1067,-1478,-2136,-1467,3161,-5761,-2167,-3840,-3732,2027,5400,-1492,5683,1002,5517,-3242,-4868,-6704,-1719,-5595,-413,1658,380,-1279,-2496,471,-3642,-113,-4108,-7856,-401,1417,-2054,1175,-6621,-155,-2612,-977,-1125,-6796,-4519,3691,-1591,-4250,1030,1691,629,-3395,-2597,-9106,-943,-1722,-703,-3898,-1434,5117,144,1005,381,899,-5927,-864,-6904,-1105,1286,-2194,679,-2171,-6166,6938,2238,-3205,2749,-1506,7431,-3557};
    Wh[44]='{-3271,-6044,-59,3796,-3996,-2534,-3747,-914,-1286,-2939,-1497,121,2028,376,-2739,-693,-2614,-4396,-1983,4414,4096,-1012,5903,655,-6166,2646,779,-1905,-1635,1838,4206,1069,-3176,5317,-632,2011,-2651,5917,-1904,186,170,-931,-4775,872,1079,1564,2915,2376,-3552,-10869,-334,2260,847,-934,-1791,-946,-14,6918,1020,-2824,2817,1433,3210,234,-2651,3303,-1315,-1479,2163,584,-3950,2448,2922,2109,3864,6142,-5029,2961,1630,730,-571,3432,836,3581,-726,-567,418,461,2517,-3332,-429,-2244,7260,422,891,-3286,-5102,-5419,459,1362,2915,-5839,661,-4775,-3159,2451,-829,2802,-713,6577,1491,-8193,-15625,-885,4211,-12,4274,3981,-2531,7324,1124,-2988,943,-6030,-1855,-13828,1539,6689,8637,-6308,12275,-9819,210,-2260,3564,-4843,-4421,-4523,2440,2668,319,-2270,-443,-5722,-4372,-4296,318,-2465,7700,-5190,1232,2819,10205,-3186,7333,-28,-729,577,745,-13457,3483,3710,-2702,-1298,175,-7065,2641,2370,-557,-1322,8208,-2023,5737,-3461,6630,3261,3364,567,-4616,2009,5688,-1229,2587,-2094,2283,2988,9057,2729,6103,-7519,-338,-2279,-1492,3134,-4621,-1018,-6977,-5737,3164,-870,-3361,7700,-18,4182,-1677,197,4436,-1013,2678,-1666,2763,4826,2529,-249,4211,9057,6704,-381,7304,3596,3742,4599,7500,-6201,3828,3476,745,2514,986,4599,-457,888,3415,5102,-674,3332,2242,3288,6113,-3557,-7612,1169,-1227,3991,3486,709,3200,-4284,6293,-3056,-140,1784,1599,-99,-3,-2198,-1106,-4641,968,-2124,3298,4355,-6591,521,5859,1009,-4101,1056,836,-1999,3095,484,-607,1002,-1479,-8901,1835,8012,4914,1829,-2792,3154,-1538,-5278,3364,-1083,1409,4323,532,235,-2418,-8242,1331,5053,6542,5419,-1409,2315,2083,-1972,-1132,-1712,5532,1812,-5185,-1080,13007,-3173,1425,-1078,-3068,3327,4733,-4121,5791,-6083,655,2541,1347,-4396,-1223,3676,10556,-6308,1285,4257,3056,3757,2331,1679,-7031,-74,-670,2038,-2246,7856,6123,5883,2792,-28,-931,-1189,-3408,-881,7172,-3354,5556,1459,8090,-4145,-4226,1013,-5864,-5727,-5395,-401,1750,3967,-6596,-2382,10859,7158,-420,-3999,311,748,-601,-2275,4921,4938,5654,2658,-1079,-2008,1877,1102,5737,1073,1077,3916,2822,-745,4304,3928,-1811,551,4284,2939,1807,4924,-1843,-1765,-4589,-7163,-3229,7099,-5566,-599,9262,411};
    Wh[45]='{3789,-3420,2875,766,1806,-1651,2221,8383,7285,-543,-6376,-52,36,-625,3464,3908,-1938,-3427,-5097,581,-1123,1285,-1035,776,127,-6220,611,533,2675,-1157,-449,3681,3842,3515,-2344,-1419,-1467,653,3554,648,-4086,1553,1073,-562,7504,7236,548,6264,-804,-72,-5092,4350,4951,3784,6186,-2666,2900,-3430,2453,-6635,-365,530,-1730,-2209,-798,-3449,220,-947,160,-2437,2452,-1019,1555,-3652,-1800,2648,5883,-658,1842,-3740,-315,-259,1741,3037,3474,-53,-1868,-87,6123,938,-614,-5039,-4438,5239,-4855,654,-1056,-1193,2133,5112,-2600,-2880,-2442,-3132,2829,3154,8457,-196,204,947,-2585,-2336,4804,-2551,-2937,-3115,5864,-6240,6801,4101,-2033,-643,9882,3881,-3740,49,-2524,4250,1723,1162,-716,6206,-5087,4821,2507,1804,3500,-2700,6083,-3044,-5493,5073,189,-2230,-2507,648,-9672,7929,1397,-6752,748,-2592,1943,-3337,-4042,6572,1639,3386,-8261,-888,3652,-2707,582,4807,869,7177,1437,1139,-3427,-562,-1264,-1959,-10966,6601,-8867,-2426,3146,-1512,5620,-2322,2034,7573,4523,-7416,-638,-965,794,-2325,-8344,-2785,1009,6855,1989,6669,383,-2802,-2687,-1593,-4636,3444,-4587,-968,3999,-1898,-846,-2600,4125,-5756,5791,4233,2368,-38,106,128,-2912,-10957,3867,-5004,1059,13,-895,2543,-2744,-2457,-938,231,-181,1036,-1883,5488,-984,1109,-3796,-7685,-4084,-3371,2851,2805,2144,-3452,3503,-1970,1406,-2377,-4389,4470,-783,1412,4770,69,-2307,-4604,-2470,-3239,5859,-1096,-4565,236,5380,136,6240,3579,-3178,-200,-2587,-982,-63,3410,1489,390,1040,747,-5249,-243,697,-2602,-2116,4960,2336,105,-1779,625,-52,-5869,-5039,-1846,2612,432,2827,2609,-2631,-1987,-503,-1508,4104,6069,204,728,279,-2590,-4150,-9394,1701,1273,1145,-3276,5849,546,3134,-3393,-2812,-1054,-2347,1951,985,-6074,-8994,-3432,8818,3967,-30,695,-1107,1613,3029,-1650,1812,1213,-3088,-2302,2636,-3999,4450,-2504,3410,1839,-2614,2337,-1204,-3542,3666,-1162,-1728,292,3,-5747,-272,-1611,4174,-2476,-7656,-627,3339,3903,2861,442,1285,-2687,-73,-148,3474,-5019,-1071,-6494,-5737,-1783,4824,-5336,473,-8857,-2619,-1500,-3608,-1331,3278,-2492,74,-1800,-836,-72,2731,-3581,2231,1851,-3833,1782,4489,-1752,3986,9194,-3862,2878,-985,1275,-5834,466,487,-4804,2885,2846};
    Wh[46]='{-116,-1818,-5136,5087,-6611,-1828,61,-3500,-416,2301,3947,42,-953,-4050,1193,4130,1925,-5688,147,1617,-3986,-1569,-2512,-2242,-2344,-1667,-608,427,-1794,2464,2120,1461,579,-6772,-8500,-2189,-3698,-2169,-2922,429,-1774,-810,1480,2070,-3845,-3535,5473,-6723,4091,2116,150,-323,-10302,-432,4550,-14804,-11191,-4702,-16,-21972,2587,2854,-1374,-3337,-1895,3173,-6230,10390,-791,-4963,-1729,4465,1914,3884,-1231,1118,-2971,-4819,2322,4047,1688,-189,-7407,2741,-5078,1604,1049,2824,-2902,-811,-2863,2897,835,6137,1430,-2486,-2147,6772,3942,-1268,3859,1979,3601,-4562,-2387,414,110,4768,-1303,-7690,1431,-7651,1767,-1041,2263,-2368,-1711,4545,-2130,625,1571,8320,8383,3581,-5742,-4638,-10117,-9760,4331,289,10234,-2415,2196,-960,4445,-1,-3879,-6821,-2358,-16,6508,-824,-180,-1157,1306,-1522,1732,-2309,-8198,-6743,3364,-54,-5156,-3554,-545,6508,-1605,3110,1929,7670,-740,1571,-3054,-5112,800,-3750,-3132,-697,-1564,-3254,5839,-2076,-1535,-4416,-1506,3215,3298,-1540,183,5029,123,1601,-1496,3464,-3298,-663,1211,8793,9628,-450,-7099,2993,5751,725,-2973,8071,4787,-2829,-4111,-7377,2207,6328,4389,5537,-5258,2993,-2143,-1545,-3022,-7353,-949,1259,3933,-2780,219,-2016,5991,3723,-420,8676,-1173,426,-101,-914,6176,-5927,3395,-4067,-5048,911,1665,-2922,-1992,2514,-2158,1054,-4047,3066,6855,1888,-3825,1227,1359,1809,-2252,2291,-417,94,3381,2285,-3337,-5571,2670,-1638,3798,9541,-302,-7421,241,-4707,-580,-4396,6894,4143,-2783,-671,-4533,-6567,-4995,699,-1030,-7143,-2198,-1199,-255,-668,2314,-3596,1572,217,-6860,-1143,3256,-8417,4584,-3310,2340,-2866,-484,401,7368,5092,2360,-952,-383,-2049,3227,223,-7255,342,-2059,-765,-8120,-4675,-2746,-1174,-3715,74,-181,-1928,7592,2028,2408,-7524,3295,-1683,3911,1281,-1229,-256,-4008,2563,815,3171,1250,-361,1260,-1192,-1291,967,-4155,-704,9331,-3154,3134,5244,4987,4155,-794,-1892,-2454,-858,-1964,-5053,-2880,559,9375,2496,1602,-1010,-4182,-4611,-3237,-4011,8583,4406,2141,-2829,-91,2010,1335,-107,129,-3637,-1199,4729,-5249,2883,509,-846,-5073,3544,-7880,-5615,2568,-1932,1352,-3044,1157,7158,-932,204,10283,-5986,-4731,2736,-3503,-6669,860,1262,-870,200,-3476,144,-1489,-233,-3359,-9199,2119,1873};
    Wh[47]='{-6025,5302,-1981,4028,3371,-1656,8037,427,1095,2058,4055,-637,-678,1579,3942,1254,-426,5307,-3774,-3225,1513,2324,-2395,3666,-4282,2028,1259,1109,1333,-3859,-4953,-699,-5761,2592,4179,2110,-1347,-1020,2263,971,-244,437,-1634,2985,650,600,698,-2319,-3662,-1838,1213,2399,4589,2607,124,398,436,1844,1710,2147,44,5644,-1760,878,-1926,-1502,3840,1070,-3730,-3693,-690,2495,-2714,1632,121,-7812,-3776,444,-3740,2561,-664,2932,-4042,-3613,-1408,-1253,-3220,1320,3293,3225,-3850,-1118,-3083,-2266,-393,3227,4272,5405,-1417,26,384,3618,1685,-3952,-40,944,3562,-3879,4895,-112,3830,4887,7875,4179,-1749,900,-4987,4721,4348,1685,-1960,3168,-3793,-1210,5141,-2297,-670,-2011,-1995,-2207,3679,2724,-195,-2795,1057,-1078,9096,-2102,1916,-5434,-2919,1898,-6992,986,-268,7343,5253,-3959,-1384,1687,2695,192,4372,6708,585,-3330,-2805,377,-2438,-2917,832,5727,-517,3513,2216,314,-1435,1538,-3957,573,-1096,892,-1684,1254,-2619,1998,-1245,-1472,5112,-7104,5615,-2401,1507,-5922,5444,1860,-2900,4777,-2418,-4423,632,753,-2432,-3244,780,5395,-332,-201,-2106,2121,1173,-3879,396,-4692,-2304,-2531,-1298,-2261,4375,822,-964,-2282,-3273,-747,-1979,5898,-1718,1755,-6005,-1137,-748,3491,-102,-339,2978,-766,1464,-590,440,1842,-6386,-2213,2548,-1751,-2529,-1678,5727,-4592,-2081,1409,-3410,-1680,760,-3283,-957,-1741,891,-11103,-5180,3015,-777,4038,1729,-2364,1196,46,-3896,633,-825,-2812,5756,1928,-659,5419,4284,-1516,-1529,-1868,1468,-7031,1040,-1253,2512,-980,5419,2137,2634,-1640,1230,1759,4257,-903,-1018,5415,-4531,359,-4521,-2568,5366,-3051,872,-3056,-1728,-6635,-689,1743,-4257,5634,-9101,-5600,-4565,4050,-794,-1207,-5009,-1433,-4450,-3989,2252,-4523,-2321,-4765,3842,-2403,-353,-339,-3254,-4274,-3698,3208,-347,5161,-5278,4714,3017,2354,1962,-249,3454,-64,1759,6323,-331,789,-3725,5092,-1293,-2807,-1933,420,-2785,3908,1475,-434,-2447,-2900,-853,-4741,-4035,-2026,-2553,-824,1055,2226,-4770,-3395,-4990,-5029,828,-2333,-701,-8310,-5415,2095,-2489,3088,4353,2993,721,-385,-4230,-62,-701,362,9570,1304,4111,-2205,-569,-1992,99,-1254,5532,1525,-1194,-3068,-4294,-6474,-1578,-601,3776,-1789,-2829,-1052,-7338,917,4880,-3813,-839,-499};
    Wh[48]='{532,1602,1838,-5200,-508,596,-984,8100,-3276,723,-247,-670,3825,-3142,-3867,2198,-154,-1978,-35,3847,455,-1553,-399,-608,-1730,5229,-770,-1015,2580,-2922,1381,2661,715,-1461,1318,-1043,-4274,-1600,4057,-548,-631,-6401,2795,2612,6723,2327,-1473,4162,-247,-2717,-1817,1461,-3417,2395,-861,3845,-781,-1885,1691,7402,3427,5410,-2468,-265,-6772,805,1002,183,4797,1464,-1712,3996,1074,-2714,2590,1838,-2871,842,4538,3227,-1687,-1401,-1302,-1765,2814,-852,2502,-3691,-524,3303,1722,7172,2192,-124,4377,-532,47,-1840,60,3383,-4472,2031,-2648,-1447,2478,-190,-6064,183,-9218,1754,-2340,-1039,-8657,-181,-6787,6552,4233,-13027,-29,-488,-798,-725,9921,-2954,-1621,1568,755,-698,3857,2239,-3129,-690,-6,3520,2298,474,55,2100,3859,2218,-5424,-443,4079,2447,753,-1467,-3869,3015,-8872,142,-5458,957,-1166,-3720,1538,-4909,5493,-2191,5844,9409,-2250,-1761,3464,-3339,6352,-2512,-2310,-401,-1157,2056,996,2976,7910,3024,1512,-2912,-1040,-1525,3701,6264,2797,3684,-1245,991,5566,-78,1820,-7861,-2592,-1311,-1273,-659,4294,3164,2143,2045,-5219,1329,5688,-2524,-1246,4318,-1397,-3872,3015,-368,4343,-5454,-3608,239,3132,1557,-4565,617,1217,-6015,-1436,-6191,4411,-76,-614,-1701,5258,-7309,-3342,-1329,-144,293,-3085,474,-1038,4387,121,-783,2612,-2322,-282,1403,-765,304,-3913,-799,357,6752,1574,1347,-1734,298,2641,-364,5878,4199,-1370,2185,-5014,-9296,-320,-151,573,-2963,-58,-4729,-2675,-790,604,1253,-2500,414,2712,-439,-283,-4284,5405,2209,-1811,-3833,345,2563,-2308,1905,-4462,9326,-657,6220,1699,827,1221,5073,2319,-2312,-8549,328,-1106,5815,6347,1779,2578,-3471,394,-49,-3010,-10097,-4169,-4006,-798,-4528,-4826,3332,1541,182,-522,-1342,584,3654,-218,-1214,2274,-2368,3083,-1372,-588,2329,2331,2602,-2565,6899,-2390,-983,2239,7329,-2729,-4741,-340,-1156,2285,-4946,5039,-6337,5166,-4023,-3405,-2382,-621,-1213,-167,-1912,7919,3310,2009,-953,3803,741,-3596,-224,-20,7846,2392,3110,-4184,-4855,2145,84,484,-2064,-1705,-1412,-2937,-123,-609,-5068,3181,366,-2626,-6206,-6303,1328,-1330,-2448,1656,1779,-6718,621,-888,2437,-3376,1241,1674,1672,2199,646,-3513,728,-1170,-5532,-1215,2043,-83,4995,1979,1546};
    Wh[49]='{-2374,-1043,729,-484,1795,-838,-781,689,-1865,1262,5361,2995,2600,1668,2032,-2971,682,-383,-2651,830,1282,78,89,-499,425,5659,505,-726,50,617,5820,1936,1607,2156,-1079,664,2770,1776,1496,4138,77,-1574,3317,1582,3435,-1579,320,1130,924,-2758,-1669,-2171,-2766,-4228,2111,-2341,1970,326,1695,848,-202,-1761,1884,-707,-883,-3696,-481,1256,1069,-49,2282,1547,-302,-825,932,-256,-3261,3049,1389,2404,316,2141,-864,1354,628,-270,1198,-181,1010,428,1176,1216,4514,3149,4562,197,-142,308,1052,2656,204,-1357,-1416,-304,3142,-542,287,-379,435,-3022,-4458,-3315,4670,-669,325,161,4440,-1156,2932,-1512,-2440,-1031,-3515,825,711,6791,-2092,1339,-2585,-387,-252,-2937,-86,1932,579,-1583,-458,-3076,55,-952,1166,211,1390,1569,-3647,-3437,-327,657,-1582,-6347,-2203,-28,5200,2133,-1889,-319,2546,91,4138,996,-2238,2009,-588,1677,-703,995,-1372,1676,957,3122,201,1107,-2,545,-482,419,-555,3012,-3427,2257,-1274,-1191,1971,-1105,-276,2280,748,3049,-837,-3776,-490,251,-2873,1741,-3479,-1074,2734,-1145,781,166,-866,1372,1300,2622,5820,-372,612,-5,516,572,-514,886,31,1660,-2049,945,-1340,922,1545,3666,1083,-1437,945,1140,-2081,617,4025,-3112,4843,-1290,-3046,1418,834,585,2333,-800,1312,1468,3366,4016,-1754,1354,-3269,1381,2575,1767,126,3256,-3173,-617,-2154,-1995,-7456,4570,1661,1046,5371,4272,2148,1459,1918,4113,-3000,1043,1517,51,1983,4101,2614,-112,1285,1322,-1566,-1055,849,38,-258,1154,182,-2700,3244,2993,5000,2355,885,1374,288,7543,1343,-1685,-2661,1003,775,-451,1430,5297,657,1884,390,-1077,2384,3845,79,3793,583,1173,-563,17,3352,-2386,1883,-1193,-3186,2285,3933,485,5258,-606,1759,997,-572,527,-751,-913,-2313,3032,-3742,3825,1315,2471,-536,3032,805,-2258,3969,2939,1489,1934,1932,328,2575,-892,4858,936,-1395,-53,3212,-663,1574,-2639,578,2836,-3298,3708,-1782,2031,59,-1138,-3383,767,1508,3862,3083,4221,-3823,-1971,295,2288,2890,2042,-6259,-585,1177,2091,1010,4028,-1505,-115,-7519,-1160,4763,4216,248,1287,444,817,-235,2390,1394,-1179,-460,3461,-992,253,1195,-648,3500,-1423,-703,1273};
    Wh[50]='{-1906,-2778,-2529,-4387,1053,-2426,-2722,-639,-6098,-2330,-8300,-4743,7128,-5146,73,-9995,-4362,-8105,625,2182,-638,1352,-335,-1049,-1108,772,-153,-1237,-2351,-1503,-1038,-1816,-5561,-1619,-1555,5458,-1284,982,165,2144,3752,-1070,4023,-82,4460,-2636,-8422,4235,458,2414,3623,-4738,8652,1588,-6059,-4895,-547,3002,3208,-2229,-1702,1990,-4328,-455,-5234,-3610,585,1492,-1274,-1350,1405,4895,-167,-1795,-3447,-3513,-705,-5297,483,-2497,-4926,-305,-2751,1697,-6748,-2059,-675,-369,2558,3674,7163,1379,2797,360,684,-1666,3994,2861,-235,-4565,1416,-1516,-427,-2514,3266,-1690,160,-526,4704,-1544,7353,-784,2885,2009,-7416,884,3803,3659,573,465,2303,12558,830,4687,-4780,-11601,8920,-3918,-6743,4455,5390,-1916,-7944,2220,-3186,3901,1638,1319,2666,1885,-4194,-362,-11875,-5688,-2479,4743,617,3725,-1588,-2285,-5273,-320,1134,12783,-1679,4072,-1500,-2277,-5581,-6000,-4448,-102,-3137,-7446,1,6464,4357,4997,-2399,3359,2156,2658,2293,-2137,3937,319,2814,-5917,5268,-7734,-495,2001,-1296,2551,-1447,-602,-1361,-44,-6953,-845,967,-1958,-10361,3608,-5664,8725,2073,2416,8549,2521,778,3178,-4052,-4450,1124,3012,2829,5312,-5952,-491,-1431,-586,-4111,-264,-2883,1445,3505,2524,527,-6269,3903,6250,7319,-2003,-9702,1898,5009,-1137,-1571,6728,-4475,8886,-3491,-756,-3137,-3293,-1529,1508,975,-12763,-4333,-1802,-2614,-1057,-2817,4450,-4099,2022,-910,1209,4973,3664,2465,-4982,2910,8842,-4768,-4885,4985,7368,-3808,-3923,-673,-2348,-5292,-1796,3259,194,-2304,-365,-1242,-4616,-6440,-2741,-5126,-3527,1616,-1346,-399,-797,2883,-4843,2553,-1173,7021,8818,1623,-1907,-6181,1249,4455,4873,-533,-6865,450,4599,-299,-2939,123,-1427,-1185,-2268,-2580,-4956,-6215,-600,-2548,-3579,-5341,-6201,2010,-2824,-2008,-6469,2381,-6259,-14638,-8413,-1839,-2194,-684,567,3083,309,-5283,3063,5390,3156,-4499,2766,-12226,-4294,-271,-1079,-1468,-9965,-2844,2467,-238,-3964,1817,4802,1507,3259,991,-1807,1712,733,-7294,2230,1710,1798,2321,3701,-4199,-147,-7128,-9497,11298,-3713,-583,-7465,2303,-6752,-5214,2502,3139,-416,1772,-2401,3547,4335,1572,-5429,1236,-7827,-4409,-7270,-1058,-423,6547,-7075,-1354,-1351,4345,-7968,-2714,5937,-3232,3688,-283,-1828,-2883,541,-3591,812,985,-1550,3029,-1761};
    Wh[51]='{4392,114,108,858,111,395,239,-3786,2315,3686,2651,328,1815,1423,29,-1796,8735,-5502,987,2971,254,547,3134,2073,-184,5458,-1099,859,394,3493,-3500,-734,5356,-2373,4216,-1898,-1012,-616,-3320,3215,794,-6596,1660,3181,-299,-1650,2187,-4436,2734,-1315,-6250,-2617,918,-3764,-4018,619,-661,1408,-1553,3388,1831,3901,-121,-147,2364,-2575,3208,-1760,1960,3254,-4768,-814,7924,-6225,-550,-187,-6928,-637,-3173,1546,-2255,-4763,2044,-9116,1896,-3024,250,-1107,-2088,79,1339,-705,4453,2998,-6723,3830,-914,3586,-928,3178,-5541,771,2164,1187,3764,631,-2065,10527,5180,-2347,4443,2763,2990,-5073,5146,5678,4492,7890,154,-2697,-897,-3405,1292,-924,1776,-3359,7714,2780,-3676,-6362,-3208,-560,-2866,1459,2128,-921,8256,3337,11406,-1274,-1828,709,16162,4504,-2391,3952,-1705,-9672,3740,4948,-1625,-4465,-339,134,5327,-3264,1435,1704,8168,-375,3972,1363,456,2434,-2399,-6533,-217,6977,-763,-555,-6210,5136,15175,-2919,-4306,-327,-878,-3549,2758,-3188,-9204,3125,2442,1536,-6650,3410,3447,3857,-5576,-3942,1348,-2695,-795,3623,-3449,8432,-3562,-354,3046,3742,90,72,-1206,1751,-3134,-925,3334,-4860,-7895,1212,2073,3852,4873,1282,3132,775,2780,-1500,-1756,-358,546,-3173,1840,12,-4843,-385,5253,2183,-1082,1407,2802,1433,-4255,2812,101,-4101,227,186,4929,3051,-2337,4116,5532,-1345,-2239,1347,3107,-8886,-1042,1944,-224,5185,2709,25,-1090,1939,3383,8027,-2019,-1812,-2854,-831,-385,-6093,330,-1425,5478,-564,-604,-156,180,2030,-1362,-5747,-1422,-447,-545,-3698,2993,-3122,1851,4482,4367,-177,-305,6914,-1773,-265,-5126,-2211,1425,5483,-1192,-256,5947,-5449,-904,-2008,6621,405,1646,-3139,5327,-8125,-2692,-1193,-5083,5473,1813,-1413,924,3723,-3125,-6708,-4941,3095,2651,1538,-3852,-3625,7836,446,2340,-1940,-3603,6196,-1635,2231,-3781,3027,1693,3244,-972,545,1287,-9013,-560,3217,-2961,-362,2303,3833,-351,-3754,-78,5839,-14589,2924,-5415,2124,2517,-131,4765,1783,2396,4245,5297,-8666,-886,8232,-1301,3813,-704,1889,2354,3171,1596,-5224,-1038,-4790,4565,4191,12041,-7675,-596,4157,5703,1308,1079,933,-1146,2634,-2932,-1739,1783,-2548,3527,-3020,-2934,1932,-194,-1979,-2333,5742,1331,-196,626,-3728,2905,-1798};
    Wh[52]='{2208,-1138,-121,-7099,-1254,-810,-685,828,-1516,-2388,-123,-1776,-561,-2954,-1920,-6562,-8,-5078,-1811,-17,2192,155,3527,-2216,-926,417,-1374,-3808,-3134,-569,-789,-372,-2326,-1574,-755,-2158,396,-1416,-2215,-3649,-1604,-3305,1367,3325,3508,-5415,-805,4528,-3852,5708,1247,-1357,122,641,3276,2932,1763,4807,-6381,1322,-2113,-3605,-2344,-1010,620,1773,1147,-3977,3239,-1318,6,-6000,-3879,2191,-5498,-2958,-3850,-1937,1585,1319,1527,592,2078,-6625,-1828,-1380,3630,-1392,3247,4206,-1893,1549,1376,-2587,1739,1334,-1687,-6,1011,4082,2288,-2152,-4848,2105,-2357,758,-1519,-1459,-3193,3007,313,5878,-3173,3962,2944,776,894,-376,-2919,793,35,5693,-1124,4152,-2387,1473,-38,445,-823,5961,-4699,-882,-1408,4453,6079,115,-1206,580,3291,-1518,-2463,3234,-2136,2966,1920,-5913,-4511,7622,-623,4323,1417,5786,-11279,-7045,-5253,235,4206,117,3728,-2452,-3310,2257,1118,171,-1733,5170,-3820,-3112,-1031,-370,-5156,-2907,1218,-2178,68,-3776,-96,-167,-6655,-1290,1418,1101,-2437,317,1252,538,-5756,-5063,-2382,5317,112,2404,-25,2264,-1540,1502,-520,-599,6494,3837,-889,-1953,2844,2214,-745,3220,1927,3251,3928,0,3703,-682,-7299,-2441,557,2258,-1212,957,764,1002,2006,-10,-1309,-3093,-3645,-1516,453,592,668,-610,1772,-1181,-2546,739,-573,900,-2746,848,1151,4421,-1807,-1854,4650,3251,-491,141,-759,3051,42,895,-2905,3103,-265,3483,-5424,3002,1138,2536,2147,-1809,866,211,-894,3647,2937,2027,-983,-417,2352,1925,-3437,3288,-3691,-1628,-1680,986,1938,6054,-5791,-1518,-1813,-48,938,2457,2214,-2856,1948,-2580,1558,761,-5249,1390,6694,2186,1317,-572,3647,473,-2469,3288,-6206,1746,-2893,2243,3063,-1267,644,-2232,437,654,-158,-647,5292,-2181,-1739,-184,2120,1123,-606,-857,1678,414,600,-3559,-2575,-3222,-1923,233,3884,-7495,-2076,-224,-440,-2924,3532,-3256,-3354,-1013,495,-209,4580,-841,2604,2993,1992,2587,1304,995,302,-3820,4484,-4858,-1900,253,-474,-1279,2666,-7641,-2094,-2028,-4711,2349,722,2697,-2687,-7065,-1434,1558,2495,-5156,2209,-1770,2275,628,-3503,1004,-2014,1828,-339,1032,-1619,2047,1734,-136,-52,1888,1915,3281,-1553,175,-1011,-1126,1094,131,-1754,7192,-681,1195,-3156,861};
    Wh[53]='{-3225,-412,-139,939,2181,-1264,-1662,-1688,575,-203,-3784,-1734,-789,3923,3513,1665,-127,-2597,-2529,-1757,-1983,2556,722,4357,-885,6289,310,2459,-5322,-1028,-1823,-561,3444,268,-892,-2233,598,172,3200,1756,-4921,-2880,-3962,1771,1948,-1990,-1676,3596,2257,2397,-1666,1638,2315,5449,7670,2631,1876,-3005,4826,-3156,-2427,4792,4758,-5346,-1990,-1051,-1972,675,-1628,443,5546,4235,-2546,-2419,-1826,-3874,4025,860,-167,3999,2153,2490,2868,-2186,2800,-4719,1767,-1328,-927,169,-5458,5195,-6865,1248,2568,4208,-779,415,769,-2327,8623,4016,-2800,-249,5273,2032,3078,1102,3186,-2347,-3862,-6982,-1535,2181,-3320,-1401,-360,455,8579,3093,-3159,460,-3537,-5473,2648,8237,-8315,2178,1368,-87,-224,-3210,-875,-2301,-2966,701,-3735,1777,2792,87,-1948,4255,7172,-1376,4860,2336,-1380,6835,-2014,1409,63,-1510,428,-7211,-1183,3251,-2272,-3525,-875,3908,-2368,4807,-1409,6860,-7646,-92,186,1833,2036,-2379,1701,-954,-7412,-1560,-3869,2788,-2243,7690,-1112,-4003,-525,4506,3881,-2397,-114,-2619,2668,545,-10400,-903,-1877,1075,-1036,-6752,-2304,339,2359,877,-4147,-115,-3308,-760,3134,8354,2717,-99,-4218,2302,-899,-2951,1710,-5312,-1564,-178,-4628,-5141,578,-1667,-3732,-954,-992,7338,-859,-2012,121,1849,857,-1589,-4931,-3930,2988,-103,1527,869,-5454,435,3845,-385,-1671,-1628,3925,-4992,-2529,-4616,-4658,2585,-3332,-439,-1840,1178,-2176,-4968,245,2003,-610,2595,2277,-1434,345,1341,1011,-4604,-2573,-3879,-23,1084,-2425,-1572,-3852,3737,244,6005,-223,-333,389,-2915,-2651,-1006,107,1582,-4616,1402,-6899,1209,-1795,-2406,788,-3864,51,-1043,3493,989,-652,-460,-2658,-673,-2418,-124,162,-3754,-4313,-514,3076,1136,1172,3032,-1284,-6352,859,-1633,-2055,4257,-3066,-2824,3728,4223,-313,-2177,1712,6528,6313,1961,-5698,1065,-1361,4301,-828,4777,-1380,67,-342,-2888,-263,-747,-718,1528,1616,4450,1796,1910,3706,-401,1187,-2198,-5517,-466,-643,-4165,2220,-1177,-1242,3901,-2578,5175,4599,-3786,-1500,2932,-3073,684,745,-3779,-3513,4604,-11679,6669,4206,-793,-774,6435,578,-1276,-2963,5107,-1372,-4177,-601,-3417,263,-127,1100,-2373,2496,-1531,406,-2042,3764,-3024,2211,3991,-2590,360,1386,-651,-3913,-1131,5395,-6030,871,256};
    Wh[54]='{4870,6557,1606,5068,3947,-745,1873,2971,4062,3554,-578,1394,3671,2418,3173,-2441,733,3730,2758,3149,2042,2012,1040,2592,593,-236,2340,-622,-278,6088,6010,1108,4101,4824,-6323,2607,4506,2519,-1264,1579,7182,452,10351,-307,8315,5214,2724,1706,2113,-4245,781,2983,-2141,3249,1219,4631,4396,491,3020,5092,2629,350,-289,4252,-7832,1940,4538,5288,714,-549,503,578,4853,2714,4431,9707,9160,4306,416,2851,1667,6733,6254,1821,1268,957,-2188,2436,-7998,-1539,1387,-520,2116,916,1640,4064,-2536,6967,1884,2509,-6645,3295,2235,14511,423,3730,139,-3691,1105,347,2854,-3945,2937,-822,-3088,7255,7875,11083,1490,2110,-4123,-913,2415,3100,1118,-1628,1479,4143,-2082,-7167,2434,2509,-1436,1823,-501,2844,3374,-5415,1729,260,-1328,-2912,6381,-4357,4511,-690,-464,-1859,-3698,2462,2225,3564,-2849,-5068,2844,6547,6206,2707,1795,11875,8183,1066,-890,-6440,2985,2399,1917,2553,-100,-3259,1258,4980,-808,-2058,-3151,-3054,2746,-4135,2253,-725,-1730,321,-7963,-504,-8383,563,5317,-4323,93,-6313,5864,-3305,-3110,-2546,-3298,-9946,-6308,267,-5898,1430,-723,-1237,-2702,-1573,-1514,-2187,4572,-276,6293,4333,-2614,3215,6220,118,-952,-577,180,7583,3911,993,1392,513,1994,1220,1766,1879,708,2054,-1357,2266,3552,-2465,2181,701,-6806,-5937,3999,128,-310,-4750,762,-2507,-4841,5776,-2961,1264,1263,-4501,4753,-795,483,-2459,3933,5556,5058,-463,-888,-3515,6230,3254,3334,5361,-2893,1057,-2670,-3234,4553,3962,-1552,-236,2749,208,1737,3903,4028,-1831,-1855,-2191,930,2231,1510,1529,2385,-1102,-974,6865,2082,1021,5566,-4157,6801,-50,-724,1238,-1381,-5278,4174,-7792,-899,3999,7993,-7714,2836,2878,2242,4348,5419,4421,3564,4675,-37,5273,-1624,5268,575,-1505,-5717,7592,1577,5898,4699,-664,6640,-1219,13,-2763,-145,2573,-785,4228,4641,1301,-1578,3359,-1937,231,1391,1044,2954,-9257,3789,-4335,2924,890,5688,-5551,-1036,4389,1752,2617,-2418,523,-2480,1788,-1602,70,7412,-3203,2425,-3620,8422,386,364,-2261,1517,7514,7451,-809,-115,-6386,7236,2536,-192,-4865,3242,-1914,-472,-1242,2646,3935,4699,1103,3403,-2846,3916,-4858,4946,3559,1746,315,21,3337,4206,-3574,1745,-7290,870,2407,214,1816};
    Wh[55]='{3784,5961,3996,-4636,-2473,-3364,1242,371,-5668,3200,-1262,-1768,1109,-1464,3710,741,-58,-3037,1575,180,965,159,2495,3090,-5498,3127,-1227,-2683,-7319,-1621,3708,502,-2553,4375,-16660,2225,-10761,6010,3073,-105,9414,4704,2687,546,-797,-3967,-5112,-2241,145,2457,-2044,1243,251,6328,-1088,-4104,20,2614,-744,-12041,7705,5361,3684,-4553,-6357,-875,345,-4733,2995,906,-3977,737,2230,-897,2875,809,4658,5825,-2297,-2003,3269,4975,4765,1896,-154,-2687,940,1480,-441,4230,1605,-635,-468,6357,1411,-797,1738,-1680,1822,1944,-3383,4870,-2917,-7797,-4111,3676,5288,2604,-4509,516,-2663,3708,-2139,2060,-1269,-3215,938,-3632,-6083,-1467,-3342,4895,-1867,-602,-7207,2526,-616,-2778,-2900,3645,632,-402,5927,3593,15634,-3957,-6772,6474,-1669,3630,-6201,-2277,-1893,1317,-3256,-4060,-457,3789,5810,3195,-4645,2407,2624,560,-6562,938,1505,-281,2636,11923,-3437,-543,-184,-4985,-1916,11162,6811,-2111,206,-1527,-2443,1130,952,1045,1149,1612,4812,-1195,-3200,-924,-5,-3881,-3190,3349,-2807,51,1169,1085,-2404,1179,-6518,-2198,-3115,-1287,3505,3684,-428,1019,890,6279,1157,-1308,-1092,-2415,-4101,-2006,1162,-264,1687,-5654,-1749,4377,-5156,2524,-2775,2127,1684,4328,-562,3132,321,1141,-1434,1457,-2489,2071,2631,-7529,1539,1606,-2929,-1125,1152,-2009,4738,-4631,-4504,-1386,1126,-4355,-3242,3469,603,5224,-1634,-424,5249,1993,-1683,2761,4829,655,-2008,-2746,345,-8276,1232,-3789,-680,5302,-452,-3415,-4323,6386,265,-333,-5322,2478,2092,220,2229,-6821,2318,-2114,-1175,-3552,-2575,-178,-1146,-2612,2322,-1748,-5576,-11806,1233,4548,-443,-7919,-2841,4599,7172,-3928,3669,7719,-2871,1842,4013,843,354,-700,-1121,1468,7319,143,-3544,-1383,1549,-3562,-1483,1612,3559,2257,2110,-1993,-1149,-8891,2617,7265,4311,-2783,3217,-2536,3200,-1550,-2054,4711,2583,2360,-255,-813,-3686,880,-4565,-2976,983,-7519,-7387,8344,4978,-722,9658,-1864,5234,961,366,-1606,-457,-4179,-4489,287,3386,-728,648,-3564,5478,-6665,4208,-4304,2780,-8095,545,-579,2410,-4753,-3002,-8339,4809,393,-501,1683,-6162,-1212,-2266,4204,1993,466,3391,-1590,-1370,5053,303,-8720,2617,512,781,31,809,1242,-10576,6381,6342,-882,280,-545,2724,3356,-565,481,-3723,-2624};
    Wh[56]='{-112,1662,-1029,-3530,-2127,-764,1037,-5024,-138,878,-8637,-1243,-5083,-2032,3039,-2331,2863,3283,-848,1407,1867,2279,82,-2902,-3745,1341,-2514,-1711,343,-1062,-59,-3649,1007,4240,939,-3925,-1085,-1148,-327,-398,5668,75,636,-2349,-941,2770,1181,-3918,-803,-148,6464,-2277,-4582,-3903,-2534,439,-3166,-2297,999,7202,225,-2751,1756,-3588,-2369,-2529,-2225,-344,879,403,2451,-4011,412,4167,-413,3664,-5439,138,7036,1001,-1834,8349,4355,-3662,-575,1693,-1004,-1056,-96,4082,2465,-3889,-5087,-4328,-2291,4594,-2653,-1649,-2324,1250,1932,-3164,-526,-949,2824,14,-1176,-11640,1685,-797,183,13867,-7890,791,-45,-2164,-1706,2438,246,-3911,2963,-4912,5327,5893,-2500,-5576,-3125,-4084,6459,-59,4494,-4489,5625,-245,440,-4580,1322,3439,2700,2119,2827,-3969,-792,-1799,952,527,-3327,-626,1297,-2629,1636,5039,-4416,3105,0,-405,1446,697,-1182,2165,2946,-4228,-5576,-898,4716,3835,-1330,370,-5737,2076,-1990,-4389,-1586,4289,-847,989,736,3630,-971,-44,-2551,-913,-3596,1467,3330,-2714,1618,7465,4724,2059,6699,-1422,1994,3964,3640,-4965,-2041,-2866,-2335,2490,-1481,829,-1574,-3776,-4924,-660,162,113,-4697,-93,4724,1431,-3366,5410,-1788,146,-1962,2790,1211,425,763,-4323,-5864,2202,836,1003,-2749,-2001,-617,2729,-2008,967,106,-4238,2490,1082,-2440,-255,1619,6552,-531,3701,-3085,3603,-383,690,-210,-375,101,1189,-1872,-841,173,883,3903,1993,-2064,-4128,1412,-2556,-8081,-139,1584,2098,-463,-67,-4846,1163,2078,-785,-666,693,-2534,3662,-795,-1739,-2253,295,-1237,-1370,2086,-7807,1403,5498,-2724,-459,3635,225,-783,1111,-2371,2065,1921,3061,4880,-2690,1632,1341,-1178,-794,548,4348,-2095,3244,1274,-3129,-3994,-3410,-9316,2181,-1817,-1633,-558,-1787,-1483,-1484,4890,3449,-5478,887,-327,-2912,-3581,-3295,-3400,-7348,-3334,-2070,3898,-1214,-1702,2261,486,272,-177,2463,-2727,-3937,-3889,981,-2746,-1875,-220,3684,245,729,474,2998,-3867,-2543,2253,133,-4858,-2183,309,-6557,-806,-6596,7700,-1211,-3872,1447,-369,-4096,875,-3027,-1098,-5405,-1951,-6777,-410,-4924,-2244,3723,-1545,-1503,-1251,-121,139,-4548,786,2700,1636,-5161,2727,2849,947,1111,-2,-1274,4020,2741,6718,-408,952,-2209,860,5126,-1286,3325};
    Wh[57]='{1638,5859,466,-5527,590,-2553,-11728,4699,-2263,-855,2341,337,3852,2551,-4479,1352,-1647,-2592,-1580,360,-2058,182,1907,-1768,-121,2413,1865,472,-394,-6796,-4689,-5659,10,2451,-3254,4191,2355,475,-3378,3789,-508,3459,-4079,5214,3771,-32,-3117,-2644,-4697,1225,-6918,2069,529,-945,-2447,-2939,-712,4570,-1375,2412,-3183,-7231,314,-1375,7573,-2358,-2006,1239,-1042,-1057,-951,126,-2164,-3022,-246,-1772,-4357,3610,599,537,1560,-5532,5844,-938,141,1286,2937,-1463,-98,-1350,1833,3786,2233,-484,-1499,1644,153,-164,619,1875,-1501,-707,2121,4057,-2268,2507,-3132,-14414,-380,-2403,1560,-596,-3359,-4147,-5576,-2253,-7797,-11718,357,-1878,-3366,-152,1673,-607,4379,2731,-1680,2702,1390,31406,-3076,309,-3239,2839,-354,2585,-1488,-236,-3188,5297,-6093,8359,-7539,-1557,-849,4306,-1734,-4306,-172,925,-2966,2644,-1215,-3676,-739,-5175,-9375,1907,-5322,7182,-6801,2117,88,-209,-2932,185,2023,-3034,4323,-3339,4541,1710,1766,-2053,-1877,-4284,-4118,-6796,-11,-155,292,7993,-608,442,-2060,-4853,3806,-5502,2243,-4445,2795,-1779,989,-1033,-4475,3593,4560,5727,5263,-947,-491,3725,-298,-696,-625,675,-5693,-8735,-1622,-178,8007,4187,-242,-1721,4729,-2325,-3588,-5507,-1746,1739,-856,-1403,-644,3723,899,3632,397,80,511,3049,2534,-5869,1100,775,3530,-4775,2514,593,-3762,-3828,-1339,-8408,-2878,1212,-3273,-661,-2756,3149,-174,-359,-3679,-3112,-2687,312,4895,-1710,-4509,-470,-222,4062,5224,1029,3110,648,389,-1823,63,1256,-1480,2651,9443,4108,960,-1580,-1150,8916,4162,-1296,-1558,103,4587,-619,-2109,-10595,-1213,-4819,-1369,1335,-1837,2900,9814,-14140,-182,-3962,-7797,6752,-118,-2276,-1806,-4567,3823,11542,161,-540,642,1139,-3239,-1866,-5864,1706,-1287,1091,2990,-6777,-1646,-805,-7939,-2658,6308,2178,3623,-3937,-3991,-34,270,-8,-5058,3132,-1437,-1071,2248,-3056,1364,87,1752,-6142,1550,8344,5864,-3161,108,836,-2484,-3574,6533,396,-1510,-5629,4458,-2856,-2392,-6108,3125,68,7211,-3259,-4685,16875,9770,3027,-4772,-3662,-1776,3178,7387,4440,4501,-603,1290,4882,-736,-4899,334,1174,-3862,-3334,-7895,-3410,-3242,-7758,2626,-2546,-6591,-4462,3376,3171,3464,7602,-6337,879,10683,-13359,7626,-5185,-4519,10410,3913,-2636,-4392,-140};
    Wh[58]='{5073,869,-814,2622,548,-1136,4038,-358,-4135,4047,-1087,2939,-1368,-298,4274,-85,-241,4890,3530,-1888,-1322,1915,-605,4731,-371,3801,-1444,170,2761,4375,5424,2242,-1041,4904,4145,3054,2458,2761,-1100,2145,3005,443,3742,-625,638,512,5678,1029,-1613,1342,-1904,-1522,-2753,-2185,-8212,-4934,1436,-8867,3571,2800,-655,1121,-44,-809,-5263,561,-869,2165,4169,-961,-2058,4448,-409,2106,-309,4135,3342,1475,1846,158,1477,6430,-2399,3378,1678,-1184,-865,-2437,-2658,2425,4038,-175,2119,-1436,7397,3725,373,111,2307,2851,-5834,-1840,1378,3171,-4326,1835,5117,5859,1872,983,3920,858,-624,2406,2310,-2805,1518,8754,6015,-5927,-2751,-8691,-1556,8051,377,2359,2021,223,-3000,-8041,4020,3405,-2321,-3188,-6157,4165,5068,-5966,3635,1450,850,-2819,6494,-2447,-540,-1365,-2648,2144,4902,1833,-1888,5097,3708,-5009,2946,-6015,2880,1220,-2000,-8803,762,4487,-585,-3554,-2003,-2792,-671,2573,4704,1696,-2402,-2509,-3208,3898,-2961,2442,1916,5014,-5664,2083,2905,128,30,2683,-5063,-3010,696,3847,1250,-1165,-3229,-2941,661,4592,516,5297,-3117,-2900,506,-3869,-1429,4990,-4631,1790,4099,607,-1796,5957,472,1701,-3784,2602,9150,-4294,4467,294,-1075,-415,513,1595,4394,6025,2861,-2462,161,1221,3271,1890,1726,-2683,-394,-1673,8085,-736,5571,-577,-344,-1679,6723,473,2841,-369,3159,-974,-972,392,-1065,-7026,1788,421,3261,952,-1374,-891,-1932,3354,5283,-1572,4660,-4001,-2612,7158,5195,3684,-1773,-462,-153,5761,-364,-2658,-2141,-5322,1855,-88,-1574,-7260,2309,6596,-1052,457,-3876,-609,4570,4287,-2307,-1540,2442,2519,377,-2019,3500,7866,3825,-1281,1136,3898,1123,-700,5703,-1832,1468,-6362,-1557,2873,2081,-651,5761,-705,1309,-700,-2038,1866,3598,8007,4462,2873,3066,-1822,-1453,6113,3417,5063,1717,-1540,3852,3139,11650,3681,3950,4821,-994,6704,2756,-1699,-2578,4489,3090,2961,1667,3774,33,773,549,2276,3271,-3457,-5151,2849,14218,4904,-2883,2253,-2105,-2541,-1750,586,7553,-1647,60,173,8237,7456,5327,1405,-4626,-3625,-321,2054,513,1219,-1315,2214,-987,6005,391,4858,5522,634,-1934,5097,2651,-1039,-338,2966,-10,4724,3994,-210,663,4333,-1156,3188,-7670,-435,1795,-7055,-1502,251,4665,1948};
    Wh[59]='{-3686,3286,-1697,-3012,58,-1000,2261,-1268,2341,-3596,-5878,-3425,-2390,5136,-845,-1210,-9721,157,-221,-784,65,1265,1956,1126,-6704,1113,-2296,445,-906,-2097,2602,-781,-2792,-4560,-13935,-4250,-7080,5209,-1082,479,7612,-2255,1633,-2619,1579,966,8374,-1351,-3544,718,-2626,-8320,2021,4133,1718,9267,2502,4704,1745,-10146,5327,-112,3359,-6904,-6079,123,-520,646,-275,-3977,3354,1291,-3671,1475,247,-825,1257,381,5800,-9687,-1905,3564,24,-579,3808,-4562,263,-543,287,-1203,-2332,-7426,-366,4875,-572,-2113,-504,-3510,1342,-1219,1898,444,6914,1146,-1826,-14,4125,2663,5498,-1264,34,-3605,-2089,1226,307,-10908,-3527,4777,1839,-12558,2844,905,1685,2065,-11796,-4174,8881,-1175,3154,-619,1141,-4431,3151,2751,16904,-1026,-19208,5336,323,-253,-1311,930,6201,-132,1022,-1218,-1284,-1813,1799,84,-1770,-48,1596,314,-3859,5048,2834,-1092,4519,-15722,-5786,-1850,-4191,-1900,-5488,8671,1612,370,-6708,-2435,2839,641,191,2817,3701,95,468,4401,573,-257,-1937,-7539,1744,1527,-2426,794,2751,-50,193,5205,-4074,-488,-1651,-1390,834,2988,2170,-3234,-198,-2125,-4655,4152,-2344,2485,3642,1408,1848,-877,-2080,-4401,-5053,1173,-348,515,1516,-5429,-1326,3562,-3029,-1468,-1304,-1590,-2108,7656,4372,-1668,158,138,-2044,-2783,-2091,-5019,-1403,-5229,3610,-1206,-8388,-1295,3149,2504,-7924,-1610,-470,4309,-3710,-396,821,-3083,-3142,-1904,-6586,-2539,1589,-2113,-3601,-7812,3959,3906,-671,1865,-1671,-5659,2124,-313,-5541,-5615,-2280,6650,-2397,-255,-7026,2360,-3620,-3405,-8413,-2490,-3366,-2218,-4138,-2236,5346,-7802,-5771,-670,-718,-915,-451,-1228,-2479,2724,5820,129,-3662,6079,3537,7827,60,-1330,3076,-371,-1582,-3059,3771,1840,2237,-6293,-432,-5917,829,813,-3437,-2646,1334,-721,381,-744,-415,1451,-3061,-3457,5346,-3693,3808,4187,102,2614,1209,-3132,-37,362,3742,-7636,-8315,-13681,8457,-4218,7421,7851,-4294,5712,-1451,346,267,314,-2578,-1340,-7568,5527,7075,-2014,-1084,-6772,755,-3425,5922,4243,5722,-2624,-55,-3286,-651,4794,-6728,-1434,-5815,-9394,1578,8857,4482,681,-1743,-938,-1530,-1545,9018,363,3999,-2111,-611,-2741,2318,-10449,3681,-5732,2910,2958,1711,2517,6420,-1783,6347,-7182,758,-1289,30,-2978,2812,-194,3071,-2880};
    Wh[60]='{1503,2810,3540,1229,473,-1613,5205,4501,2318,2604,3964,3535,-3459,534,1879,5097,1049,1234,3281,2266,1500,-4499,-6958,-185,5551,4797,4733,1027,2678,4428,1839,-761,7661,3271,3820,50,3254,-4194,2326,-711,6264,414,2705,-1782,-4194,1905,749,1312,5561,-9580,-712,4421,-290,4736,6557,-3652,797,3564,6152,-145,17246,2073,3432,3730,10341,3925,1730,144,235,1594,4941,-3605,1457,1602,4458,3850,1687,-5209,-2932,-5473,1413,2045,341,-2519,7475,-1357,3994,3452,724,8090,3461,6230,4255,668,-880,-2144,2810,-2609,1442,3708,-3430,1907,-3623,-2514,-643,-14,-8007,1614,-9501,3464,3613,2814,5781,-958,1674,2434,-4965,15214,-4030,-1361,-258,-2005,10214,34,3762,2053,-4218,-3618,1372,4167,9291,1654,1539,-617,1667,-2193,-4853,-1992,-6162,3801,792,-2398,8115,-3498,-2371,-4074,-2049,-9985,-6250,6455,1501,2556,1259,-2988,5771,4279,-6235,603,-4445,10410,-3085,3322,2338,-2482,2812,-1375,15,-4082,-1882,1685,10546,343,5976,-869,-1130,-6459,-4287,-8725,-7133,267,-1878,-2614,-131,3037,1195,2961,-3393,4406,-1854,1900,5014,2229,-2924,-27,-283,-1589,-2402,-1953,-2563,1901,5859,294,1320,2109,2636,151,321,1044,7080,171,4968,6459,2359,2037,-995,3740,5239,3923,4011,3989,-107,-4006,3635,4421,3374,6782,1552,-706,6328,4453,6909,7021,-349,6333,7988,3483,274,648,-2006,-1795,2485,-1420,2399,4294,3659,4504,592,4616,-1021,7597,2303,2800,3784,180,9467,-3569,408,-2005,7124,-2939,5664,9331,8520,-589,-1828,3305,4113,4135,415,3581,6718,1513,1850,2374,3049,942,-1431,3850,7363,4899,1947,-4360,-1442,444,1862,3945,-132,-3603,-634,-180,853,3488,7626,2397,1348,625,859,-3059,-2253,-5771,764,6064,5830,558,2022,1655,1978,2810,4379,4196,2653,6591,4758,2159,6474,4499,1361,3945,3056,-2775,7412,-734,1839,-1286,1843,2626,1140,-4108,3322,4062,4572,2316,1898,5585,-7348,-3261,653,-164,8227,1923,2336,2423,5224,-1676,1492,-3322,2841,5278,733,3500,2614,8896,564,960,-1966,-5444,5097,8603,6596,4916,15361,6943,5629,1297,4470,7504,6513,2951,3032,6689,4741,-3752,941,9326,5141,7280,-336,5141,-7109,-169,8857,-9248,5419,5107,149,2673,4489,5312,-1776,-1211,2012,4621,8193,-3208,-5639,192,2126,-13,2058,3894};
    Wh[61]='{-5117,-176,4321,-1307,2056,3681,1080,3618,-699,3095,202,-397,-942,1654,-4248,505,-3051,-900,1015,-3188,2824,1195,-3117,2556,-9,6870,9414,741,6704,5771,2558,-5014,3920,1524,3110,-2939,-274,-121,1837,1752,88,-3063,1984,2244,-139,-1022,-915,-3728,3469,-404,-213,5834,-4824,-1733,-1977,-2812,153,1795,3249,8994,2376,1398,1209,2279,2199,6264,-3403,-2758,-527,-4877,5478,4465,-919,5527,-255,102,3125,-1365,-1728,-4343,714,7768,3107,4543,516,1513,-57,-2125,4370,5869,-2600,-5317,-690,-1141,-1170,170,-1505,3281,1805,4074,-2196,-162,-6127,-1050,4680,-2156,-3356,2907,-2646,3217,-680,3715,2010,-1276,3913,-247,2609,1511,-1401,-3625,521,6708,-1646,5439,4506,-8925,894,-3615,6420,-653,8383,2858,-5419,4304,673,-4372,-758,1887,3493,4057,5927,2636,-1658,1760,1233,4851,3498,946,8359,-4143,0,-2446,6518,4689,1889,-1257,-2978,986,1231,-3557,119,-4870,-3039,4277,2971,-1676,232,772,638,-805,4282,-209,-10947,209,6870,-1215,2431,2258,-3566,4304,1832,-10888,-1188,-399,-385,-392,2553,-1226,-1517,242,-1898,40,-1777,-21,-711,2053,90,-4865,1932,-405,2797,3142,689,8164,2343,555,2060,1384,4099,-1721,5161,4523,-2259,2216,6513,3635,2113,-816,4777,-42,-1014,5385,4091,1374,31,6284,-4011,-360,4086,-157,5590,2934,-4924,1630,3234,5795,2824,936,6953,1706,-2126,2059,180,4392,459,34,-1740,-3193,2888,2089,4785,949,2985,1693,-436,2775,574,1547,2832,-2629,1231,977,-1276,2770,-2939,-2639,2176,2656,709,-1850,2169,-5454,3500,5517,6210,-2264,3015,-1162,543,-974,651,-3129,2968,4428,4333,1123,480,321,-1071,3435,-2241,11376,-2071,1728,396,2983,-2233,3039,-1081,-2602,-1128,-158,2069,2147,-344,5083,-1397,3574,2998,2187,2648,-52,-2073,1325,-4116,-861,-434,1435,-2854,-7626,2622,7441,-3337,-3488,3972,6376,2653,1119,4748,1986,-1166,-1545,2362,1237,-4819,4809,-308,-3664,2316,15,-3417,4799,-193,3903,3146,-1611,3186,-121,14238,586,626,8330,-1853,2653,-3537,-1439,255,7485,8735,255,2529,6210,-279,2878,4667,-1322,2087,-3725,326,-2519,6728,-1469,-5385,11894,-895,1644,1370,5727,1795,-4863,3754,5073,-363,-1007,311,4274,746,1787,1030,-1105,1141,-773,4099,-5200,7031,843,-2944,529,-3635,1369};
    Wh[62]='{4331,-600,3085,-458,1258,-980,887,1541,4289,-1032,681,845,-650,1166,-2812,-2666,-897,1160,1070,-2194,-3645,-1124,1387,-2208,1121,-3671,57,643,324,-1914,-672,2215,-2998,-3706,2741,5229,834,566,-4829,-1660,-3869,297,1024,1250,82,1199,-1457,9926,-2583,-1459,2509,-3674,-4104,-4958,217,-6142,2937,-422,2983,7846,6582,3835,996,3393,4182,1402,637,-1312,-1212,276,6933,-1020,-100,-2110,553,1933,-2604,2624,-942,484,436,-2255,1767,-870,1707,951,-2946,-2805,4184,-276,-2449,7075,4736,-808,-2521,5722,456,-1962,1917,749,-709,2697,289,-8325,916,753,-4675,1730,897,6132,5620,8618,-3554,-1750,1242,4672,2386,461,-2434,-6250,-761,-3442,1320,-2834,1680,911,2294,942,53,-3637,-6884,-763,-1132,-493,1586,1218,-3266,-3488,-2500,-173,-3515,3093,3151,-2534,-2130,-4389,-870,-7163,2135,-8374,-2017,726,-5390,1456,-3791,-3034,-2424,-1336,-164,14531,-1138,-4323,-925,2602,3159,2775,3107,2856,484,-393,-1273,3244,943,2269,-116,-3596,2075,-5473,631,4526,625,4135,3425,-1033,-220,512,2113,-7138,6513,-922,757,-5600,-5712,5024,-616,-3645,-3945,4912,1045,5268,802,2275,206,2229,4362,-232,-3615,5917,-783,3256,1431,3146,-1810,3332,-400,-2946,-1353,-2548,1413,699,1194,-1114,-4575,3498,-1096,6933,2004,2773,1214,-989,5703,-1111,947,-1950,-284,1229,1495,261,-4096,-2138,-3103,-112,337,-2094,-1726,-3703,735,-6137,4443,-629,-2414,101,4162,-231,2077,1746,1341,1304,-322,812,-2641,-408,-1923,-4233,-825,1351,1284,1137,2421,-1582,631,-2214,4448,315,2592,-3935,-922,-4118,3381,-578,3720,268,-1065,-5019,-269,-7714,129,3017,-2145,-4897,-2807,-28710,-1674,-7602,5351,374,-6567,756,9238,-7622,2583,1558,886,1124,1475,-1752,5351,-3298,-470,938,4179,3862,-4111,-1333,-39,-4062,5937,7749,1268,-109,-491,1097,2344,-5083,-615,-2890,-1872,645,-1090,1771,6450,-902,-1005,4904,-1815,-5332,4172,-154,2749,2504,-3791,970,-1756,-3669,566,4343,2493,1705,-3291,-2031,3793,3581,1972,1533,760,4047,177,-736,867,135,5336,4020,-4528,843,181,938,-874,2120,-1024,4428,1326,-7456,-851,-4111,-7661,-364,5864,2180,-2322,10283,495,-212,-5087,-1442,-3708,2365,1905,3557,7216,94,4531,-871,7187,5146,8696,3344,-3173,7700,3955,-814};
    Wh[63]='{-4086,4523,-2303,2131,4084,-577,3283,-2553,1733,-2121,3740,-3061,1828,-2988,3164,-5703,4313,-596,384,-18,-2795,2543,-284,4057,6479,8530,2044,2169,-1798,2010,-2329,-3208,9931,-389,-255,-377,-1245,1774,4365,2047,-2534,-792,-7963,297,-209,1856,2197,5922,-702,2169,7543,-393,1488,-5351,-681,3654,4074,-1494,3242,6962,-7749,1568,1474,12763,8769,-884,1680,2824,-2037,2156,859,2719,-2069,1896,3005,402,211,2369,-1741,-1846,3151,2150,-795,-957,-1840,2315,-672,2583,7,-2719,171,-808,664,-889,1163,1362,-46,3405,-555,-2678,13496,-1414,2087,2673,-3503,-828,-4370,213,2739,-4389,-1627,-4321,6528,193,-657,2142,-725,6367,4975,-4414,-1806,1008,520,1200,5375,4707,-82,-2344,8623,458,3681,-2045,-2080,5585,-1755,8168,6586,-63,-1330,-260,-1052,1385,1217,-7329,747,6591,-4377,-4133,2736,-470,2438,-3840,1155,8623,-11269,-5102,3049,2534,-3217,-4389,-4121,-1694,25,-685,-6230,-5224,95,5073,173,1810,5034,2507,314,1982,-3508,-4418,232,-2425,1072,-75,-648,-1920,-2524,-2470,-6992,1320,-4528,8090,-16171,-1367,1580,-803,-5229,4182,-434,2675,3579,-2109,-1342,4020,-1214,-4648,2436,595,8583,-855,5839,985,3701,1053,-3017,1270,10019,-895,1839,-772,-1632,761,-579,-5390,-4672,-2431,-2390,-3129,-7387,3852,-3735,-504,6708,396,-2399,3876,-1988,-406,-2089,2773,-1859,-3171,-2250,4243,-313,3891,3483,2091,-425,5214,1154,-1060,1782,-3662,-1575,-2312,-1823,-5966,4082,2352,4145,-5375,2568,1923,-101,-1160,-1455,447,761,625,4313,2091,-1610,227,-5039,1473,4042,-755,1866,-3520,5439,-1519,-7324,4545,2912,31,-446,-938,2963,-4079,2000,-5131,-3293,-1876,5927,6801,-937,1652,2622,2636,2617,138,643,-1428,4755,632,3525,-4812,1148,6904,5351,-3129,3061,-2880,-2224,-1235,-2418,2739,3608,-1523,-1174,-7041,6962,-3422,4873,-2229,-3020,558,-2253,1660,495,2247,-539,-4411,-2888,-2037,1511,827,257,3200,-144,-3303,-2517,-102,-4838,-1861,-1466,3164,-6083,-1453,2045,4997,1248,-5961,2442,2656,-1741,-3281,-2128,1667,8510,1075,5283,-6044,-7861,1102,2476,8750,-5976,5473,3127,-1956,3693,-324,-1428,-888,2008,2663,-1871,-722,-4079,-476,-2851,1151,4694,-3881,8046,-2736,-957,-754,2644,1082,311,-1343,-2362,1207,3784,-7622,-1126,-2178,1322,-2189,930,-4921};
    Wh[64]='{-1295,-3400,3623,-1960,355,277,944,7182,-1093,-3115,-8554,1396,2082,605,-103,-4284,3852,1585,2316,2418,368,-3986,2622,460,-2539,-6430,1019,-5000,-3071,3071,4853,-3164,-9453,-25,114,-441,-3845,76,-11,929,-909,-2053,2873,-588,-2568,-905,2746,837,-2250,2066,1685,-1163,880,2402,582,-1710,-2059,4113,1057,1572,1202,1322,2404,-2717,-4528,2139,-5283,1276,4501,-1479,4965,-892,7182,-955,714,-2751,-2563,-4692,3095,-1700,2893,7700,-6083,3554,493,2249,-2336,841,5683,2091,1583,687,5122,-3178,-2493,-4523,562,-574,2646,7514,4655,166,-328,-4094,1206,769,1904,7236,-7949,5649,4567,-410,-10087,-1828,1809,240,903,-4865,-3559,5927,-2614,-6127,-4204,-2861,-12216,-4316,97,3942,254,-1882,212,-4060,285,2602,2602,229,-3593,-1101,-1458,-889,-8374,5854,-11181,-702,4729,1172,1616,-767,10595,-1196,-2022,5185,-4050,-9550,5317,1855,-3715,3476,-611,-8178,404,-277,2268,-7656,-5307,12744,7075,-819,-282,-2410,3767,-2219,606,-3432,473,911,-2259,3093,5952,-3601,693,2861,3869,-4130,4777,942,4851,-4880,3645,1884,-3544,2885,-9926,2268,-550,-5380,-1823,3205,1119,1047,-775,2236,4167,-5722,-1069,1218,124,-5175,-52,-2541,-2354,-1021,-11953,-1492,-622,-4313,-2254,-6254,3649,1993,426,2331,-1184,104,427,-2431,-5014,-1810,-6279,497,-2088,-7373,-12685,-2308,-1221,-354,3330,-1025,-3181,-3178,-1105,-4528,-979,224,-6093,133,789,-1821,1329,3574,-4472,1993,-5537,-2232,-383,-7988,-4128,-5336,-2727,5424,-672,-3281,2824,6318,1939,-3371,-4497,4116,1722,-5751,-2731,-2279,-1190,-2827,-6699,3125,-6293,-4306,-3007,-3791,-3339,2612,-5156,1372,-4291,281,-6655,2636,-1335,-2670,673,-5693,2927,-554,1788,-2504,-1988,-99,-355,-6567,732,-9340,3293,-1567,-1975,3579,8305,-4455,-5991,616,-3947,-853,-3647,-6503,7539,-3991,7504,-2115,6328,-1695,-4360,733,10478,-3967,6923,700,-586,-4489,5249,8261,437,-200,-2320,-3913,-639,458,-410,6293,4548,-8750,1719,495,2719,-5932,21,-698,5722,-9355,13427,820,2827,-4128,479,-375,4841,-3183,-3601,-5776,-1450,2038,5136,2064,-2412,-5981,-323,-4582,-2692,-2392,-2426,6347,4040,-6030,-706,-2702,594,-6723,-2531,-6118,-1682,2205,520,-3583,3876,382,-3010,3869,-3085,1975,3403,5581,2497,-5932,-1096,9428,-4570,13476,4265,809,-1232,1148};
    Wh[65]='{-583,4846,889,-4108,3791,621,-5937,-2335,-1368,601,-6064,-4401,-841,2592,958,2349,2266,609,-1605,-2917,1220,-388,-4770,1680,-2116,-4592,-2663,3254,-2651,-496,-1799,-2866,2268,-1614,-2797,875,522,-1138,-383,-167,-1936,-1082,7788,1429,-7768,3662,-6875,-855,-248,631,2751,-1855,-3110,1879,-4138,2507,1378,1571,-1033,5268,635,-675,-3442,-1485,5297,-2458,-1446,1989,1923,-706,-1636,-4069,-588,145,-1268,-883,-1076,4680,-1903,-299,-697,326,-5341,1658,-2795,2281,-1994,-1953,2827,-1486,-561,1925,1065,-2451,-975,-1053,-2961,3205,1192,4296,3664,-3796,2290,-5483,-325,1074,2683,7485,-13037,3161,3442,-994,3129,-1530,3271,3422,-1263,-7353,3708,-2729,-166,-519,-877,-999,1759,-1921,3747,-640,-880,-6064,2426,-1342,-2780,-7504,897,-6777,-6250,-425,-3811,-1396,2026,-148,1555,2717,-277,-5087,-2873,-973,-1468,-3715,-4943,-3200,-6806,-4355,-2780,-7021,-2006,1464,-2724,5356,3723,1067,1550,4868,-1770,479,3083,110,878,-791,10107,8100,-4355,-818,-7426,-5839,3061,-409,1988,303,925,-6611,6855,-726,-1206,3786,-1701,-97,-5288,-196,895,-1429,952,-1722,1687,-4011,-2917,-2507,-1699,-5180,-33,5087,-717,-2095,304,-968,-1641,2426,6987,-2163,4165,1135,2269,-1005,-1500,-3410,-2856,-3310,-466,-484,466,3300,3212,6059,319,-1612,821,-858,364,2958,-3586,-3349,1021,408,1644,1061,-199,894,-5107,-3181,659,-3559,4516,-5053,3784,-198,957,1495,1575,4084,2746,-2496,-4028,-470,-4675,5244,2479,-1622,-467,-9677,-4152,3032,6611,519,1130,-894,-628,-7333,3029,-308,1182,-589,2519,818,-1165,-4609,594,809,1805,1074,1155,-5703,1467,-8627,-633,2817,-2707,-85,7,3530,3374,-1104,1286,-4697,-3942,-3208,-256,-1368,5751,-2006,-1883,-1259,-2437,-1391,1347,176,-2371,-1085,2387,925,-1983,-1724,125,-4794,-6503,1437,120,-2626,572,1901,-2788,2641,1256,5273,-330,-5917,-2302,-1170,-138,-3017,-23,-70,-9033,4006,-3952,6831,-860,340,-2127,-4299,-5327,17,2761,-3464,-7392,7758,946,-1082,-787,-1109,2225,-3381,-2937,-180,-1733,10029,4670,3259,-508,-3520,-696,-460,159,1824,-1021,-361,-131,99,2315,-364,4587,-326,4184,-4343,-1181,-3090,-438,1436,-5532,3703,-31,-4792,455,-4963,-2222,2907,-1115,-4931,-2700,1077,991,-5185,148,-6503,-5351,2060,-2790,-1427,2607,1395};
    Wh[66]='{-1252,6699,4204,-485,1043,-1062,-5727,-4377,-2678,2293,2644,-531,-1889,3344,5126,-8520,5932,2153,2893,-1263,-647,850,-597,1217,-1994,2607,525,-1529,-1901,-458,2145,1561,1188,-108,-1901,-1002,-4538,2451,-2335,6879,-1901,2197,-1993,2288,-863,-1776,-5014,-1574,1105,-1008,-8681,266,-703,1102,636,-3759,2470,-101,-1295,1779,-913,-2347,2033,-68,-1227,-411,-5625,6391,-419,-19,-2692,-840,1987,-78,3120,527,-14,3435,774,-3164,1719,2910,-3559,3032,-1073,-1121,209,1022,-5844,-1328,2814,2849,-1408,3854,-1806,-3500,605,-2192,3212,-2493,-2785,2910,373,6318,-4804,3862,1900,1724,-1001,732,2072,431,-1995,-1602,5092,519,-4121,-3071,-1840,-3041,-2548,2032,-188,4536,-919,4746,-278,-3537,-5039,-6054,811,-2498,1303,-1440,-3872,-628,-6215,3269,-4543,-2398,-3835,2331,-5253,3901,2790,-7031,437,-4875,1591,-1082,-8823,-20,-3347,4345,-1430,-2500,-3581,504,-376,6738,-2426,-3959,-1953,-892,5888,-1431,2481,2178,-121,-1149,130,10009,687,-403,3073,637,764,-258,1284,2281,-3789,-1986,7207,3752,-5107,1708,-518,238,8300,-3986,-1732,-89,5371,-1054,466,767,474,1250,-185,-392,-52,2541,-1034,3913,2167,294,-15,2048,-1654,544,646,897,1513,3762,-2648,828,-870,-4331,89,-4758,-1353,3085,1892,5756,-3212,-5712,3637,543,-8535,3405,4589,3999,5664,396,9228,1008,-459,2182,1143,-5361,-1002,-7099,3684,2841,-3249,-14,1668,-4592,-1842,3413,997,-1462,-1981,-4042,1324,1821,-1392,2551,-5629,-410,1411,1407,4375,4624,4501,-1733,1702,-747,-1280,-795,-2004,-2423,1386,2467,-842,-3708,236,1112,1020,816,3422,4533,-720,-6342,394,2810,-784,4809,2578,-358,-1155,-1813,1169,1174,-3955,7924,-23,281,4233,-5771,-15,-26,2424,3200,-206,866,3522,-4672,838,6831,1771,6723,-1954,-575,-1457,-4011,-1461,1989,3388,-1466,-4250,4384,2644,3884,-4409,-1972,6367,-764,-6499,-3471,2380,-2773,3286,3156,2076,1345,-1374,3645,3991,-942,-5273,357,-975,-702,-6562,4279,-9125,-3229,7543,-1873,-3649,1279,-1047,-3547,6162,3344,-960,7026,-3322,1920,-1150,3276,-2507,-1981,-3144,2844,661,-721,-2937,8793,697,5942,1536,-1606,3464,2420,-963,2001,341,251,4145,-2985,-2861,-38,3383,1741,-132,4729,-4819,529,-1538,-2949,2292,-1389,-249,1669,-5141,-3530,-1078,-1827};
    Wh[67]='{4428,10537,-676,-3161,615,24,-3142,2768,6157,929,4082,8120,5058,-2617,5678,9907,3688,15000,7319,-336,4052,-207,-3037,828,1419,8461,1916,3125,-1525,1733,-1307,-8232,1806,833,-1999,743,1802,5,-3498,78,3510,5190,10800,2556,4077,3410,-769,2413,-637,3920,-171,-4235,5068,-387,10869,4479,-2055,2578,-5971,10507,-3557,3261,-1177,2189,6254,-971,-1035,-4462,-2021,-592,-1226,3488,3332,451,3354,-2551,-770,7553,5522,1362,-1827,4365,1503,4472,-3872,-6899,-711,-2792,5869,3249,7797,-4226,4060,-3188,-6557,48,379,2219,2597,-913,522,4797,-1730,11035,-2330,-2202,-1007,5332,-3708,-1950,-566,-19677,2237,1721,-920,-5854,6376,-2512,-2222,4116,-1013,-2136,8901,6103,1802,2152,5141,5234,-6499,6972,-3542,2624,276,7011,10273,9306,9296,1030,-3212,2546,-3317,-1468,-3251,-995,910,-3637,2303,-4189,1168,767,1345,1302,3112,-2619,-865,-3342,5136,-4130,-232,17910,7880,-1108,548,-3610,3120,249,1434,108,1110,-113,2492,-224,2094,2685,-393,-1448,-920,-1437,-445,4812,3520,8837,-5439,-1040,-3461,-2130,7045,-6508,-13935,-2219,-131,-3212,-3085,8818,3793,10722,1413,2255,4804,1205,-1953,2100,-3547,-8745,2973,-1445,-623,-5039,2376,3696,-165,-867,6030,-8769,2597,-5078,-3420,1646,-2218,-3769,2290,1364,-3400,-357,-4306,4931,-2167,-1376,2609,1342,2401,2362,-733,-1730,-6679,-2379,-6748,5463,-5502,3193,-1445,946,-6245,7578,-4003,-647,-7138,-3168,-255,-3635,-5590,-2846,-237,-1267,1003,-2687,-1966,-2373,-798,-8500,-2181,-5673,9423,-1081,-6713,-6865,-3422,6909,1333,-3588,-2626,2768,-986,1194,-2465,1608,3349,-3522,-356,-4357,4416,-3322,-1630,3078,-3564,2180,1195,-4265,-2705,372,-9863,3864,4990,-969,-2658,1898,-4353,-5161,7041,-202,-310,2445,-4460,-1774,1868,2366,1258,265,2976,3684,-2558,7382,-5312,-603,2836,4741,-6381,-1303,-2030,-4836,4064,-6459,1002,-5117,-4160,-431,3808,-3181,531,-2661,2325,-6977,691,-5092,5463,5283,2680,1157,-339,-4140,-5502,-1589,-684,3896,1258,-1501,5727,2875,7739,509,-7387,-4113,2607,-5834,-2191,868,6630,-3884,3923,-2293,2922,3635,350,-824,3095,2551,-5151,-189,-5234,-13574,-3266,3972,-2541,-2139,-7749,-3403,-1569,6147,4604,2988,7514,4089,-2758,1140,6093,-6098,-2203,1331,9414,-3093,-2352,-7050,3203,-2770,270,-2763,-2963,8339,323,-2187};
    Wh[68]='{-2016,5141,1257,-3120,3161,-93,2282,-5239,-661,5180,4987,178,-6069,3066,5517,4780,7778,2592,640,-1115,-957,1291,1105,691,2609,-6362,-2673,1032,-4345,4287,-40,1673,2727,974,-5097,-2072,-2531,606,1099,852,237,5253,-7900,5307,-3024,-1697,242,2902,-1469,-1146,-7299,1386,-124,10185,-5766,-407,-161,-457,689,2253,-2438,886,3364,2692,2563,-2038,-159,1655,-1127,-1273,-5810,3127,-1525,6831,6582,-4599,3251,-3476,-444,-25,-112,1738,-3496,6816,1701,245,106,325,-1491,-3906,258,5053,-154,-2476,2036,-3105,-1340,5092,2261,5673,5678,-3132,-2448,-4406,-1508,3393,4089,3547,-896,607,5864,2656,592,1920,4599,-2639,-2239,-4169,4580,-1145,-2629,-4016,1276,3469,4416,985,3188,-653,-3017,-8618,-2384,3684,1237,880,-6757,1630,358,-3566,-1910,-2418,-2314,722,2038,-4440,-1663,1135,-635,2293,-2066,-5454,-3569,123,-10673,1785,-684,-1850,-7792,4233,3676,8569,-2126,-4291,6889,1122,2020,311,-630,5253,2917,-116,5151,6240,-6547,3815,-67,1708,4360,-6479,8105,-2653,-4870,-13662,-1162,-3015,-739,3457,-728,561,-1188,-3273,3422,3205,2443,-4074,-2364,6059,-2293,1949,-3232,2486,3479,-3547,-1145,-243,382,-1530,681,-2683,983,6411,-4873,7250,3044,-445,1484,-83,-847,995,2609,-3811,2329,2868,-2187,6845,2653,5893,4562,184,3188,-18,7177,-7680,-3666,-909,2316,3415,2788,-466,2084,238,-1107,-7856,2568,920,1661,-3225,4460,2401,-3068,5781,-1,-1822,-2619,3037,809,-1348,5229,-91,-215,-2425,9506,1666,314,527,-926,-4392,705,4929,1408,1473,6484,121,5600,1939,4958,1040,2467,5727,-2644,2156,6767,-3127,-1628,-283,-1859,-1286,2067,1427,7539,1041,4616,7558,978,-7373,-1217,-4113,4160,-16,3164,-1182,-737,3732,3688,-972,-23,5737,2985,811,-1007,5039,-4592,4711,-1425,4055,3432,1713,-188,-1113,2788,-2443,8203,6855,26,3596,2360,1722,6318,-1862,-1593,-6782,8540,5844,3862,4721,-3205,6342,-1365,900,108,-4558,-3730,-4855,-37,-1712,-8710,-233,-2629,-220,6166,405,-4699,-3964,1306,4538,-1322,-7314,5751,13134,7270,-204,-1658,2700,3703,-1143,-9775,1762,5927,-3559,-3098,5068,1586,-5224,6367,4377,4726,-1284,3271,-495,2211,-2272,2702,-1029,301,-578,-1685,-1231,1044,-3913,-610,-1661,-3642,5468,4899,-7358,7670,-1286,-1684,1643,4306,-782};
    Wh[69]='{105,-4511,-866,-2175,-1981,3417,-1649,-1097,3552,-4438,-2354,-723,743,-1661,1154,698,-3835,1334,355,-1282,2868,-1752,-2352,1120,-365,-891,-3354,2810,6132,2968,-493,1625,-5000,26,2102,1134,-3759,-1984,-196,-4394,481,-3649,8925,-3332,2469,-1166,2770,4291,-102,1210,5219,-1485,-3271,-4023,3945,-5800,-2902,-2324,406,3,3439,36,-1036,4091,1976,3007,1658,8471,-2030,1265,1613,85,-2458,437,-2519,631,1646,-1883,-4448,2053,-4096,3447,1602,-7226,3073,-2442,102,1267,-1920,2058,-1975,2172,-2482,-2602,3317,2612,0,-2868,-5600,2990,-4291,258,-296,-7358,4611,-1678,-5976,-2036,-4045,-5981,-519,413,5029,733,-4116,-4338,5419,8725,-308,7558,1722,-3862,-1953,-4643,-1645,3461,-5522,1297,10039,1890,-3095,4235,2990,3461,-4096,3464,5766,992,1380,78,-1849,2907,-4270,-1303,-2058,-4130,8774,-965,6547,-1921,6435,-5063,2012,-3630,3918,1722,1807,-5278,-7329,1068,5410,6870,239,2122,-4565,-875,-2023,2274,-3317,1622,-968,-8569,-4748,-2949,898,-1564,1702,7158,-3173,752,558,12480,-7011,5849,7124,-2763,-3854,2883,-4204,7080,-1791,3195,-6796,2199,1334,1527,3479,-4042,-3608,-937,2491,4714,411,44,-3041,-141,-501,-3342,-1239,-1052,-772,-2714,3110,-1212,3684,758,-502,-1519,-2775,5068,2097,-778,712,-286,-9755,-1909,-177,600,-1341,-1209,2409,3593,8198,-991,-11093,-1791,-1571,-610,-854,-1445,79,823,3881,1234,-983,-274,-155,282,374,-4758,3828,5737,-1806,-455,1287,1055,-3557,-3784,742,-5478,-2219,2626,303,-1817,1186,3989,-686,-3305,505,286,-2509,-5854,-415,-23,1895,-1520,-4184,3937,-858,-3073,-5185,-757,-568,2252,2255,-8466,2414,-5097,213,466,-4323,3110,23,-605,5712,-4719,-2766,2678,2031,1087,-3588,4003,-8540,-930,-5083,2258,1115,568,2663,-1838,2319,-6523,4794,5629,7050,2388,-1077,-832,-7270,1868,1989,-749,1816,837,-3330,-5703,-253,1052,5947,6069,-3073,-1674,-92,348,-6743,8232,-698,-3251,-1326,-659,610,-2763,-235,-5297,3811,-4934,2144,3295,-4084,332,8940,5576,-2016,1691,-4760,6743,-4291,-4370,-3503,1253,-2824,-1459,1278,-1102,5078,5322,-6972,-2457,-3315,579,3276,-3210,-5761,759,-4106,-2546,3247,-1429,2495,-2352,-4929,4926,-1062,2797,-1481,-4587,-3679,-3166,2502,-1706,-3071,8583,-3215,1351,-1860,-4360,435,778,220,4990};
    Wh[70]='{-166,2390,-647,2220,1374,2142,3808,2685,4724,3476,292,-1357,-7021,-1192,4611,949,2919,2341,8681,11699,2951,-1645,1452,1416,3969,-1818,1660,-1055,5444,1635,3061,-3728,1307,-1669,1,-2573,-1098,318,-4240,-102,-354,319,-6030,4770,-2087,1831,13,-2042,8344,-3823,-3813,-601,6909,5405,-309,444,-4338,6889,4580,849,11435,6601,-5166,2661,-1137,2536,1174,-2470,3083,-5224,-520,-3762,-44,1300,4287,-3144,2551,-1453,1060,-842,1000,337,-2277,-2753,-1774,-3261,3823,430,209,-1116,6298,895,-3666,-836,-1005,3229,946,-1071,-563,-1102,64,2675,-2241,1190,3002,-2095,3654,-3437,-7871,1292,-2590,-3869,-2546,1811,1735,616,-191,3237,-12890,2337,-1778,2073,3444,-1202,1021,5893,3596,-3146,1864,-5576,7353,665,98,-786,628,1784,-1988,-5,838,-548,2166,-2298,-6054,-50,1319,-3979,-2277,-9399,-385,3366,3679,-1590,-7797,775,12832,-2995,-912,1593,-8408,2944,12783,1881,-674,818,-1488,2580,-3969,-2115,1496,-778,-4946,778,3005,3115,2524,349,712,971,4230,-179,2824,1491,-2988,-2163,4289,2846,-3173,4704,4934,5952,118,2077,720,-2707,-473,-6518,-2022,-3647,-4562,1556,3586,102,1823,7031,5937,-1442,-5434,-1318,71,7792,4960,2025,8134,7968,2932,-2143,963,3039,2115,2102,-1015,2152,2403,7714,4633,4492,-1749,-2498,1756,4116,2117,1817,-2819,-1434,3239,4667,387,-2119,856,3027,3815,-3037,9682,-4670,3269,6967,-2210,-573,3935,-63,-3061,2447,3845,-437,4582,81,-3293,-6376,5488,8422,625,1909,-6401,2719,-612,4667,3088,1756,1488,-2094,1656,-1176,1723,1994,-1069,1724,54,-116,3085,2624,-3886,1168,432,-320,-583,-3281,-1525,-3229,318,-4223,-3232,4157,-2727,2487,3195,3398,-124,-2529,-2973,3703,4592,0,-438,-1868,3942,5161,6127,-611,7622,4616,-4709,2281,3693,7319,1478,3142,-2102,-963,2456,-4260,-2561,3803,-570,2211,7153,12753,9599,-5039,-1629,-1333,980,-258,2749,3508,-257,4130,493,2846,1193,701,728,1936,-5517,-350,-917,1093,1992,6196,1798,-178,-2352,5830,510,3942,-7631,-4812,404,-1790,546,786,13076,1140,785,1795,1708,6782,2485,-81,-251,-1178,3154,2175,-851,714,7504,5361,-2546,1588,1433,-1197,-1708,-3674,-310,7211,-3666,-1667,977,-1284,-5180,-591,-9047,5917,9057,-681,-1942,-7407,-3762,-2871,2768,905};
    Wh[71]='{-363,-1726,-3273,4760,-168,-1087,2653,-5747,2022,1372,3774,-248,5620,8486,-1640,2736,1447,-2242,105,1222,-5830,153,3852,709,-1583,-5195,2158,877,5258,3732,-3139,-1939,5185,2227,-479,-1746,4028,2546,5375,-1854,236,1113,-1204,4138,-1547,-3923,4169,-2912,-2491,-1995,2580,-3063,1638,-5415,-4091,5278,-3984,-1536,-2322,-3103,-680,-1201,5717,-1304,-602,2183,-3120,-5571,891,-4824,-5517,5122,1162,-2680,-150,-3349,1877,1244,-8779,-329,207,-721,-179,100,328,362,941,688,967,-1787,-3315,-3754,-3752,3210,-2426,-3952,-1800,-3828,2325,-2658,2031,-795,6176,11679,236,643,538,465,-2541,3615,-274,1826,-6782,-1314,5346,-2476,-4606,4731,-197,2575,-5126,-5019,-3576,-1470,2000,7778,4580,-2153,-416,-462,1217,-1,-521,-7202,2875,3427,-3623,-3854,3139,1763,-1350,1378,254,-2105,178,1262,1672,-1007,-1549,1192,-2434,2000,-3513,-2895,1128,-6298,-5844,1324,4355,-5629,-1978,-253,3403,7636,89,6718,5336,-3867,728,-562,-7089,-606,5727,820,-798,969,1372,-6948,-1859,298,9165,-6406,1760,-3615,-2358,5649,1568,31,-1589,-1701,94,767,5732,-1129,1932,4887,-1116,-195,-6245,3327,-997,-1058,-3601,-4401,8608,-1440,-1093,5068,6469,2807,1723,2792,-1986,-2578,-276,5961,1221,-579,-2700,-1694,618,2181,-6923,-2016,4221,1282,459,-2795,3051,5180,-853,738,4401,860,3020,7680,5766,-183,-1323,368,2178,-6835,4091,1871,-61,-1668,-1889,-5024,630,1342,629,-689,1171,-1043,1343,671,146,133,-4245,-2031,2197,2012,1039,1535,5742,-3410,-1315,1750,-565,-960,3479,1326,-1782,561,-3132,422,1530,963,2856,336,2573,1091,1697,2099,-4492,5590,5024,-1859,-1811,4804,8725,-5615,1923,-9677,-9746,22,1061,645,2966,5039,1824,-5683,-1304,6547,434,-1456,3117,-3125,-1947,-1431,-6992,-79,-3459,-1677,-3120,-5292,3015,29,5239,2342,-2298,4042,1424,-3549,7412,1567,2226,-2053,2724,1948,5239,-1079,-3618,5112,-3518,733,-1358,6694,-4545,-208,-1171,3376,715,-3186,-7661,3044,-1083,-2822,-3342,-3061,642,-3005,2337,-2839,1909,-1970,2587,56,-2286,-2331,-866,-3312,1933,2166,-1967,4616,8696,-996,-945,-4052,1222,-6928,10166,-8662,7089,1318,1466,104,-2597,4555,-3293,2617,5576,902,830,3225,2871,2631,-2233,7080,-3579,-7802,-301,6245,3322,6357,1719,-2215,1128,3891};
    Wh[72]='{993,-1529,-1395,683,5786,206,-1035,-2226,-306,-783,-5932,-2459,135,-4621,-6220,-5673,433,2734,363,2066,-775,-2432,-689,-1459,5346,445,92,-351,314,-580,820,-1328,1805,-1812,1571,-4135,4123,-2381,-934,-4641,-664,-1517,1745,-5947,-524,1813,-826,1184,-2006,1077,0,-2844,796,2457,1696,-4140,-3305,971,2387,-4941,4812,3828,-631,-1619,-1064,142,2315,-1148,-24,-2274,3037,-1232,-5332,-244,-2170,-2058,124,-853,5087,790,-1826,-1674,-4545,-4238,-2056,1089,-188,-2529,-3034,-1125,1547,-8496,2683,-2177,-5737,-2215,-3569,-2575,770,-3845,-3005,512,3129,3229,7099,-706,2839,5107,-1268,-2553,-237,-5034,-228,-3334,-1210,-8222,221,-1931,-1433,-885,2144,2705,-4360,575,4025,85,1707,-4172,2337,-2028,335,-4831,68,482,2941,3808,3361,-4775,-4873,-1981,2897,-3898,-2565,1250,1215,5405,5151,-5288,-5039,-838,1853,487,3332,-9858,-2866,4238,2386,-447,2810,-6513,-4174,-604,-292,50,-3752,-4484,-1281,5405,156,1278,-787,1674,-1536,-3449,2448,1502,-528,1516,256,-1337,6909,-3627,4636,2012,-74,167,3742,2751,6660,2951,4,1466,1429,4697,193,4943,1441,-2839,5234,1582,1499,4963,-541,3144,6269,342,4455,-16,-9482,-504,158,1877,1346,3518,2019,8837,1864,-209,-1523,13,-66,974,-357,-1280,-614,-791,3803,1474,-302,-2119,1604,-203,513,3273,-8125,1218,2402,3269,1326,1169,-1855,-4006,-3884,6113,-1430,3510,-4572,637,-4428,547,-3308,-2210,2475,128,3393,341,-322,4511,-383,-17,1087,-1160,544,-4133,-359,-3559,505,-259,-682,-294,-3889,5688,-6215,812,-2602,1621,3315,-660,1095,-1940,-1270,7163,-3237,8671,4533,1187,-584,6562,3923,-66,-2036,10781,66,1030,3217,1479,3859,-2941,8193,-1837,3776,2260,327,1121,7807,-3525,1457,-1550,-4050,-2651,1033,-471,-1061,-4584,-1510,-3288,823,-2182,-197,225,-9443,-183,664,-218,3149,-416,-654,-266,8037,-4270,1094,1816,-2895,6245,1568,-2507,1945,-5688,3286,1072,-2304,3051,-4199,-14,5625,1911,-1112,1495,829,-2668,352,1947,-1787,-1486,4768,-988,-1759,-3166,3603,-2498,2015,-2858,1700,-195,2121,-5776,-881,4482,917,-3159,-2617,5849,-244,-809,-50,5024,-198,915,-933,1464,-1641,4807,4941,-2485,2514,2551,-3740,559,245,-6313,-741,980,2408,-513,-6523,-2261,-4511,-2807,-5327,2951};
    Wh[73]='{-1386,-897,-1396,-476,-40,2263,3083,-146,1929,-216,6855,-4580,497,4272,-375,839,-4892,-1192,-258,1146,-3591,131,1138,2658,611,-306,-61,-2169,2028,2712,6088,4020,7421,1285,-809,452,-948,4028,-3784,-1611,1566,-3232,1710,751,3679,-2169,-3054,-2187,2106,884,2124,-1123,266,502,421,1093,4631,-3623,466,8012,1846,4272,2993,-3173,1763,591,1488,1130,95,-2136,-3593,397,5297,-2147,588,-2653,1912,-3979,1531,6865,-1520,-4357,-252,-1020,-1888,922,-68,2456,2907,880,-162,437,3325,-1711,-261,1199,1129,-406,-513,358,3857,-1251,2861,-5043,-2844,228,6220,-25,2802,-1976,1738,-6835,7744,733,3317,2266,4099,2600,1800,-186,-1298,174,-4755,110,3886,2149,3168,-524,1370,-4912,-6977,4819,-4260,-4812,-7758,2556,7167,-6318,-4155,1011,899,1072,811,-1011,-2849,4211,-3305,4643,4641,4926,-1815,-91,-547,6147,-299,-4704,-1051,-259,3867,-6113,-5249,3359,4760,1091,3950,-2841,-2049,1624,731,767,-1368,1093,6752,-2736,1834,184,-1213,595,-892,-953,-1264,3295,-532,366,1188,1177,2585,-391,-4516,1784,1341,293,3188,2066,-4338,-881,-2491,541,7695,-3020,1435,100,-5395,1159,4277,-460,501,181,5717,1629,-1774,7729,1927,-1475,239,-874,-947,-4042,-2222,-5566,-1291,6166,1512,-4892,-474,4020,6157,-3994,515,-9106,-3027,462,4218,-2292,-1034,6025,-3867,720,4431,5449,-4338,-2088,1467,3229,-3039,2211,70,-2822,2509,2890,-3652,-570,23,-3122,-4733,-6420,1368,3278,4665,-10019,1065,2805,-3610,2946,1339,-426,-621,1796,-1107,-9614,2619,4428,1950,1828,-1015,502,-2512,-2133,72,1036,2802,5361,2700,2702,1253,2885,-1185,488,2910,-722,-3237,1910,-3205,-2578,-299,-3413,575,-1015,3103,1594,2673,-4934,2006,-2741,-4096,1103,-8002,-2406,-822,-3439,-2626,-5366,5937,4470,1256,2687,5019,-6699,442,-6416,-178,3537,2302,-3864,-1246,3798,3547,-3325,337,-1462,2360,2712,2919,3671,-598,3505,-252,944,491,-3674,280,-658,-637,-3161,-2202,-2788,-422,2482,-4787,1317,-1340,734,-257,616,1879,-58,10556,4147,-7714,1745,-2919,2091,399,6918,-853,18,792,2004,-2451,-6376,-747,5263,3715,-4160,1621,-3212,3735,-1542,-1111,3996,-1781,4643,-6889,2673,-2958,-1864,-3693,1372,-562,-1805,-1364,105,-1770,182,-5532,-2216,1843,-1210,-1222,2136};
    Wh[74]='{230,-1034,-1254,-325,-2612,-1428,5019,-946,85,-961,-905,-686,2573,2744,-4208,-1820,2,3156,2012,2944,-1407,1728,3576,-216,-2030,1729,-2844,75,2111,81,-870,9624,3513,-773,-326,1345,-854,-784,3867,373,-733,-1730,3017,-48,4787,5512,-3041,902,-1333,990,678,-2302,520,2695,-922,-1317,-1221,-179,-1970,2609,3068,3767,2651,-1538,-2014,1043,222,294,-61,-115,4426,786,-498,-1820,-129,1972,2988,-1152,6586,-3793,-2155,-3969,2349,-3391,1275,170,-1006,-2062,2668,884,-126,-1383,-939,217,1967,-896,304,-1680,1435,2749,-459,2636,2966,707,1365,66,1673,6586,4711,1370,-308,-2307,3618,2186,-2741,-786,-2739,3093,-5385,-1165,2427,902,-639,-2023,-5380,-1536,-2485,2322,7451,-3078,-2998,-2083,9028,-310,3688,2275,-3364,-1893,-369,-3208,178,-764,-720,2575,4777,-567,1680,4270,-264,1512,-1673,-2458,-1097,-404,-380,1785,3269,-1312,-568,-5771,-3232,3320,-839,-3837,-1915,-509,-2309,-4064,198,153,-4936,-2285,447,-1145,-42,-1583,-1715,-520,-1286,255,-1751,-3349,2108,-5327,-977,2529,1237,-339,3688,3674,-751,1575,-2687,6025,1650,-4355,254,-5776,-427,2814,1617,718,-2135,-1387,-3752,2023,-726,758,-717,1322,-2416,590,-760,482,809,-7041,6489,56,-327,6083,790,2027,-4992,568,2570,-1777,-996,989,3627,-2385,-4350,3757,-7036,-1760,-5737,1179,1348,-521,-2261,4296,-168,4526,-1578,2287,886,1600,1064,1809,-1201,1625,-30,-3068,3527,623,-913,-1533,-299,-1800,-1485,-3476,-4968,-6860,-1230,-5703,-4426,-368,-1845,-5092,-378,969,2636,579,-4128,-284,-1503,-522,-1794,-805,86,-1119,-3542,1052,1975,4382,426,-7500,264,-2215,-6000,-1933,-5576,-2702,-412,4550,-1224,-4245,-57,-1654,680,-914,578,-3540,-1386,3034,-1910,-4987,574,-933,1322,1300,1558,1520,-1861,55,1649,-507,7871,-17,-6186,2327,-4707,1067,2497,1444,-1405,-3041,-2661,-1223,-1053,1373,-5927,1373,3063,1018,2437,-4555,208,-1810,-2143,155,-2197,-2165,1126,5170,-53,2666,7490,-3247,-3405,4074,3903,2587,783,383,859,577,-1729,-13154,-3012,1486,1507,-1761,-48,-2318,1313,2507,-4633,3225,-3471,-6230,5732,-3974,-1818,-3283,-140,-1381,5712,-620,661,574,-4826,484,6826,4450,-3745,3625,614,112,-254,1148,1624,6318,31,6323,-1505,-11240,-1284,-288,367,-425};
    Wh[75]='{1921,2963,-662,1229,798,-1553,-2521,-440,1339,-2175,409,-709,-5751,-1512,-5019,2324,-4826,968,2445,-1824,242,1423,-6694,-543,565,-212,-1669,-1838,-6391,1159,2338,2342,-594,-4099,-2232,-3796,1346,-2502,-3071,-5039,-977,-387,1680,-3481,3132,1038,2597,1450,-4611,1689,-404,3989,-9785,-1633,1336,-564,-2480,-2700,1678,-2210,-1652,29,-668,394,-5429,-117,209,-908,3874,-159,2423,-3637,3359,2302,1418,2502,-4189,2307,-127,1534,-1248,-5781,505,-7075,3820,-2731,24,578,4492,1413,100,-5175,592,-2619,2739,1069,429,-368,-8627,-2213,-4045,-704,-3088,-7246,615,-110,-900,670,1352,-2590,-1992,-10585,-463,2418,2441,2622,3803,4230,-4953,-659,616,-2479,-2093,-2568,-5927,2512,529,10947,-1697,-5380,-1719,359,1911,-938,-196,-3083,116,-1227,1152,-1711,5859,-1340,-3254,2064,1190,2666,505,-2792,4243,-4445,3615,2080,-764,4455,3359,-1883,-1254,2305,500,-1112,3579,-3593,71,-1583,4758,343,-2792,650,-6972,2196,1832,3088,4506,4016,1091,-479,55,5947,-3022,1549,5634,-2304,-520,350,1259,3193,-790,-2797,2875,803,-134,4448,2551,-4384,-4082,-297,1385,-292,-2454,-2250,-586,957,5336,-7666,353,-1301,250,429,-4448,1654,-5537,3041,-2028,-5390,-2922,-162,-3574,2459,-426,-13964,2475,997,-252,-2203,-1031,790,4262,-833,2237,-807,1117,476,3833,326,-2093,544,-1816,2207,3308,3627,10800,-1107,-592,2590,4262,-2180,290,-2971,-3637,3137,-82,4375,-44,-114,2924,-1268,1999,-2083,4626,-2580,-1934,-3405,5771,-1071,-1635,-3125,-2939,3845,-3562,3295,-2113,-737,-1677,-1763,-3991,-2103,3625,2294,4201,-334,-1480,-1771,-7792,-6137,-3083,-228,413,5141,834,1700,-4748,8349,1247,-3610,-2924,-7036,4724,1866,-6948,280,-386,-2578,3837,-3327,4741,-4086,-1785,-2692,-1070,1787,-346,-1741,-3508,12812,571,4926,-3339,89,-6235,-4248,4956,-1722,-8916,-5151,-4155,-5800,4350,2486,-1196,-4531,-5903,-1966,-2788,-1233,246,-5239,3291,-5527,5122,-469,1796,-596,-728,-4377,-311,-125,-2320,5058,2983,275,-3679,613,2744,2222,3178,-558,2912,8002,6289,886,732,428,3410,3305,335,-1719,3530,-5263,-3098,-12470,-4316,-3676,3579,-1781,-5634,1759,222,226,608,1004,-3215,1042,930,-801,-1468,1712,441,4372,-1188,-2349,-7031,-1104,3327,-3527,4152,-144,-2275,2403,-314,-2521};
    Wh[76]='{-4970,1343,3413,6181,1835,-1668,49,3625,8696,186,5415,2641,520,-2092,4384,1466,1746,2265,1611,1120,-4047,1568,2463,1213,-4221,-4013,2386,231,2612,7275,2102,3535,3754,950,1,615,-2044,-1416,1494,-2541,-6,1104,536,-1309,-5258,4592,9663,-1937,1737,2697,-181,-1231,-2807,3937,1804,1879,3771,-1055,-3173,4401,2354,-2224,783,4074,-1350,2829,-3691,1240,3007,-5019,-2296,-3491,-447,-321,4157,4816,-6181,462,-1826,-4936,-2133,1151,-2546,4716,-3627,6127,820,1993,3505,-3208,2619,2788,-1665,433,-7949,3771,-5048,822,717,-2352,4631,6166,-1779,2666,-1314,2357,3542,10390,11962,-1973,5014,11552,4853,-5532,-565,-3530,2927,17558,-1445,-1790,-3991,-6767,-9555,-1032,3337,-8750,4133,-187,2675,3923,4047,-7500,-3342,-1917,1904,5258,-8413,-575,-114,-1176,-3884,5571,11992,-3449,3945,-3583,8095,-9648,13125,1314,960,2875,-1855,5815,706,-9291,-6752,3718,5883,-2104,-7539,-5092,-2470,4494,-3801,-7871,3925,519,4831,-6284,7265,7475,-3896,2100,1760,-2954,-1149,271,7441,2033,9672,-8881,6098,-2785,-732,1541,5278,2978,4291,-7500,-8574,-3259,-1358,4528,6870,8222,-704,713,2512,-3847,-1285,3322,-475,2929,5322,-1713,-708,-4118,3315,2868,-7749,2303,-1039,7265,-4851,-2622,2797,1560,3811,350,-2783,-808,2624,-5966,3112,111,682,-2644,-3308,-3745,-912,-406,-2822,1130,-4074,1955,-7612,497,4687,-290,183,4387,-621,-540,1405,4851,2810,2213,249,-422,-6157,-2482,5756,3583,2321,-9067,-1838,-1796,176,-6411,507,889,1729,-7006,139,-1431,-6801,-3356,-2242,1484,1304,2709,3571,1557,560,-7441,2414,-3850,4367,-631,4238,4467,-5380,2629,-6650,-7978,-1248,2093,-2900,-185,1033,-7539,-8754,-1401,2697,218,-4721,-1810,-5815,46,2800,-2907,7377,5209,2595,2019,5400,-763,2810,-613,4042,6166,-5053,5327,1010,1026,9150,480,6342,2531,8100,4492,3413,-3874,3598,4265,3776,-4497,632,4626,7744,3276,-1384,1039,-2314,2071,-2398,-2373,1044,-5410,-1656,-1035,415,-4453,-4758,2539,-176,-1490,7377,-3105,-2299,-3886,-830,-924,3176,2441,1983,-2247,2357,4731,-711,2622,787,2800,-4553,4870,6118,6528,1669,-4299,-1828,-2988,751,2310,9692,-42,1203,-1398,-4987,2495,9736,3652,2183,2731,-7475,4204,-3134,-132,7280,-2814,-1240,-6992,1067,221,-3244,4321,1442,1322,-1119,-3503};
    Wh[77]='{-3835,4763,-5991,1262,715,2283,-5097,-2758,-3027,2238,9311,-1701,964,103,-1616,-5195,4047,2020,581,1458,2849,898,-167,108,888,-1012,4619,4538,10195,-2817,-2452,2453,807,-485,-2282,-833,-3430,2423,-2404,1066,-404,2709,-2203,653,-2169,-3476,1788,4633,140,279,3371,3710,101,-657,-1401,4094,303,-8232,5019,-6235,1817,-1244,-2832,-1770,1250,-213,-695,-7949,-6059,1342,4411,-7255,-1392,734,-1281,1311,836,-3491,-2973,924,3051,-3459,3828,680,-6826,-1976,-1227,-3769,3122,-3830,5498,110,-1676,-4350,151,-1367,-41,5322,870,5659,6352,-4360,1193,11093,1513,-3625,-5180,-1243,-6372,-3791,-2153,-519,-1160,-1213,-2158,3266,-2480,-6791,4135,4145,2163,3823,6547,-5649,267,4531,-10791,-11416,409,-315,-1771,4528,6049,-6035,2658,2181,7036,3483,2331,-3005,-3564,-3112,886,3266,-135,-350,1375,8686,-192,3369,1707,2113,-1907,4270,-646,-4187,-364,389,1444,9331,-1304,1126,-4006,5805,-1705,-4106,2281,-1658,-1419,1043,5000,1551,3979,-5898,-4284,859,-4174,462,1246,3227,2353,1191,-2202,2319,-1402,3359,-197,1536,-5551,3769,6010,1499,-1525,1702,1284,8383,1291,-1408,-5234,-249,3247,-1589,-1666,5703,-413,660,-2651,-4902,-2648,-1710,2438,-297,-829,3881,-2430,3583,-406,-7675,-3554,-1085,-1263,-825,2785,4431,4902,3706,-1549,-2741,914,3666,5058,-5532,2425,4013,-84,-1232,3686,103,1383,-1068,1617,-1624,356,-3562,-1945,2431,-4511,-3315,3337,-494,-623,2568,784,-5815,-1027,4245,-3776,-5747,-6430,394,1074,2346,-5278,-1071,-3352,1180,2171,-836,-440,-1078,294,-7119,-752,-2939,1794,-870,1700,-2342,2795,488,-2243,4191,2203,1019,4550,2980,-2265,-6625,-2875,-1965,-2690,4645,2775,-9047,-4233,4038,-4953,-2910,-1906,1145,833,-997,-5317,3127,-5644,-5722,1561,-5317,-6479,6645,581,-2070,371,-1447,-3652,2269,-3874,-2001,5332,-547,-549,637,-6777,2408,3662,5053,6376,-1724,2025,2125,3190,-1545,-3508,1994,3747,3237,-496,1940,1424,-2634,657,-5634,-2081,-327,-3305,1000,26,9707,-9296,-41,-7319,-2836,-2570,1966,-944,1485,-2177,-2690,2543,-3205,240,4235,985,2237,-1068,1258,-1210,-2585,3339,369,-564,912,3315,-2829,-2792,-1195,-2346,-993,1436,-6669,-4829,1182,4501,3225,3186,-6005,-10,-3977,1756,-734,232,1966,2648,-597,-2812,-1362,-2243,-508,-4855,1484};
    Wh[78]='{-6972,192,-2509,99,-705,-1370,-2546,-2261,-268,-611,-5053,-6162,-1968,623,1228,1181,-977,-3393,-5053,-6474,-4099,-1622,3496,-4758,-2565,-7231,-740,-1367,-3540,-1643,-6157,1534,-2626,-4528,-2413,953,-2232,-755,-2451,-3366,-2019,542,-290,-4790,6938,2268,-673,-1373,-2590,9716,-607,222,3349,4687,-2459,27,2108,-2447,-1195,802,-5004,-2644,-2687,-182,8198,-6992,2607,-1204,-4707,-6474,-3991,-4357,1447,2121,-6562,-75,-1834,-8466,4228,574,-1065,-3793,-2026,-2362,922,3833,46,-3027,-307,-2399,-2216,-2187,-1943,-5195,-4204,-2200,-1037,-618,-3029,988,2320,5908,3891,1634,6718,1046,5410,7783,1527,-98,-982,4477,10390,4809,-709,-885,-734,-2369,6284,579,2048,5351,-10312,-2255,-1900,-1027,-2739,-3144,-6665,7011,-6835,3811,-3413,-1795,-83,1018,2346,6054,4755,-5981,4423,-2431,-392,-1229,1308,4299,1279,2851,1594,-1025,-4479,-1192,-24687,-431,-5649,5156,-920,-3344,-4748,-246,-9868,-5229,9155,5756,549,7314,-2282,-3664,2186,-2719,-3208,-2966,-1889,-2467,-487,-2246,3000,-2658,-11220,855,-1873,2634,2160,-1483,3452,-3186,-4736,-2749,4877,1550,-7158,-2885,-7778,-1073,2104,931,-1816,-2841,193,-423,570,-3737,-832,-3181,4453,-1043,-2663,-2188,-290,-3256,-3503,3603,-6645,289,-3620,-8920,-3815,2927,-5424,-6445,845,-2666,-8374,1900,-6254,-11777,-3415,1067,-1285,-2141,-3837,-631,-5825,-726,-3454,1490,-3847,1222,-5576,-125,-452,-2932,-758,-3247,-9692,1579,-2440,-1934,-6308,-5751,-5717,-1359,12675,-7612,1458,607,-3593,7812,218,-2476,-4675,-6450,2658,2854,-6982,-8139,-81,-4841,-1098,-4892,667,-7124,-3173,-690,-3583,-4572,833,-4653,-6757,-242,-2193,-1508,-6855,3789,1682,-6606,-4086,-9204,-3386,-9692,5971,-381,-2224,-6455,-4824,-3620,-2500,-3486,699,-7099,-6997,2543,-792,-8325,1597,-1593,-10693,-8613,1823,-884,-5039,-9775,-11503,-4113,-6025,-1407,-9677,-4929,-4592,3483,7158,-3664,-13994,-1700,4899,-2526,-8452,-578,-5327,990,-2685,-2746,-318,235,-5424,1021,-7651,1052,-2287,-4721,3417,1816,-5551,-1871,-8066,-2451,1611,-8251,-4133,6459,-2152,-2464,12548,6918,-5375,-3713,-5776,-2160,-2104,-3398,-13027,-9536,-4895,-1028,-7089,-5454,-4287,-1660,-2153,2020,-6567,-442,1893,-2076,-5014,-6333,-3415,-3198,7875,-3820,-5297,123,3093,-2307,-933,-2827,-9765,-6948,-5668,4482,-838,-3452,2529,1394,-5292,-1263,-1912,-2763,-9355,-4768};
    Wh[79]='{552,424,-745,-1556,-5131,1430,-2437,897,-2902,-1431,4436,2006,5341,-947,-3669,1622,-5117,-2895,-3366,-331,2387,-4841,3442,82,742,-968,-3283,-2163,-3063,-5336,214,1955,-5273,2653,-2183,-5078,-5556,-2093,3239,203,-1573,-5688,2386,-946,4045,-1032,-4291,4055,-2059,-211,4023,-4794,-200,541,-1555,-97,-2998,2966,805,-2069,2531,-512,-547,2368,-1522,3872,-1831,-4990,-2687,-229,-1850,2492,1132,-726,-352,-2347,1160,1540,5712,80,-791,-7456,-433,-1872,-710,818,-1364,1424,-1085,1427,-3129,-5434,3088,1678,6303,-3305,-2753,-2998,-1048,-3066,2707,-945,538,7128,-5336,-12,-1608,1518,-2719,1395,-6445,5292,-3405,1104,514,11,-150,-3166,4816,3615,2971,-1271,7705,-5390,-890,-6337,-3496,-2763,7006,4177,2939,-2893,-1785,-2432,-3220,-2939,-5214,2731,2322,5595,1379,-1417,3247,-4001,-3020,-3305,-1702,687,-3564,-1931,-850,-1342,-1434,-3007,5136,2426,-5751,-2841,3007,-1948,1971,2976,927,-3256,-229,126,-675,-1335,5292,-1181,-6616,-4531,-6250,4990,-133,-4592,140,-1706,-3518,-1723,1151,-558,-867,-279,4516,2231,-2080,-971,899,-2651,-809,-875,-2149,282,2648,-9111,-118,-4851,-5551,205,-4716,2271,740,1855,-1230,370,679,6489,-1190,200,-2424,1646,-2469,-1922,5673,-3229,6264,-5214,3027,-1553,1627,3432,-3549,-376,-4685,2568,-5131,1496,-6005,624,2137,-3291,-484,-3430,-9731,-619,-6459,-364,3881,-1801,1520,2047,-5595,4252,-4450,-1531,-345,4238,1928,324,692,-2966,-749,2954,496,-527,-2286,-2117,-2122,745,-1218,2770,2261,802,1987,2521,-3225,-6083,-1372,-75,-2797,1517,-1262,4006,29,4511,-2951,-605,3483,-1121,4602,-2084,-200,-734,-1490,1621,1519,3251,-829,2697,-2019,-4479,1372,284,-2722,2675,-4091,798,-5024,3647,433,-181,102,967,-3493,-1423,3635,2391,-3720,-154,4245,696,1739,-6411,-713,-4226,3994,-2014,-3781,-3405,-4094,-567,-1895,-1062,-1329,2171,-2976,-4267,3176,-3881,-3205,-2780,-2326,564,-461,110,-2753,-2164,-1046,3801,-2995,3452,-233,-118,186,3381,4240,-2221,613,5283,6401,1389,3981,2358,2656,9213,-1435,633,-4941,713,148,4287,1342,4841,592,4638,-801,-582,-5927,-5336,-148,1149,-3510,-1177,-5483,-1802,994,-1036,-1468,226,1217,4013,6674,3706,-1206,4953,-2183,1704,2509,3166,-2131,420,-673,5415,-236,3339,-986,1065,185,-722};
    Wh[80]='{327,661,-4270,-3264,-709,2039,-677,-2374,1418,-927,-5175,-135,2236,-3266,-6840,195,-5610,-4338,-221,-786,-1949,1152,3845,-1958,-61,-3103,-3420,-949,-2105,71,-2851,1859,498,-560,958,-3044,599,-812,-1078,-2524,2166,-3007,3540,-6157,1712,-268,-2780,-24,-1864,1417,-3056,1331,417,-1409,629,2912,-221,714,-3549,-3208,35,-1613,-176,53,-5327,899,489,-2900,-2585,-885,271,764,399,-4453,-375,-2481,-3381,-3601,1239,81,4350,22,-1359,-3286,-2031,1084,2539,989,2822,284,-3491,-1561,-570,5366,-474,-1077,-1157,-5268,-5761,4057,2658,3286,2807,-7314,-1608,-3740,-4531,-692,4904,1679,-2473,-3657,985,-2192,-4211,265,-1697,-3178,-202,6406,4116,7280,-316,-416,-1254,-253,-7612,-791,1917,2302,1677,93,-1024,3366,1588,3791,-2663,1619,-2480,599,5034,1962,1300,4211,731,-3613,-2075,-6411,1376,-2409,3012,-1356,-293,-4650,459,5737,3522,2761,-2425,-9155,1435,5664,-2033,-4326,207,-2099,-2227,-312,3994,-421,7490,-2069,-1776,163,648,-3854,-2722,-1280,2078,776,-3593,-2927,-1915,-3420,328,2595,-4748,-2863,1435,3674,-1264,5058,-6210,-455,-3188,4511,-89,-3342,-353,1243,44,-930,-1092,-529,-452,1816,-980,-8315,-6772,87,-1538,4553,-2369,1113,38,-4526,1343,-2607,-2128,320,-3269,-1531,7187,2709,1114,-1972,2005,-3320,-1398,-4160,712,-1093,-6396,671,-1359,-1435,-2065,369,871,5180,2758,-2307,2827,-370,4147,614,5756,-227,-2430,-531,-1195,1998,866,320,390,-424,-770,1369,-713,3930,595,-6894,4992,-434,-3627,-150,391,-442,-3962,-1407,480,5991,-909,-2310,-3364,3896,-2687,769,-2322,-3388,1152,2030,1262,-704,-2227,-1395,-1408,-4758,-221,-1276,1647,1445,1972,2288,1632,-6054,730,-3256,-1846,1687,2504,8227,50,-491,-469,-3308,-6396,-2426,-2968,-2100,77,-1683,-1314,-4885,3698,-3857,10781,-7622,-428,-3527,1402,-1201,579,1535,960,673,-4433,-581,1,-3403,-3264,1359,889,-879,-1450,5053,3986,-8535,-2047,3361,2536,-5458,2458,-9028,1600,3701,7036,-2067,-8017,-2536,836,-2041,-5439,-3779,6977,3046,1096,8823,-1693,527,328,-3486,-1599,7963,-1181,5883,-1224,6738,-5239,-994,-4270,-1015,-3381,-3381,-1262,-4233,5292,1024,-3251,-3281,3989,4868,326,-1593,-4101,1705,-1545,-1580,2108,-487,692,136,210,-4672,-1380,-961,7509,-2856,-2756,343};
    Wh[81]='{716,-975,-1533,1987,-2010,-2902,-7338,4003,-3723,-193,-4375,-191,-2612,-1650,-7094,-3383,-10126,-3796,-5517,-284,3293,-4533,-3769,-1552,1101,674,4074,-1591,-5869,219,2252,3837,-380,989,-5322,3310,-1079,-4365,48,785,-3254,8569,914,298,-2008,-1466,1354,1408,3959,-1249,-5351,6821,3300,5219,1585,-9125,-1751,1813,-1026,-24648,-2514,-5039,3317,-6811,-1719,501,-1831,-7456,-4536,-151,-2268,-4082,-1306,-4982,-3410,-4167,-6386,-5122,-3657,-225,592,-487,-3457,9096,-9599,-5415,1697,1282,-6489,-4887,3352,-9423,-5307,3535,2366,-3586,-2797,2348,1204,1816,11005,-3728,216,3950,-3420,-390,-1971,-3515,-8413,12119,2402,-170,823,-6142,-593,735,1949,-10087,-1486,2575,-18,913,-2856,-5463,-8496,-1223,-9702,-7001,4753,-6601,9179,2810,3342,-2277,2445,1135,6616,-628,-6845,5400,6582,-538,-2194,1594,603,2304,-1503,3242,5810,-3266,-3862,728,-6030,2224,-4645,15625,1861,6430,-5883,-11347,10966,-469,625,730,-1805,-7836,-5029,-7192,-2401,-1031,-5468,487,-795,904,-3457,819,-1214,-208,-1420,-310,2152,-122,-4248,2709,3640,240,534,2095,20175,1265,1517,6562,4553,-7109,-1284,-1788,-3913,-3110,-6357,-2741,-2489,-751,6870,-1311,-709,-1128,1821,3442,-708,-7353,643,2484,-1972,3100,-2226,5844,7207,-6381,2783,6860,1756,-3535,-1080,-1026,2685,-621,-531,1263,1821,3356,353,-2785,-3903,2308,-1495,-3901,4956,3696,2338,-3515,1604,4340,-1268,-747,3442,-687,-1252,6489,8315,1479,-833,4699,-2595,-4628,9443,977,4172,-1643,1663,6708,-951,-2333,9980,-3833,-2117,3427,3376,-1561,-2570,2839,-2031,-1636,-4794,1433,-2148,4135,-3715,234,499,3925,-7167,-6772,-1588,3869,4978,3623,-450,-4621,7890,4565,2080,-4924,2570,-1711,-2915,-487,4069,-1884,-503,-964,-6982,5766,2164,-3371,1231,-8740,1022,-1163,-3164,861,2727,-65,-1093,-3898,979,-8588,6596,-2409,-1512,-5170,-444,-7050,-2132,8339,3447,2043,-5800,-4611,-3315,-1685,-4687,5161,6777,732,-571,6997,-4853,-5727,1184,-4431,-1882,-7119,-4741,801,251,-1844,2819,4660,-6645,1726,-2939,-4165,211,497,359,3007,-2604,4804,-7114,-8071,-1442,-14062,1579,-741,682,2543,-1910,2479,-670,-2529,-390,2282,-12050,-3808,-1011,4243,1737,-2758,-3862,-7475,-3283,-2854,-584,-820,2722,-5102,98,-1833,-1018,1145,-2220,7089,-45,-368,-974,-204,771,-4985,-1573,-982};
    Wh[82]='{-112,2634,-2678,1950,-203,-1629,-2639,-912,110,119,-3945,-1226,-2534,-3872,-3378,-645,-864,-1464,-858,2998,-2247,1831,3281,-1820,-2145,-1336,-6303,-180,-3164,540,-568,-9560,709,-412,4111,-2004,3908,-1436,2192,449,-708,120,-944,2261,1857,502,2910,-2463,369,-1477,758,1260,-1550,4775,2355,191,-1944,-2727,-2731,2761,-835,44,731,109,-11259,-2011,-1840,3569,-2196,2049,-1796,875,839,-3469,-3259,3369,3139,-3012,-2172,-7714,-2180,839,844,-4245,668,2602,2337,2587,2500,5766,-386,-661,1793,4489,3400,-611,4799,3293,-942,-194,-1706,-1030,2819,6665,621,3837,-3999,1089,2597,-2142,-4013,-206,-6723,-5361,-1979,-8725,1578,9501,-296,3400,-1252,-4606,1069,1055,-1151,-6162,4655,3791,-3000,2462,-3391,3874,588,-1054,-6059,-774,-5053,3552,-57,-3134,-3291,45,-2856,842,-618,2351,3781,5610,-2785,2795,5058,1307,-674,2871,6430,-279,600,-1364,-1385,-1621,-1030,3293,-2770,-5903,-4985,1696,3366,533,460,2524,6210,93,2048,-2099,-2509,917,-2165,-268,-1535,-4006,-1235,1925,298,-4638,103,-1464,5317,-1016,-221,-1150,-2121,-345,341,-2880,-307,96,-3142,-1556,2109,747,1275,2130,-48,-1065,3984,-1227,3369,-2739,-1834,1557,4785,3249,-3547,645,-1068,1223,3068,8891,-276,2092,-2897,-4035,-3142,-3215,-1486,-4091,-3137,186,-629,1925,516,-1348,-3415,2166,1209,-5883,-3039,-935,-3144,1796,5747,-790,2091,-1855,2600,2709,1806,-950,-4675,3137,2932,3161,2384,-2954,663,2266,-3386,4296,-791,2934,1518,6279,-959,1003,-121,-1518,1156,461,-1030,1883,1824,-190,-1939,-1158,1466,-4819,10029,-3786,34,5805,-1834,678,5327,-1339,-395,3457,1166,1154,-3813,175,2919,1828,-2416,275,-228,-2202,597,1329,-2504,-634,3171,-425,1260,1331,-1387,5708,-2285,604,-848,2651,-1282,711,-4458,-3642,1790,5615,-5600,-1328,3234,-1306,-3198,-5004,-2946,-2565,1929,-949,-1423,5219,-4365,-1632,-1822,-2019,2249,3671,3903,-7661,-3576,-762,-3403,-903,-262,2761,939,-3574,2585,-334,-6416,-3007,-2427,134,-517,3835,5161,6450,-1018,-3728,-286,4985,3298,4919,2482,-1654,1855,1246,-3098,3691,-1966,-4108,2199,2973,-1773,3864,8071,3308,2590,3149,-4304,-958,2060,2900,-2296,-5371,5205,-1034,2352,-1028,4047,3698,4724,3203,4494,-1663,1871,-6059,-2504,3535,2399,-4448,-3039,6186};
    Wh[83]='{3012,5683,2176,-2802,1644,697,10468,4553,461,-78,5273,-3449,1542,-7524,138,3447,-4177,3117,2238,-2429,2034,-1632,1857,858,-1976,-2277,-1921,1235,2032,1831,5712,-3098,11132,3984,2054,-1152,2524,2927,3200,-88,4318,-1047,-157,-2059,108,1228,-2895,-6533,786,-106,2441,-1007,3833,-1030,919,-422,901,-457,427,-1984,223,2502,2438,6689,1111,602,7436,5083,2775,-3710,507,-8300,2471,21,2299,524,8437,10205,3469,1988,-4096,-2014,10283,-6191,7241,282,-2026,-2062,1779,4252,-3181,-605,3632,-3332,963,-5971,1507,-8637,495,1722,-14814,416,-2132,2386,7895,-342,1678,11093,12929,5615,-651,16132,6689,2824,-2087,1893,232,1223,-6088,-6333,5639,-7363,546,-340,9487,-8237,16748,2401,1174,-335,-404,3000,-2239,706,-3769,-1161,2944,3857,1802,2512,-9047,-4645,567,1490,1617,-1104,2027,-2403,11308,2332,-5688,-3481,3278,2766,7729,-1774,3193,-2313,3696,8940,-3835,2486,-4770,5771,3378,6313,-1932,3874,-2915,-3884,547,-1333,-2005,5351,2165,772,2445,1641,-1440,-3627,63,-642,-4353,-4645,-1176,6645,3393,-4672,-9033,8334,-6123,-5541,-3208,673,6040,-8310,-4772,6748,8618,727,1199,7055,-3408,3364,5185,-2065,323,-3581,-411,10605,-1518,1397,-8325,255,-5410,-4643,-474,3063,-6840,-255,5424,168,255,-1610,-5000,-1744,-707,-3039,-1864,-711,-6,-1591,1381,-2089,-3974,-4328,-786,-5019,1976,4250,-3134,203,-1138,9702,-2459,-1909,614,-584,499,405,-925,3449,2382,-386,-5708,650,-786,-1523,-236,-260,2829,6811,-6416,-4379,2778,4406,4206,3618,-1855,-1982,2413,875,4936,2912,-640,4433,572,-381,-298,-1120,9462,3483,2829,-3139,-2971,3933,-3645,9399,-3955,-8027,-3215,-1419,3188,4377,3083,2636,974,374,-696,-5917,6728,-7646,2578,2707,-2612,4040,7666,3259,2763,-2775,1282,453,-2954,10419,-2476,4873,2536,2109,2229,4602,9921,3581,1429,-3525,-260,-4638,4475,770,-964,-394,2443,4355,-3237,-807,899,-4904,4086,-691,-4685,-4895,2028,3454,-1636,-5664,-1590,-8154,-5903,6083,-287,961,398,3562,-1407,-7646,-11328,-3176,4394,-394,3876,2595,-3493,3920,-886,2312,3483,-3095,260,-2983,-2004,-8417,5258,-1679,3676,6958,839,-503,-4294,4255,4387,4279,-1147,1754,-1671,-4089,4245,4326,-2978,5986,-228,1070,1486,-4580,8427,1175,6015,999,1921,13457,-646,-736};
    Wh[84]='{2399,-9931,-1389,-409,-3188,2797,1556,4177,-1322,-44,-148,-239,987,407,5488,-4260,-3669,2230,-1452,944,-32,-1547,1750,-2536,-1771,-1041,-920,-3352,49,-6982,-1975,-2296,-7753,628,-629,-3745,1376,-2592,1011,-6064,908,-543,-1680,-1351,-3862,-38,-1068,-3710,-1350,322,-497,4370,2479,490,4165,-1697,-2934,2607,-157,-9697,6640,-2219,234,-696,-528,-704,6923,-4772,-1181,4255,2451,-788,-7,-2861,-4189,-4750,-2360,3237,3303,-566,-2792,-9443,2604,-2653,2861,-1368,-2438,-96,-147,-247,-6503,-10556,-5576,1866,-1944,695,-3332,-100,-1898,-3513,-3391,-1551,-1695,-5952,-1577,587,-3789,7221,3750,-5883,-4916,5844,6357,-1818,-4970,-4301,1452,5078,-3869,908,3571,-1373,1890,662,-648,-3100,545,1826,-3508,7504,-3012,4875,1702,3676,7338,-3952,2027,2548,3608,1197,-1112,-498,4926,2526,-3269,-37,-3710,8349,-6035,936,242,-2299,4636,-4504,1345,5371,-3068,-4477,4353,-3107,-2868,-1529,2841,1047,-5117,-268,-5375,1632,-1667,4387,-7128,-2521,-1716,452,-1574,-1909,-2204,4184,2744,-2036,-1038,-9257,-1342,-419,1149,329,350,-1173,-1989,2043,1093,3588,-2021,2009,2399,-392,1433,-6259,-3056,-989,-1183,-1566,1672,3381,-426,1420,-854,-2141,-2927,902,1154,-2453,-6557,-3618,3530,2978,8134,2243,-872,-1118,1815,-7758,-2937,-989,-1750,-4645,-9877,-2005,-2346,496,463,-2092,-1072,-969,-12177,-719,1627,-1912,1168,-934,-28,3559,-3601,-2971,-5356,1660,-3859,8378,-2036,-5561,4558,-1624,1001,696,-1376,-1090,-3276,3762,1495,-3984,6386,2259,-4921,-1005,4077,-1405,1788,-2941,-1268,3864,4506,-5400,-5517,-77,-2902,3105,-1224,-1250,-5795,-1666,-2607,494,1710,3029,800,2792,2033,1668,2749,-1144,-2590,941,-2398,5024,523,3745,4233,-735,-2727,1737,-3308,2629,-1490,-887,-1100,-4829,3991,2460,-18,1762,4160,3557,-42,4682,1481,3208,-5371,3898,-4426,1582,-2178,-3193,1077,-2170,-1676,-765,-6171,-5244,1514,-1885,-3652,57,5585,1363,1074,-7241,-928,-219,4565,-1535,5424,1416,-3530,2797,-4042,-5239,-1556,752,-3674,-289,-3518,728,2724,2768,-2514,-2434,-5737,-8867,-3894,-1519,907,-1600,358,-5693,-1575,-4975,6591,2453,-3435,-138,-2294,581,-4768,2293,-2639,-621,1649,-703,2055,3498,-257,2070,3957,4902,-5112,-4858,-1801,-1784,-878,1372,-248,7055,1095,-567,-2844,-7001,4916,-1489,-4108,-945};
    Wh[85]='{1375,-6132,-1386,733,2893,505,-3200,-3154,-2028,334,10996,-1666,1903,4636,-83,-6,173,1171,2249,-148,2763,-1296,-4689,3662,1804,-6479,6826,4592,2442,-414,1501,3391,1811,1203,235,-1007,-110,925,-1237,2043,-3056,4042,2318,-4462,3588,4279,-4902,-576,-4536,1457,-337,6391,1807,-3293,-97,-2900,3129,2142,-3684,-544,-1700,398,4421,-277,4465,3920,1099,631,-5634,-761,-5029,1386,-2541,-120,3317,7285,10117,-2108,3603,-1689,-1801,-5766,3591,2983,-1200,4855,47,-891,2396,317,1557,6694,575,7592,1155,-1295,390,-327,-1838,-4675,8530,-4221,1744,-12695,-4458,-459,2034,-1898,-2622,1030,-1870,14355,6635,82,2360,-3562,1654,15,3161,2092,-6196,1887,4697,2819,6601,-2651,-1149,-4514,9487,4301,39,728,2504,-5952,9804,2568,8701,440,3935,2695,-2834,5053,2736,-4641,1175,-1748,-4140,2641,-1011,1129,-4555,-5117,-4663,6796,7397,2006,-1457,238,-3237,-600,140,-283,1984,7338,2363,-107,-5097,235,4633,-429,-3125,7304,-7895,1192,-6767,-2648,5849,1938,509,5327,6318,131,-9809,3601,1912,-550,-4306,8627,-8515,-930,4162,7729,-5366,2293,6430,-10458,3369,1200,5156,437,-4501,-2900,-1224,-7622,-188,-744,303,-4887,14003,-2883,-6381,3596,220,6743,-6298,-1340,7158,-343,4504,8041,-1118,6660,9511,6479,861,3281,-848,-2954,4062,-4929,1229,-4692,2687,-7592,1783,1140,141,-379,440,2817,5410,858,-2382,-96,1549,827,-59,-50,-1207,1367,-3505,-2239,-3747,-1739,-2220,-1406,-6733,127,2050,-6586,3454,-476,-5532,-3806,1424,-651,-3940,-1513,-2556,-1047,-629,-2695,3735,-775,-584,437,-2467,-3461,-2077,2053,4067,-902,-4506,-8232,-1697,-1511,2607,-6401,15312,-908,5751,8198,-957,624,2442,-5649,-632,3701,-2766,-1070,-615,1572,-719,5800,3249,4089,-4687,-2207,426,-5029,9291,229,-3764,1339,-2556,-3088,1644,5888,1784,3981,4514,6586,7065,-2583,1895,1185,-2360,-485,-853,631,100,-1462,-690,-2612,1563,6069,-553,-2609,5766,138,672,-4121,6,-670,2648,3454,-404,-3959,-4599,1078,-853,-3266,1304,-1176,4401,-529,2832,-2414,-110,575,-5991,776,-1160,1300,-4257,994,1668,-692,1435,880,39,-4702,431,8647,1159,-2445,3986,4831,982,-7392,14638,-287,402,9682,-3361,3635,2000,-3942,-151,-6000,-1270,1611,-66,-8002,-491,-714,3256,-7651,-271,-4079};
    Wh[86]='{-1676,323,-372,3269,1354,-699,-3623,-2602,3518,1628,3620,1069,1308,-4399,-5434,1981,-163,-609,-4685,2780,-1608,1560,6860,-784,-1556,-4511,776,-428,-297,2015,1069,1275,-697,250,-12,-458,-1535,-166,-1086,342,2729,1931,-2355,-1081,222,-3225,1503,3974,-33,-2335,-3879,1423,-2851,-1205,-2653,-4812,3171,-3889,3449,2229,3137,3710,-4003,-6562,-8461,4147,258,4394,2454,-1768,668,2036,3330,7,1002,2338,5727,5249,83,-1015,-2724,2432,-7084,458,601,-4094,-703,-2761,-503,2709,1434,-886,2458,-1500,2697,1975,872,-667,2922,299,-3867,-2291,2934,1431,-894,-1267,87,-792,1334,-1278,1979,2174,-5166,-390,624,-200,-1658,1690,5288,185,-1425,-2868,7988,-592,3291,-220,4257,-388,1633,-4211,7260,-535,1384,-2702,-3464,749,-1151,-4550,-3688,246,284,-1768,-2998,-7285,-1379,-1337,-688,-370,2978,-5991,1666,-3039,-3308,2150,876,-294,-1971,1923,5073,-5175,2722,3251,-1462,-3278,2028,-4113,2807,4492,1341,-139,3010,3454,1882,969,-84,877,-792,2249,-2117,-418,-551,-579,5278,2951,114,7211,2279,2968,1052,-921,4343,2258,-3129,-1556,-5781,696,-1751,982,679,-3889,-627,2558,-778,2880,2135,-1719,1246,2119,-442,-676,1569,3740,5742,2702,2210,2460,2189,3071,4155,-2291,-673,210,-3579,762,-1188,5737,1909,1427,3608,4038,1840,910,-304,2183,5615,-2156,3430,2048,5000,1211,2003,-6376,82,-3352,-822,-266,3020,-8100,-2362,-164,-2386,620,-2988,3994,-3117,4572,-957,-1026,52,3442,-2661,-58,5458,-1208,584,784,-389,-2531,29,-1424,-2362,4536,-371,-2138,-2529,1785,1871,3256,676,-643,-725,-1011,-141,1994,-449,1155,1951,-11,4147,2270,2749,2785,-4865,-1978,600,-1984,-2631,3339,6596,3200,-179,-712,512,2856,1763,706,-3515,-2196,1340,-1718,554,4016,2707,-5878,1340,-1406,-5146,-797,4072,-3022,-4079,3532,1901,-56,-916,1718,4653,910,296,1735,-102,2575,-5161,480,3286,508,2763,-1940,-3920,377,766,-3339,-3195,-2335,-3266,312,-3110,419,3129,1048,-2142,-4055,-1458,-451,-1826,-6430,-1085,4340,2517,-3884,-3100,-293,1386,-1960,-456,-1943,-770,2812,-3161,1759,961,2639,3845,-3713,-531,717,-3928,-485,5146,6259,-1474,-4960,1607,-8432,-525,-1304,4213,878,-861,-1877,1025,590,-5854,-2653,668,2700,-2973,-4133,2780,3559};
    Wh[87]='{1759,967,1506,-2121,-711,4704,-4001,-3125,1734,-2788,798,-363,-2093,1651,3420,911,-4794,-5664,2258,-336,1018,559,-5708,-823,-451,7133,3388,614,4267,81,-622,1060,-1571,-899,4299,-1584,2536,1397,-482,-3496,852,-581,4919,-3212,4873,3032,563,68,2937,-836,1804,-3227,-4313,-698,-723,-1998,-2067,316,-691,7617,-5644,582,-3334,531,3762,4667,3842,-576,-1184,877,-2695,-4067,-230,5869,-545,-3786,163,5297,3137,286,-634,-4560,6352,-1712,983,-381,-1296,-2141,-1335,2785,6054,-756,-1,-3059,-2446,-2152,-1578,3068,-2746,1233,3554,1738,494,-288,469,-4665,-6025,-657,-4409,-3500,2469,-2634,1229,-2800,2514,4580,2009,-1779,-5131,444,911,8037,7553,-1063,-5493,-6215,3303,-789,-992,1578,910,834,2215,-1690,1711,4440,419,2731,-1818,1662,-1958,1560,310,1528,163,3686,6040,-3491,-2030,-1083,2229,1872,2390,5415,2253,1319,1519,-3513,-2265,10947,-3784,6367,-1352,-2465,2556,-2191,1301,-2407,-867,6684,3305,7475,-2415,-3322,3803,-2124,2023,-240,-2253,-1662,-2343,-1513,-3005,-426,5209,2890,1423,-3369,2700,231,2683,-1862,664,-2218,-2731,4929,391,289,-5961,1687,3085,-1027,-1320,-3046,-938,-966,528,1939,548,-345,-1479,-695,-1398,-3967,-480,-5493,1625,5312,1336,503,650,-1754,-586,1118,-4775,-1302,2048,95,486,1572,4072,379,3635,485,-3688,1347,-2810,3015,-4226,-908,-3627,-3623,2196,3969,-2237,-1500,5781,1602,-33,2042,-1911,-917,-1422,-7426,-508,-3354,-2396,-6850,-597,-4338,7949,-1857,4157,2165,-218,-148,189,-65,2385,1151,-1419,-939,3959,-1685,4707,2619,4628,-258,2890,6064,281,2445,4436,-2822,3205,3618,-848,4582,3342,-3828,-2449,-1802,131,-1868,1716,-183,3359,2644,-3657,2746,186,5786,102,4409,-1258,4245,3405,-4396,510,3676,-2839,1779,-4465,1660,4760,-2239,5839,178,6083,-2622,-2158,-890,-1994,-1894,-5576,3217,-6113,-1781,5327,3225,3315,3732,4414,2998,-3977,128,-422,-1264,1062,-2739,1594,6162,1730,-719,5141,-4802,5112,-369,5937,-3356,6816,2805,-2841,1927,-4138,-2575,3061,5498,10214,2939,-407,-487,-211,-4868,-205,672,-563,4572,-1928,-1254,-3776,3508,430,3090,1018,2924,-246,-2260,2401,-1862,1968,1978,2949,1911,-3901,4958,-176,2158,-3813,-2468,1268,110,-7919,-5224,-4682,92,-1018,114,-1534,-97};
    Wh[88]='{2714,353,152,-3442,466,2019,1462,-1127,-2683,-1217,1236,1879,-7158,1915,2702,847,1658,1121,-346,1049,-587,1889,-2462,1575,-351,-673,-1755,944,-2385,-2670,-593,1772,2644,4567,-4038,-1336,-1287,-4050,977,-1162,-397,568,3786,-3139,519,-1589,-5083,185,-735,4416,-2333,2917,-1148,3234,-241,-1282,167,4826,-227,456,2011,4299,-1625,-2113,-3493,-4936,1076,667,-1804,-1033,6674,-1623,532,1635,-239,-3044,-92,3679,2729,-1495,-750,3,-6337,1774,2702,1735,2512,-1485,7919,1345,-679,4909,332,368,3566,-2310,892,2491,-207,1528,-1855,1612,1185,-2208,329,141,-1926,-1674,2983,2364,-2438,-1591,-5283,-2443,1241,7163,1594,-3339,3820,-5727,356,-8017,1444,806,-2340,4262,71,4201,-89,-2316,1262,566,-2478,-2084,7153,-531,5371,-5927,-1129,2214,298,-254,385,-2197,2486,-3215,767,1180,-603,-1811,1466,2011,-2705,-5581,-2656,4479,-4870,-297,-715,12343,-3615,-2939,1062,-5537,725,-2937,-2185,1671,1754,2130,4328,1922,3886,589,-302,416,-537,618,-2288,2739,-1196,3093,3088,2827,-4057,1004,-390,1995,-4448,-4240,1499,640,2900,-1413,-2015,568,-3864,1290,145,-242,-1172,5034,-684,2800,-869,2912,-1522,5200,2305,502,-947,2062,2612,-2958,3144,2937,3312,-646,-2478,2753,3244,876,587,-2626,3413,1676,3430,-188,269,2897,6660,-3395,1894,1444,-1013,1384,599,526,-1973,-415,3254,-1156,-2966,-1469,-1372,-2264,1229,1298,-1518,5,2152,-2968,-1166,4624,-1411,-1280,1459,2636,3608,-4438,322,-2331,1744,-2465,-1336,-47,5429,1683,-620,-3527,-3864,-2351,-1138,1361,774,4604,-930,552,-1767,-2427,74,-2075,54,-3156,-1884,1153,-1474,532,2015,822,-2288,1091,2208,-2531,4118,2199,-188,-2148,3850,-1295,1132,3378,556,1608,-631,2258,-3305,2912,-240,5258,117,3923,1078,2337,-2114,-2507,-7275,1927,3459,-2707,-1422,-1232,-3405,-4577,3127,-228,-1437,2390,-8125,-1671,3679,1984,4201,455,5083,383,1488,-1953,118,-1798,-1091,-1346,-1787,-312,2093,-1372,19,-2700,1093,385,-3674,2009,1821,-795,1702,2482,1315,-517,1059,4541,4802,2429,3303,2322,-3764,-785,-739,1630,-192,1337,4975,2047,-304,-3168,3386,3894,795,-197,-1148,2663,-3903,5942,1250,3398,4091,-3808,-4089,1265,6132,-5253,233,-226,-465,-769,-1271,1697,2817,-2498,1622,-380};
    Wh[89]='{4338,1990,-2924,1013,-909,2098,-4758,-4350,-2093,-2531,913,-1522,439,-1662,-1683,-3833,-446,3691,-591,-949,1524,-1132,-4865,-1513,-3359,1212,834,257,900,2414,903,7919,-6386,-1710,3420,-1041,-303,1041,4060,-3498,-1657,-1993,10683,-1798,-3757,-2220,-3818,4082,526,3103,-3117,-3281,4558,3049,3549,8007,-29,5434,1621,4279,1383,196,671,458,3100,740,-3217,-4621,-339,1900,3193,3105,-1004,-3083,-3605,575,-4924,-3103,4533,-377,-1353,-1069,-2294,399,-486,-1853,-2797,-1212,-3095,-2531,-1735,-3312,-2132,-2666,-3676,-571,-7211,2878,-1260,-4177,-728,-7480,-6416,6186,-1805,-2778,3837,4985,-6342,1446,99,-6000,2875,1837,-1427,4511,119,9072,2438,-1842,3952,-206,-2254,1940,-5053,-1569,-7290,-1350,-566,-14589,-700,1647,446,2802,2941,1959,5078,1346,5947,-2019,4416,-3364,8300,-1282,316,-895,-6059,7792,-368,-749,3283,-1391,3457,562,-3112,14121,4633,-6499,1072,965,3212,-30,3403,-4726,1569,-2541,-2573,-2832,-5161,6225,-1939,-3469,-1135,-1004,-673,1579,-3867,70,-4638,3747,-4277,8779,-5717,3354,8388,999,-7709,1505,1407,1110,6708,9687,-3549,1278,-3613,-1101,-1198,-1639,-1733,-325,-1293,-2512,-401,476,-1843,-157,1663,9711,2297,-3076,-2629,-3120,-2115,1451,-2083,-109,-4777,-8857,-1250,-1335,2219,-3869,-1334,523,-4287,983,1563,1939,-2022,2849,-1451,1604,-221,-1339,-1095,435,-5693,1734,5268,-800,6445,4843,1707,4792,3962,-698,2875,988,4995,-3981,6337,342,-3259,4182,2463,6816,2763,1453,-725,-3017,-9106,-946,9409,221,-2558,2783,1473,-192,1892,1475,-335,2958,-3425,3320,-3063,-4479,-2426,-502,-4645,2502,-4709,-1604,202,182,-1132,-537,4331,-2707,-1309,3115,-10791,6777,7182,-3662,-8281,331,1445,-3991,7729,-3361,-6176,-441,-9980,1856,2700,-7348,682,-531,1098,-2849,1558,-8071,1115,430,-3576,-2261,4592,1079,-10068,1259,-6582,-1707,2822,-1268,-2656,4960,-1256,-971,716,432,-7021,3696,2753,2678,-5214,3811,-7172,2648,3955,-163,239,4821,4448,5532,757,3151,-4084,-1216,3391,718,4555,3891,-529,2309,-1072,-1834,-2639,-9936,-8525,-856,2910,3437,3862,-2199,-1987,3273,-997,-4667,-3417,-1614,7646,-467,-2348,-3793,-3205,1798,4145,3247,-4079,951,2424,-1773,5336,4333,-3391,-322,756,-4118,-3640,9501,-10742,3706,-293,-3681,-1918,-5839,-3271,3251,2385,-3017};
    Wh[90]='{-1010,466,-256,3769,-1439,-1043,3210,-1049,-1068,1256,4567,1824,1064,2915,-995,5244,4912,4150,2612,-3146,1838,-2055,-295,1541,-2366,4924,1259,57,144,6474,-20,4780,2990,1656,3891,1239,1655,-118,208,3955,11,5000,-1596,1655,2045,2573,960,-3588,-102,-3957,693,1040,-2183,2326,-2912,5737,2462,-2885,4016,8247,-1274,3474,-2110,-1683,278,1065,3039,9096,1726,2675,1066,3662,4543,157,1095,-2741,4748,-955,-2363,1528,581,386,8222,3427,177,-120,166,5034,1342,4050,-416,-117,2661,-3867,5258,5541,-1205,7749,3503,1718,-3283,-3928,-1820,7045,-6748,-787,806,6025,1224,5263,405,3276,2038,-1025,-839,1815,1717,-5771,1818,-3718,-4265,-5537,-3203,2009,-606,-392,2177,-2083,-3105,-12324,-1894,1997,3310,-3188,-4899,2668,1475,-2604,3408,1840,-828,2473,-3146,-1586,49,-1726,-3740,2407,6445,-820,-4663,839,-642,408,2196,3984,-552,-1046,6030,8974,554,-737,396,791,-1132,3325,-2512,2854,1161,-516,-168,1499,-1347,-1245,-394,1148,-7646,4196,-2612,2827,-2016,2656,-1945,556,3762,-1899,2003,-1337,-6572,1877,-1207,-4755,4479,-190,2729,-2145,-3857,787,-5883,-2215,3881,3986,-1069,-2209,-1943,-1431,2077,3837,-4890,5605,4245,1160,4689,-4453,760,2408,-3830,2261,2729,-3039,-635,1148,108,-1850,-2471,4548,1802,2358,-1206,-3134,-1727,-942,474,-4555,-1263,-970,24,1251,4118,1318,-357,4694,-908,-2,84,-1212,-7338,-111,5537,-1535,4206,1384,1517,231,-3425,2602,-21,3286,1490,-6762,-6215,5961,2371,6777,-2844,2070,3349,290,3483,-40,800,-9716,3769,4628,6835,-3142,1398,-248,3840,5888,-111,-878,4516,9008,-1351,-13,338,1564,584,-690,-399,-179,3300,-2322,-4650,3784,4772,298,4257,-2629,2861,-6538,-1087,588,-3308,10166,2722,207,-1828,1992,812,5209,2257,-807,-3298,-197,-2360,2988,-605,4785,374,1638,3015,222,-1223,1741,5327,2971,3732,7480,1177,-2369,2192,1982,-1057,2145,-150,6035,530,-2565,301,3771,2844,4938,2995,285,-5478,2145,7192,1624,92,-253,770,-2247,397,-3479,6215,-689,-2392,-117,4145,4807,-1206,311,-2036,4978,-484,-2790,4511,2121,5566,-567,2397,1903,3544,1520,-1761,-601,3715,1409,2039,7905,4333,-771,5585,6,897,3903,1566,7138,-7114,-3044,2626,906,4326,-1684,-2907,194,6430,-3427};
    Wh[91]='{-1303,-4248,3586,-3193,326,1168,-5185,2680,-2597,1248,-2939,-1071,-1551,681,635,-96,166,-5253,-230,-5312,3334,-1647,1322,-663,2032,-1106,-480,135,-13906,-1311,6362,-7685,932,-588,4418,1258,1463,669,-176,10791,-1557,-8945,-3635,684,-2216,-177,2924,867,-504,1055,-2106,-17,5078,4260,-4738,1557,-2086,5961,1105,-7041,737,5668,2272,-3737,2235,-1915,573,2092,2149,4868,-872,-2775,5009,-2976,7221,3698,1120,5541,1333,-4645,-54,5419,-1204,-557,1166,-4291,153,1028,-547,-1353,-6958,-1470,2504,2254,-1099,-525,439,-9340,-4746,2176,-1019,-4460,-2481,7509,-2026,-1934,-3381,2639,-10380,11406,-2464,3325,1380,3986,23,6328,-9218,-14091,-13525,-18105,698,7402,997,-4506,-7631,-991,7607,3330,-1435,-3435,772,707,-1956,7382,-2783,-3527,-5693,-508,40,-2067,-6352,-553,-6508,30,-4580,1103,-5273,771,-6904,67,-1853,-3806,2019,-1655,4121,3857,-4501,-785,297,14707,-8579,-4199,261,-1365,-1826,7656,1972,885,2023,-548,994,2854,6918,5561,1193,-2841,281,-1214,-158,1306,392,-3962,5698,-1542,115,-3164,-1706,-3090,-6782,-3867,-1649,-5927,520,2055,1909,-13906,-9575,1518,389,-936,-3452,3750,1364,6123,4113,1987,4248,1245,-495,-884,10341,2783,7041,286,712,3850,-831,1467,2257,1257,2905,-6547,-5385,2985,-988,-3686,-4543,3422,543,6523,531,1705,471,-3806,5009,6772,754,2027,-1238,-1839,-6337,4667,3181,3562,-175,-2932,-2188,6494,3295,-1486,6914,69,246,-4130,4011,-583,6816,3107,3447,13525,5371,491,-1287,762,1354,4711,5766,4758,1904,321,-2854,-5458,-505,2124,3937,4133,-547,3303,1524,3388,382,-454,3347,-5590,3605,-3310,4326,955,-12089,-5869,-9746,-8056,550,5380,-12,8081,-1143,4394,3876,-1801,3825,-88,5458,-95,4187,8535,3259,341,844,3615,535,935,1295,2448,-4167,838,-2888,-366,5688,-6567,-9663,-1791,-4772,565,-2276,-2578,-4440,-1383,3684,-1763,-1345,337,-2846,511,-747,-3110,-3437,4792,-3581,3491,-2423,-2294,1125,725,29,-2690,-3002,948,-9926,-568,1209,-4768,316,1313,-7119,-3466,516,9355,1109,-3408,4628,1850,3007,-5229,2756,-5322,-907,-4379,-1542,2222,560,-3017,-2028,-1607,374,321,-8823,1596,-1899,-493,-3239,-7607,-429,1149,-561,4150,7480,2985,-3427,-2218,-3276,3085,4272,-1489,9096,5278,549,2956,2512,831};
    Wh[92]='{-1851,1235,-203,2871,-133,1516,-491,-3330,-1760,-2517,1693,-155,388,1352,2222,871,4396,-867,2941,229,419,2196,-4333,-133,1331,1446,1362,1029,5434,111,-1329,1285,4536,1450,1193,836,-775,1877,-1143,1057,-1455,1467,-1005,6054,-1361,3427,1606,-597,5537,965,8203,-782,-2379,1816,6743,-5146,-472,-5019,-1575,-2332,-747,4484,842,2766,4597,-2661,1218,4545,-4023,-2983,1001,-4345,-977,567,1489,7094,7504,3994,-1683,-266,1065,2502,-632,2382,-2432,3051,-265,-4628,2834,-2160,-822,-2570,-850,2800,-817,-570,-1307,-662,2844,-1810,2727,-4299,615,-742,-580,-1845,4980,3315,17265,1176,194,-2376,3041,-1545,-4785,-1550,-654,4921,-4265,3291,-206,489,3295,-2702,6494,-4140,-4162,2937,1849,2937,-3505,1619,-3354,-1654,-2897,-1235,-227,1431,-474,-4055,695,-3281,-459,1574,-2697,-2138,103,3984,-56,1440,-433,-3161,-444,173,-3557,2432,5341,-2344,-138,-41,-5385,-1210,5263,8515,-5561,-260,3000,1518,-3398,780,1708,-2343,6577,-5097,-2612,5478,-1868,-5322,-1374,2851,-1088,3244,57,-709,-1490,-278,832,-3063,4677,-3535,-3586,3632,-1564,-2819,-3984,850,-1912,-473,-5180,-6845,1188,-1165,-3066,4890,2426,808,-2338,-5244,-1579,-1206,933,-3461,3852,-552,-1419,-2846,300,3967,-2990,-665,1468,-1590,-4262,-7553,6137,6206,2834,2384,-656,3532,747,-508,2199,-3249,-6552,-3476,1501,-592,-3103,1292,6645,2551,608,-5815,2661,4731,2731,622,-655,-1406,768,-7290,-1240,-3417,-599,1859,-2227,1765,4257,685,3806,1364,-10292,-855,-4401,-2526,61,182,-7265,2413,-1206,5000,4831,723,-4394,-2008,-1923,-1423,-639,1638,-1923,2237,2810,-3415,1180,424,313,27,-2341,2343,-4909,-4177,3903,1248,654,5083,-1610,156,1828,988,-4309,290,-3520,2880,1597,943,1844,-3894,1226,-3381,-2258,6064,-1536,1601,1564,5395,1352,-847,2332,5268,1292,-2487,-1628,961,746,4069,-1026,4248,-4396,-1157,5131,2410,-1284,572,2319,1205,-59,1037,-3647,3669,802,3027,-1101,-3874,-795,-1478,-4091,-478,5854,1555,-2585,5336,3513,1524,1735,-1691,1340,8540,-8676,5263,-3393,8032,2868,7231,-7631,2346,-897,1110,-4921,-4855,707,-281,4533,-3095,738,1936,-960,2871,-3310,1599,-4458,1636,3889,-2519,-3361,-4731,819,-4794,4575,-3554,-2277,-3552,-2785,3464,-874,4643,830,-4260,3134,-899};
    Wh[93]='{-1640,-1614,-1881,-128,-4182,3315,-5834,922,-2595,-3334,-5390,5180,2844,-152,-3691,5048,-12382,-974,-3076,-3374,-2714,-3725,352,-4680,-3688,-4650,-575,-2293,-8666,-4309,-4621,-9980,-12812,-3061,8789,-1188,-3134,-4536,5156,-331,2452,807,38,4536,-6484,-8681,-848,-4980,-4028,6381,1811,-10078,-1834,-2863,-5278,-3168,-3752,6269,-6411,18183,3867,920,-4523,-3483,-5698,-4631,-1693,-4577,476,1884,6118,2308,-3012,-9311,-5600,-3764,5957,-5590,2087,-2521,-101,-7373,-5166,-1337,534,-2403,648,-3239,1721,3842,-2834,-11542,-6328,-5541,-5336,-892,2897,-6381,-5336,-3229,-6191,-3881,-5766,5244,-1424,-4169,-3151,-10126,848,-4379,-2927,-3027,3105,2846,-4091,5141,-7607,-1674,243,3703,5219,4907,1712,-2298,-1931,625,-8291,5947,4326,9892,3017,2832,-824,3625,-3200,-194,-7856,-826,-748,2,-1256,3376,-6513,-2386,-352,-4167,-3999,-509,-11503,851,2232,1552,2929,-1849,-1768,-7441,-10839,-3452,-8476,-31289,4555,2963,5371,-921,1527,-681,197,2413,-5327,2182,-2423,-2866,4060,2556,3591,1976,-1220,-3718,-89,870,8549,10859,4494,4765,6972,-567,6469,2790,902,2188,-2575,345,-2985,-232,5390,4233,6767,-3144,-5083,272,-2371,3168,3400,7968,-3435,3120,5244,5004,-5590,-6982,4609,-10878,-7216,-4001,-1064,4177,2910,-2121,-5239,1319,452,-10117,-643,-6069,-4843,-9785,-3645,-2988,4665,3161,-3811,9389,334,1896,4831,-986,-3630,-3630,-2517,2073,3469,7832,1971,-7539,1666,1868,-4704,-988,-1840,-3447,-2612,-3281,388,992,293,4899,-989,894,-1712,-6376,-6987,-451,4904,-164,-2152,1865,2196,-2993,1429,1191,-1105,7695,-9355,-183,-3029,1428,-8500,2150,-841,2927,-2644,2329,5883,9223,817,-3181,-897,3815,-7260,2866,-2724,12021,-3908,5385,-2976,698,-2697,1506,-2048,11132,-9296,6596,-9521,-2587,-751,-5043,4189,-901,-5537,-3796,-8081,-7441,-1012,-1949,988,7661,9404,-2714,-12714,-10224,-10234,-11660,-2663,-406,-215,331,-2998,-2104,875,-586,-6801,3605,-1147,-597,-8549,5380,-1035,-8349,-2885,7548,1124,5395,2166,13554,524,-615,-1024,977,-7553,1234,9882,7983,-5000,4611,-3706,1235,-5278,-8481,-1820,-249,-508,6040,-117,-3728,3422,-7543,-1329,4497,-7045,2565,720,5541,-8027,-588,-8813,4929,-309,1638,1160,-1282,-372,3598,728,6972,-5742,3527,-8544,-1152,-5981,2398,2117,-27,-4011,10166,2712,3066,-4599,4799,-6723,4074};
    Wh[94]='{-445,-4970,173,2902,-1522,-68,-1712,-3845,6635,3471,1616,2322,-2346,-101,-6938,-386,-7075,-250,-208,1866,37,6137,3654,2415,244,-409,1677,112,4201,850,3334,1591,-7656,4294,-458,1302,-3498,-2489,-4272,2369,1231,-1302,-1028,-718,-231,-4206,1973,2873,-2047,-1542,7060,139,-5288,2371,1861,-2934,342,-1226,2406,1140,4294,-2464,-2551,4448,993,5405,-2210,3684,-263,-227,-3903,-6591,-587,-2756,-710,1751,-2897,2208,-3459,3078,2998,-7421,2036,54,4057,-2912,-2851,1679,1068,706,-462,6635,-636,1058,-5288,395,1308,878,-4711,2073,-2006,9277,3698,-16386,2004,907,-2482,5688,10273,-5991,-92,-4379,12666,-7973,5830,2081,1318,5517,-3249,8364,-3068,2714,-11826,-12324,737,6176,-3830,3786,4892,-6313,-1829,1000,8623,-12744,837,645,-1184,3811,2092,1904,4682,-225,7602,-1940,1713,-10869,7797,-10234,2697,-3583,-3398,-4562,-10078,2504,-2260,-7060,-8901,-5581,-2109,-12246,11074,-1915,-95,-5209,2805,-4194,1473,-3051,1890,-5585,4763,1154,-2479,-5786,-3264,678,2854,2683,5947,-2678,2061,-6254,-183,1519,-439,376,-783,732,14189,877,-4926,-6801,-8339,1777,1334,7456,-3562,3562,-3493,1909,166,-84,-3891,5747,-4101,-451,-6586,-3750,-4409,3317,-5854,-8056,3173,4311,-419,6787,-5615,-6767,-2410,8535,-677,5742,-237,-6225,4140,6240,3842,318,1754,-2604,-332,-4934,1335,1069,-8056,-1713,-2822,-5161,-1794,3649,-4167,1833,1737,-7094,-1895,-1335,-4814,-2066,-485,2106,-1507,-2832,365,1798,2243,-2103,-4682,1021,-2254,-12050,3725,-2325,3454,63,2136,-1219,-4218,-11416,-267,-503,-684,6840,-2995,1169,2751,-5751,-2203,-342,1188,4057,-3547,-3935,-1632,3603,-115,-7460,-5771,-7202,-3876,-1238,3842,-7973,-4843,-3911,4125,-11650,-3388,-2199,-5581,5927,171,-7456,-41,-406,-1785,-2558,2285,4479,5361,4675,-5126,-1926,-1030,3659,-3256,-6118,4826,806,-7231,-2006,5258,10791,-4094,849,3144,3037,4201,2310,-1228,1585,3098,5400,-7558,-1341,57,4033,-3850,-6513,-2036,-3383,158,-3430,-646,-5878,-2387,3623,6225,513,1943,-1790,-1926,-548,-3994,1326,8330,4213,-911,-2017,4125,5605,6181,-7519,-2413,7275,-1638,1513,-2712,2279,-1408,-431,2683,4128,-508,-1896,-2465,-5351,5454,-194,21,9384,1242,6308,-3505,894,-4599,-3281,-3176,-3479,785,7211,3186,2875,-4091,2856,1851,-4870,4003,3393,-4406,1495};
    Wh[95]='{-239,-5756,2705,-4116,330,-1119,-5161,-3032,5585,1517,-1752,1511,-419,-7739,-4201,-2827,-3710,498,-172,939,193,-2144,6206,-2119,-1385,2734,-3176,1524,-1751,1562,-2597,-623,-5029,1676,-5078,323,-347,-2263,534,-3110,-7197,-3251,-7827,87,725,-5541,-3105,1684,-5141,-490,-7548,1034,2563,-689,4370,-11289,-2225,-1540,-4145,-4799,-1285,-2973,-2963,6962,-3215,-641,-888,1557,1250,405,1027,5576,-1357,3901,296,-2827,-5922,3889,-3906,2288,988,-5444,-709,934,4777,-5532,90,-3154,-2335,3652,-1477,-4025,-1038,3361,2269,-1423,-2868,3012,576,-5698,-2321,-716,-3793,2617,-192,1411,1651,1381,-3405,2636,-4587,3408,-6328,-1003,-3754,-982,-2314,1342,1645,81,-3134,-2355,4189,-1155,-5083,-3818,6879,-2429,7290,-1614,1040,49,-2504,935,-1074,-2956,-6396,2028,415,-847,3569,-376,4301,1206,-2169,-729,-26,-764,1809,1833,-2078,2246,-380,-3327,-7343,5454,-1850,-2707,3386,-4682,-4887,-5288,359,-3022,-5156,1499,2875,3928,-858,-401,773,-1885,4792,-207,1143,-1140,1536,4282,1121,102,-2344,5258,-4282,4885,1071,-1994,-3974,-253,8608,-2349,1324,4113,4868,3674,-2326,-5610,1418,-1142,3920,-1168,2705,4589,4377,-2059,-3808,-1313,2822,885,-235,-3920,-5527,2592,-3542,-2563,3676,-290,812,-7788,5200,1130,933,4211,5380,-830,-7954,1074,-1879,2231,-2174,391,20,-1112,79,703,1347,-2580,1175,2153,6196,219,1669,4509,-10468,4741,-3022,-928,-2310,-3200,4084,-4157,-1789,3576,-2885,-664,-4670,-4113,374,106,-1121,5864,-1483,1594,-4638,1855,1391,781,-6015,317,2370,1994,-3122,-78,-1362,855,1185,-3203,3635,1546,-2939,1506,-5703,-625,2731,6015,2041,-3530,2678,523,499,-3476,1090,6093,-1239,7324,2222,-2717,3710,-1937,1824,1634,2280,-2346,-1146,-5327,-3908,-5444,2078,792,-1071,-6274,4782,-672,-738,-4086,1623,-2440,2304,-1013,2325,715,-1159,-2445,2141,-889,-2895,3303,1329,-970,1934,997,-2680,-5161,703,1056,2322,-4008,-1638,-5434,423,3779,-4650,1910,-4787,1348,3647,-2529,-356,3986,1839,-3159,-4428,2044,-1390,429,2034,-1591,3020,-4873,163,-5327,-915,164,162,-4794,-2169,-5029,-4526,3374,-631,2119,1265,-2402,-1237,-3562,-9624,3706,-819,942,-1256,4038,-4641,-2714,-59,-1822,-1040,1315,3188,56,314,-2636,-1566,2078,-3688,-1312,2247,4885,-816,-2988,-177,-2132};
    Wh[96]='{-159,-3730,-986,-4277,-1562,1226,-1132,619,-4331,-267,-3281,-662,-7,-702,1325,-3247,-3015,574,569,-2702,-1877,-2250,2010,-1441,493,-2204,-3186,-1650,1885,-306,-819,-305,-1104,1058,322,142,697,2264,-704,-4572,1632,-3342,2399,-3942,824,852,464,-2780,791,434,2414,-1170,-4338,2814,1560,-639,283,580,-2744,-1464,-335,-2041,1339,-7172,-975,-2357,144,-5112,2023,-698,3454,480,-2792,-5957,-847,-4035,260,-4919,-850,-3195,2418,-4260,-4047,1650,191,-3784,1237,-552,-5439,2147,-1862,-8911,-3356,1514,-5400,-2475,2502,-2369,-1730,-494,2973,-71,-4069,-4770,5405,-2958,-2893,-4020,-1002,770,10,6523,5097,-38,-4145,822,174,1956,-4145,-3571,3955,3769,2270,-2241,3591,-3146,-279,139,2656,522,3364,510,-99,653,6787,-4367,-6884,3037,-8364,3288,-1940,1423,2233,1693,-4523,3859,571,3273,-9116,2822,-953,-60,88,-563,-4416,-3142,3276,-1458,1922,-6811,3032,-704,-1599,3151,1608,792,-624,-504,-1175,4484,2049,-3256,-4904,-3376,-1149,2161,448,-2106,1232,-4890,895,-4631,-1934,3928,393,780,-8325,-3701,-2308,7954,-168,-1106,-1281,4492,543,33,1235,-1217,-1750,3217,-1196,-2714,-525,265,-2286,905,2624,-1911,775,-2836,517,-2561,-7431,4946,-2301,637,2578,5688,908,-2998,360,-554,-1430,1149,636,-773,17,908,-129,-3305,-1137,-6508,-4333,638,-239,1789,-77,808,-1189,-1800,-1442,-2712,946,-879,3046,1026,2773,702,-4245,214,-2575,-991,-3679,-613,-134,-2252,3657,2491,-345,5605,541,2070,-3598,-1802,-1039,2858,-1569,446,-372,3159,-5302,952,3317,94,-1436,4216,2604,54,-2159,-1121,-3281,-3684,-3017,470,1918,3278,683,-4289,-1181,4282,1452,4465,-3227,-1046,-2770,-3889,-3242,-1566,-852,3808,-2502,2192,-2761,-752,-1203,-6347,-1225,-6030,-1457,-4497,-1369,-4785,-3024,-4074,-1005,-9082,1304,-158,1271,-9174,-886,-2636,-3676,-1628,3488,-2888,-4965,3051,305,657,-3845,-762,-5800,2988,162,-1506,4248,-5297,2011,310,2332,1113,91,-6098,1922,-1290,7851,-721,-9941,2536,2785,-2888,989,1968,5229,1749,1760,-755,4169,-5019,-1053,-1856,-2478,-4318,5405,1032,-1678,300,-1021,3356,-3044,-1129,-346,3232,-2128,-3283,2668,3200,138,-397,-4272,3935,-2056,271,-4936,659,-1303,-2337,-2692,-5302,1241,-4372,720,-143,480,3854,11835,-1016,-2498,1826};
    Wh[97]='{2137,767,-653,-2775,1867,1445,-5009,-6166,-847,3520,-914,-2416,2868,1164,-2902,4665,7446,6440,-3569,2783,1365,-987,3122,1437,-617,-1849,3979,1949,303,3435,-264,-282,1035,-3066,5034,711,2247,-1685,-2304,2452,-107,10,-6943,-6840,-186,-1390,-2993,-6782,-1921,1589,1301,-485,-3803,3500,596,-2343,1558,-94,-736,13300,-1655,-2915,-5043,2805,2413,518,-925,-1545,2108,-2614,1270,-92,3095,-4348,-1583,4143,-393,3098,422,5356,-4255,-12812,-2558,-2060,256,3666,-872,-542,1633,5288,-2917,4726,-540,-5273,-9272,-574,-2292,-286,-2423,-3903,-10615,-1218,908,-3896,491,-1943,4753,-3100,1205,-2941,738,-1065,-3547,-1335,-3193,-3750,3200,4699,7104,7973,783,1194,3903,5766,-8452,-4372,3696,4699,2102,2971,-5058,-4323,-4665,4123,-6972,5429,-108,-4829,3896,-5629,12109,-1213,-1701,-6235,853,-7885,-194,-10009,298,-2230,2469,-4436,2995,-7065,-1147,-1993,-266,-1207,2175,1222,13291,-2482,1453,-10371,-1473,2229,994,3278,2292,-2233,-3947,3432,-5073,-8432,-2330,4750,-3469,-882,-881,-509,-2108,1937,-4565,-299,1583,3205,2719,-3798,13154,4709,1964,1563,-3635,-3151,-1528,-4782,-2137,4116,1369,-2381,-335,2880,1799,2568,-2012,764,5078,-2203,-6191,4699,3300,-869,5712,-6406,3486,2113,-2192,-4809,-1632,1851,3579,1729,1948,995,3276,1088,-595,1948,-897,1931,-3298,-2841,5781,-1771,495,-7006,-980,-407,-223,-2702,2165,-588,551,5336,-2541,889,601,2873,231,-4948,-4,1953,2167,4318,1884,992,2448,3471,2226,-4782,-1412,8242,6381,-1212,-3078,0,-2539,2978,2247,-3129,-1896,-3283,-2592,6010,-704,-1012,7758,-1951,3723,-3037,-2709,-1488,8955,3803,2250,3122,-1875,-2248,5170,3044,-4423,11904,-1356,-2785,-82,-5029,3688,-1429,1228,3547,-1695,-628,-1262,-2937,1665,-118,-3613,-2427,-886,673,3574,-2624,1278,-828,251,150,-7451,3120,-3552,-2902,52,3281,3049,3198,-240,321,3903,435,3479,4104,-1534,447,-4709,2416,451,2912,-1450,-4177,2727,1766,2868,6123,-564,1495,1695,6943,-5908,8168,6318,-17,3693,2481,-4360,2432,-863,-589,12587,-5932,-3989,5986,-6074,5761,-4753,4265,3452,2644,-6855,2563,-7622,-2958,2734,5097,3391,-4497,684,-608,3588,1895,-1711,1530,-1956,60,-2275,1424,5356,-6230,1000,-1719,6445,-3666,-7026,-2481,-1442,-4946,-575,-4819,-8481,4943,1614,-984};
    Wh[98]='{4829,-2001,1375,-2736,-1259,886,-8310,-2558,2924,-1724,-12343,-6572,-855,-3244,4030,-5273,-3767,-3308,-4926,4675,480,623,-3483,-4853,419,4155,-4489,-103,-2785,3105,-275,-5375,-4240,-4833,2536,-2634,2958,-1508,-8515,-2658,-1494,-137,1955,-1746,2792,-1071,-2247,-5087,-783,1568,-8383,-3720,-75,513,1611,3059,-492,7509,-755,-3444,4411,4099,-2958,-3417,822,5312,-2731,-5781,2792,3898,7,-876,-1932,-4423,-1063,-6972,-4741,-2,5292,-1030,-4416,-1049,632,3332,1156,1434,-4199,1160,-3674,7905,-1788,-1408,3713,2912,-1401,-3395,6450,-2268,-4846,888,-3510,2436,-828,-4382,5263,266,-3737,3232,-1773,482,-361,3728,-6811,-349,3300,-1975,-3850,320,1777,-615,4536,-3454,-4123,-3872,-5864,-14453,3168,429,4592,-8066,5888,-3320,-2030,-2032,3173,-1771,8330,1789,-4521,78,-522,4340,4309,-552,2313,2451,3879,-2266,3249,2175,6420,2636,1800,-5219,-1223,3906,8994,-279,-95,-6191,2644,1452,-6611,-4401,1210,-4218,-2342,-3405,294,2495,2421,4096,2651,-1389,-386,-5976,-4187,6264,-3813,-1172,744,-2751,-2080,876,2663,2863,-5551,3139,5092,11162,1890,1718,-4570,2592,-1320,-5126,-5004,-6401,419,266,-493,6171,1250,1233,1754,1211,4978,668,-3862,316,-272,-2321,3601,3232,5190,-1359,2050,-2900,-4040,-1419,1383,-577,2575,7543,-733,6142,661,3559,4621,-2270,1756,-6640,-4384,2961,-3552,548,-5512,-1103,3261,-864,-497,-2230,-5131,2297,1155,1862,5283,-4291,3085,-2800,4018,1473,-3815,1313,-5351,-1635,4912,7397,-1981,4257,313,2077,6010,2744,-5834,4858,-1711,997,-1033,60,7158,8325,-1914,1060,-2702,4531,3779,1507,-1811,765,-4392,-5322,2109,-5371,-2448,1185,-2917,1071,2175,3525,1643,3664,2309,717,152,3388,-961,-191,5566,-3735,-795,1813,-3076,971,-1323,-3347,2163,-8222,-282,-2036,2553,-4672,905,-3754,11054,-3593,4223,-885,559,-992,1004,-2766,-241,348,-1156,2442,2646,-650,4531,-853,-2236,5317,-183,820,1293,2381,-3208,-1729,-905,3444,1409,-2578,3034,-5996,5268,-3198,6567,217,8295,-2658,-3867,2214,-6694,-1668,994,903,1868,3510,-2421,-1599,2241,1096,1171,517,2238,6186,-2802,4091,3771,-2397,-5307,1211,-858,-529,-4382,-4714,3767,1193,689,4223,-1634,-1520,5351,-8457,-1907,9252,-5234,2868,1418,2866,1784,-2766,3239,-6562,-1049,-3918,-438,-4501,2215,-687};
    Wh[99]='{2485,-4499,272,-1187,-1330,976,-268,-75,-7495,456,4,-4267,-4423,4475,-2697,659,-3386,378,-4489,2929,-960,-1336,-2641,-26,157,2225,-5263,-1008,-1827,-9218,3095,1143,-2150,1105,3867,2283,-3730,2398,1427,-5112,-2714,-1105,1981,-5717,2115,-3017,-3,-5087,-5517,391,-1262,-2937,-1800,1972,3537,-311,-4816,5366,-1511,2807,1446,903,-3222,-1370,-906,7036,137,899,3271,-2600,-2814,-1978,-5712,-4089,-2191,-6391,917,-1270,-949,-1221,1184,2303,5058,-4377,2414,4431,-3486,4479,-988,-85,-1348,1002,764,323,-1246,-4042,3154,-1580,-168,-5830,-10292,-798,-1522,7939,5810,1793,-1988,5336,-348,-3757,-3244,1379,-5371,1205,2414,-2932,-309,-729,-2205,5400,2489,3347,-2587,-4199,-1571,-7436,8017,1119,3383,-418,-979,1693,2158,-797,2592,-256,1403,-1802,-469,-70,-4658,1319,5942,1492,-925,3068,577,-4494,1330,-7749,795,5029,-7451,-2268,-4995,-4143,-3122,-1905,1992,-3334,-2214,1054,1716,-1061,5727,2196,2445,-5507,-754,-3395,-5024,2587,-12353,-4990,6723,-2302,-3613,-2709,-4475,-397,6132,-2320,-5107,888,-903,1286,-1245,-7407,-4184,3322,512,1486,1049,802,2819,-4721,4304,899,6303,-2626,-2064,-1428,5249,-4199,-3437,534,-452,159,-1752,-897,-3090,-5659,4443,-1246,1455,-44,2731,-420,-946,-2761,-273,-3457,-1329,1596,-588,-3537,-2939,-3603,-3186,-1463,1910,-3969,565,-944,-1184,3911,990,-2504,1676,-3530,512,3354,1105,-2702,-3037,-3796,-4184,-1041,-1621,1588,-3200,-136,5214,-3796,1771,-3249,28,6103,-3132,-1439,-2218,-1920,-3151,1013,179,-2822,-5634,-5698,-2305,921,413,5874,-2366,1126,-1805,-235,-1837,-437,2971,-4221,-1188,241,-3835,-8378,-5766,-7998,-2968,-7968,-3791,1888,-1510,-10419,-2354,-427,6645,-1700,-2543,-1080,101,-1423,-4890,626,5932,-2780,225,-1505,-2402,-2119,853,-4565,3991,-5483,2299,-5322,-5341,-502,1737,-390,-3334,-1877,-1098,2220,1043,4406,203,-2322,-2805,-2158,4272,-792,317,-1834,-4252,-1340,2883,1503,-1357,-6733,773,1729,-2661,-711,1555,-2971,1604,677,2695,-6586,3354,2156,1069,-9174,-3886,1231,4924,7866,1040,7080,5747,2712,-3249,-588,-3654,-2807,3933,-8657,-2768,2247,2012,-1687,-2612,3596,-3449,-4724,-4130,1898,4875,317,1350,1716,-3583,-2159,-252,-5664,-2050,6713,-2541,-5634,-7011,-3852,4138,2272,2739,1417,5932,2758,1944,-158,597,-1636};

    #10$display("EOF");
    #10$finish;
    end
    endmodule
    