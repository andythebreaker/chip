module mxv_TB;
  
  // Parameters
  localparam NUM_ROWS = 100;
  localparam NUM_COLS = 400;
  
  // Signals
  logic signed [31:0] matrix[NUM_ROWS][NUM_COLS];
  logic signed [31:0] vector[NUM_ROWS];
  logic signed [31:0] result;
  
  // Instantiate the DUT
  mxv dut (
    .matrix(matrix),
    .vector(vector),
    .result(result)
  );

  //dump-wave
    initial begin
        $fsdbDumpfile("mm.fsdb");
        $fsdbDumpvars("+all");
    end
  
  // Test stimulus
  initial begin
    //======================================
    matrix[0]='{32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0 };matrix[1]='{32'd0,32'd1,32'd2,32'd3,32'd4,32'd5,32'd6,32'd7,32'd8,32'd9,32'd10,32'd11,32'd12,32'd13,32'd14,32'd15,32'd16,32'd17,32'd18,32'd19,32'd20,32'd21,32'd22,32'd23,32'd24,32'd25,32'd26,32'd27,32'd28,32'd29,32'd30,32'd31,32'd32,32'd33,32'd34,32'd35,32'd36,32'd37,32'd38,32'd39,32'd40,32'd41,32'd42,32'd43,32'd44,32'd45,32'd46,32'd47,32'd48,32'd49,32'd50,32'd51,32'd52,32'd53,32'd54,32'd55,32'd56,32'd57,32'd58,32'd59,32'd60,32'd61,32'd62,32'd63,32'd64,32'd65,32'd66,32'd67,32'd68,32'd69,32'd70,32'd71,32'd72,32'd73,32'd74,32'd75,32'd76,32'd77,32'd78,32'd79,32'd80,32'd81,32'd82,32'd83,32'd84,32'd85,32'd86,32'd87,32'd88,32'd89,32'd90,32'd91,32'd92,32'd93,32'd94,32'd95,32'd96,32'd97,32'd98,32'd99,32'd100,32'd101,32'd102,32'd103,32'd104,32'd105,32'd106,32'd107,32'd108,32'd109,32'd110,32'd111,32'd112,32'd113,32'd114,32'd115,32'd116,32'd117,32'd118,32'd119,32'd120,32'd121,32'd122,32'd123,32'd124,32'd125,32'd126,32'd127,32'd128,32'd129,32'd130,32'd131,32'd132,32'd133,32'd134,32'd135,32'd136,32'd137,32'd138,32'd139,32'd140,32'd141,32'd142,32'd143,32'd144,32'd145,32'd146,32'd147,32'd148,32'd149,32'd150,32'd151,32'd152,32'd153,32'd154,32'd155,32'd156,32'd157,32'd158,32'd159,32'd160,32'd161,32'd162,32'd163,32'd164,32'd165,32'd166,32'd167,32'd168,32'd169,32'd170,32'd171,32'd172,32'd173,32'd174,32'd175,32'd176,32'd177,32'd178,32'd179,32'd180,32'd181,32'd182,32'd183,32'd184,32'd185,32'd186,32'd187,32'd188,32'd189,32'd190,32'd191,32'd192,32'd193,32'd194,32'd195,32'd196,32'd197,32'd198,32'd199,32'd200,32'd201,32'd202,32'd203,32'd204,32'd205,32'd206,32'd207,32'd208,32'd209,32'd210,32'd211,32'd212,32'd213,32'd214,32'd215,32'd216,32'd217,32'd218,32'd219,32'd220,32'd221,32'd222,32'd223,32'd224,32'd225,32'd226,32'd227,32'd228,32'd229,32'd230,32'd231,32'd232,32'd233,32'd234,32'd235,32'd236,32'd237,32'd238,32'd239,32'd240,32'd241,32'd242,32'd243,32'd244,32'd245,32'd246,32'd247,32'd248,32'd249,32'd250,32'd251,32'd252,32'd253,32'd254,32'd255,32'd256,32'd257,32'd258,32'd259,32'd260,32'd261,32'd262,32'd263,32'd264,32'd265,32'd266,32'd267,32'd268,32'd269,32'd270,32'd271,32'd272,32'd273,32'd274,32'd275,32'd276,32'd277,32'd278,32'd279,32'd280,32'd281,32'd282,32'd283,32'd284,32'd285,32'd286,32'd287,32'd288,32'd289,32'd290,32'd291,32'd292,32'd293,32'd294,32'd295,32'd296,32'd297,32'd298,32'd299,32'd300,32'd301,32'd302,32'd303,32'd304,32'd305,32'd306,32'd307,32'd308,32'd309,32'd310,32'd311,32'd312,32'd313,32'd314,32'd315,32'd316,32'd317,32'd318,32'd319,32'd320,32'd321,32'd322,32'd323,32'd324,32'd325,32'd326,32'd327,32'd328,32'd329,32'd330,32'd331,32'd332,32'd333,32'd334,32'd335,32'd336,32'd337,32'd338,32'd339,32'd340,32'd341,32'd342,32'd343,32'd344,32'd345,32'd346,32'd347,32'd348,32'd349,32'd350,32'd351,32'd352,32'd353,32'd354,32'd355,32'd356,32'd357,32'd358,32'd359,32'd360,32'd361,32'd362,32'd363,32'd364,32'd365,32'd366,32'd367,32'd368,32'd369,32'd370,32'd371,32'd372,32'd373,32'd374,32'd375,32'd376,32'd377,32'd378,32'd379,32'd380,32'd381,32'd382,32'd383,32'd384,32'd385,32'd386,32'd387,32'd388,32'd389,32'd390,32'd391,32'd392,32'd393,32'd394,32'd395,32'd396,32'd397,32'd398,32'd399 };matrix[2]='{32'd0,32'd2,32'd4,32'd6,32'd8,32'd10,32'd12,32'd14,32'd16,32'd18,32'd20,32'd22,32'd24,32'd26,32'd28,32'd30,32'd32,32'd34,32'd36,32'd38,32'd40,32'd42,32'd44,32'd46,32'd48,32'd50,32'd52,32'd54,32'd56,32'd58,32'd60,32'd62,32'd64,32'd66,32'd68,32'd70,32'd72,32'd74,32'd76,32'd78,32'd80,32'd82,32'd84,32'd86,32'd88,32'd90,32'd92,32'd94,32'd96,32'd98,32'd100,32'd102,32'd104,32'd106,32'd108,32'd110,32'd112,32'd114,32'd116,32'd118,32'd120,32'd122,32'd124,32'd126,32'd128,32'd130,32'd132,32'd134,32'd136,32'd138,32'd140,32'd142,32'd144,32'd146,32'd148,32'd150,32'd152,32'd154,32'd156,32'd158,32'd160,32'd162,32'd164,32'd166,32'd168,32'd170,32'd172,32'd174,32'd176,32'd178,32'd180,32'd182,32'd184,32'd186,32'd188,32'd190,32'd192,32'd194,32'd196,32'd198,32'd200,32'd202,32'd204,32'd206,32'd208,32'd210,32'd212,32'd214,32'd216,32'd218,32'd220,32'd222,32'd224,32'd226,32'd228,32'd230,32'd232,32'd234,32'd236,32'd238,32'd240,32'd242,32'd244,32'd246,32'd248,32'd250,32'd252,32'd254,32'd256,32'd258,32'd260,32'd262,32'd264,32'd266,32'd268,32'd270,32'd272,32'd274,32'd276,32'd278,32'd280,32'd282,32'd284,32'd286,32'd288,32'd290,32'd292,32'd294,32'd296,32'd298,32'd300,32'd302,32'd304,32'd306,32'd308,32'd310,32'd312,32'd314,32'd316,32'd318,32'd320,32'd322,32'd324,32'd326,32'd328,32'd330,32'd332,32'd334,32'd336,32'd338,32'd340,32'd342,32'd344,32'd346,32'd348,32'd350,32'd352,32'd354,32'd356,32'd358,32'd360,32'd362,32'd364,32'd366,32'd368,32'd370,32'd372,32'd374,32'd376,32'd378,32'd380,32'd382,32'd384,32'd386,32'd388,32'd390,32'd392,32'd394,32'd396,32'd398,32'd400,32'd402,32'd404,32'd406,32'd408,32'd410,32'd412,32'd414,32'd416,32'd418,32'd420,32'd422,32'd424,32'd426,32'd428,32'd430,32'd432,32'd434,32'd436,32'd438,32'd440,32'd442,32'd444,32'd446,32'd448,32'd450,32'd452,32'd454,32'd456,32'd458,32'd460,32'd462,32'd464,32'd466,32'd468,32'd470,32'd472,32'd474,32'd476,32'd478,32'd480,32'd482,32'd484,32'd486,32'd488,32'd490,32'd492,32'd494,32'd496,32'd498,32'd500,32'd502,32'd504,32'd506,32'd508,32'd510,32'd512,32'd514,32'd516,32'd518,32'd520,32'd522,32'd524,32'd526,32'd528,32'd530,32'd532,32'd534,32'd536,32'd538,32'd540,32'd542,32'd544,32'd546,32'd548,32'd550,32'd552,32'd554,32'd556,32'd558,32'd560,32'd562,32'd564,32'd566,32'd568,32'd570,32'd572,32'd574,32'd576,32'd578,32'd580,32'd582,32'd584,32'd586,32'd588,32'd590,32'd592,32'd594,32'd596,32'd598,32'd600,32'd602,32'd604,32'd606,32'd608,32'd610,32'd612,32'd614,32'd616,32'd618,32'd620,32'd622,32'd624,32'd626,32'd628,32'd630,32'd632,32'd634,32'd636,32'd638,32'd640,32'd642,32'd644,32'd646,32'd648,32'd650,32'd652,32'd654,32'd656,32'd658,32'd660,32'd662,32'd664,32'd666,32'd668,32'd670,32'd672,32'd674,32'd676,32'd678,32'd680,32'd682,32'd684,32'd686,32'd688,32'd690,32'd692,32'd694,32'd696,32'd698,32'd700,32'd702,32'd704,32'd706,32'd708,32'd710,32'd712,32'd714,32'd716,32'd718,32'd720,32'd722,32'd724,32'd726,32'd728,32'd730,32'd732,32'd734,32'd736,32'd738,32'd740,32'd742,32'd744,32'd746,32'd748,32'd750,32'd752,32'd754,32'd756,32'd758,32'd760,32'd762,32'd764,32'd766,32'd768,32'd770,32'd772,32'd774,32'd776,32'd778,32'd780,32'd782,32'd784,32'd786,32'd788,32'd790,32'd792,32'd794,32'd796,32'd798 };matrix[5]='{32'd0,32'd5,32'd10,32'd15,32'd20,32'd25,32'd30,32'd35,32'd40,32'd45,32'd50,32'd55,32'd60,32'd65,32'd70,32'd75,32'd80,32'd85,32'd90,32'd95,32'd100,32'd105,32'd110,32'd115,32'd120,32'd125,32'd130,32'd135,32'd140,32'd145,32'd150,32'd155,32'd160,32'd165,32'd170,32'd175,32'd180,32'd185,32'd190,32'd195,32'd200,32'd205,32'd210,32'd215,32'd220,32'd225,32'd230,32'd235,32'd240,32'd245,32'd250,32'd255,32'd260,32'd265,32'd270,32'd275,32'd280,32'd285,32'd290,32'd295,32'd300,32'd305,32'd310,32'd315,32'd320,32'd325,32'd330,32'd335,32'd340,32'd345,32'd350,32'd355,32'd360,32'd365,32'd370,32'd375,32'd380,32'd385,32'd390,32'd395,32'd400,32'd405,32'd410,32'd415,32'd420,32'd425,32'd430,32'd435,32'd440,32'd445,32'd450,32'd455,32'd460,32'd465,32'd470,32'd475,32'd480,32'd485,32'd490,32'd495,32'd500,32'd505,32'd510,32'd515,32'd520,32'd525,32'd530,32'd535,32'd540,32'd545,32'd550,32'd555,32'd560,32'd565,32'd570,32'd575,32'd580,32'd585,32'd590,32'd595,32'd600,32'd605,32'd610,32'd615,32'd620,32'd625,32'd630,32'd635,32'd640,32'd645,32'd650,32'd655,32'd660,32'd665,32'd670,32'd675,32'd680,32'd685,32'd690,32'd695,32'd700,32'd705,32'd710,32'd715,32'd720,32'd725,32'd730,32'd735,32'd740,32'd745,32'd750,32'd755,32'd760,32'd765,32'd770,32'd775,32'd780,32'd785,32'd790,32'd795,32'd800,32'd805,32'd810,32'd815,32'd820,32'd825,32'd830,32'd835,32'd840,32'd845,32'd850,32'd855,32'd860,32'd865,32'd870,32'd875,32'd880,32'd885,32'd890,32'd895,32'd900,32'd905,32'd910,32'd915,32'd920,32'd925,32'd930,32'd935,32'd940,32'd945,32'd950,32'd955,32'd960,32'd965,32'd970,32'd975,32'd980,32'd985,32'd990,32'd995,32'd1000,32'd1005,32'd1010,32'd1015,32'd1020,32'd1025,32'd1030,32'd1035,32'd1040,32'd1045,32'd1050,32'd1055,32'd1060,32'd1065,32'd1070,32'd1075,32'd1080,32'd1085,32'd1090,32'd1095,32'd1100,32'd1105,32'd1110,32'd1115,32'd1120,32'd1125,32'd1130,32'd1135,32'd1140,32'd1145,32'd1150,32'd1155,32'd1160,32'd1165,32'd1170,32'd1175,32'd1180,32'd1185,32'd1190,32'd1195,32'd1200,32'd1205,32'd1210,32'd1215,32'd1220,32'd1225,32'd1230,32'd1235,32'd1240,32'd1245,32'd1250,32'd1255,32'd1260,32'd1265,32'd1270,32'd1275,32'd1280,32'd1285,32'd1290,32'd1295,32'd1300,32'd1305,32'd1310,32'd1315,32'd1320,32'd1325,32'd1330,32'd1335,32'd1340,32'd1345,32'd1350,32'd1355,32'd1360,32'd1365,32'd1370,32'd1375,32'd1380,32'd1385,32'd1390,32'd1395,32'd1400,32'd1405,32'd1410,32'd1415,32'd1420,32'd1425,32'd1430,32'd1435,32'd1440,32'd1445,32'd1450,32'd1455,32'd1460,32'd1465,32'd1470,32'd1475,32'd1480,32'd1485,32'd1490,32'd1495,32'd1500,32'd1505,32'd1510,32'd1515,32'd1520,32'd1525,32'd1530,32'd1535,32'd1540,32'd1545,32'd1550,32'd1555,32'd1560,32'd1565,32'd1570,32'd1575,32'd1580,32'd1585,32'd1590,32'd1595,32'd1600,32'd1605,32'd1610,32'd1615,32'd1620,32'd1625,32'd1630,32'd1635,32'd1640,32'd1645,32'd1650,32'd1655,32'd1660,32'd1665,32'd1670,32'd1675,32'd1680,32'd1685,32'd1690,32'd1695,32'd1700,32'd1705,32'd1710,32'd1715,32'd1720,32'd1725,32'd1730,32'd1735,32'd1740,32'd1745,32'd1750,32'd1755,32'd1760,32'd1765,32'd1770,32'd1775,32'd1780,32'd1785,32'd1790,32'd1795,32'd1800,32'd1805,32'd1810,32'd1815,32'd1820,32'd1825,32'd1830,32'd1835,32'd1840,32'd1845,32'd1850,32'd1855,32'd1860,32'd1865,32'd1870,32'd1875,32'd1880,32'd1885,32'd1890,32'd1895,32'd1900,32'd1905,32'd1910,32'd1915,32'd1920,32'd1925,32'd1930,32'd1935,32'd1940,32'd1945,32'd1950,32'd1955,32'd1960,32'd1965,32'd1970,32'd1975,32'd1980,32'd1985,32'd1990,32'd1995 };matrix[4]='{32'd0,32'd4,32'd8,32'd12,32'd16,32'd20,32'd24,32'd28,32'd32,32'd36,32'd40,32'd44,32'd48,32'd52,32'd56,32'd60,32'd64,32'd68,32'd72,32'd76,32'd80,32'd84,32'd88,32'd92,32'd96,32'd100,32'd104,32'd108,32'd112,32'd116,32'd120,32'd124,32'd128,32'd132,32'd136,32'd140,32'd144,32'd148,32'd152,32'd156,32'd160,32'd164,32'd168,32'd172,32'd176,32'd180,32'd184,32'd188,32'd192,32'd196,32'd200,32'd204,32'd208,32'd212,32'd216,32'd220,32'd224,32'd228,32'd232,32'd236,32'd240,32'd244,32'd248,32'd252,32'd256,32'd260,32'd264,32'd268,32'd272,32'd276,32'd280,32'd284,32'd288,32'd292,32'd296,32'd300,32'd304,32'd308,32'd312,32'd316,32'd320,32'd324,32'd328,32'd332,32'd336,32'd340,32'd344,32'd348,32'd352,32'd356,32'd360,32'd364,32'd368,32'd372,32'd376,32'd380,32'd384,32'd388,32'd392,32'd396,32'd400,32'd404,32'd408,32'd412,32'd416,32'd420,32'd424,32'd428,32'd432,32'd436,32'd440,32'd444,32'd448,32'd452,32'd456,32'd460,32'd464,32'd468,32'd472,32'd476,32'd480,32'd484,32'd488,32'd492,32'd496,32'd500,32'd504,32'd508,32'd512,32'd516,32'd520,32'd524,32'd528,32'd532,32'd536,32'd540,32'd544,32'd548,32'd552,32'd556,32'd560,32'd564,32'd568,32'd572,32'd576,32'd580,32'd584,32'd588,32'd592,32'd596,32'd600,32'd604,32'd608,32'd612,32'd616,32'd620,32'd624,32'd628,32'd632,32'd636,32'd640,32'd644,32'd648,32'd652,32'd656,32'd660,32'd664,32'd668,32'd672,32'd676,32'd680,32'd684,32'd688,32'd692,32'd696,32'd700,32'd704,32'd708,32'd712,32'd716,32'd720,32'd724,32'd728,32'd732,32'd736,32'd740,32'd744,32'd748,32'd752,32'd756,32'd760,32'd764,32'd768,32'd772,32'd776,32'd780,32'd784,32'd788,32'd792,32'd796,32'd800,32'd804,32'd808,32'd812,32'd816,32'd820,32'd824,32'd828,32'd832,32'd836,32'd840,32'd844,32'd848,32'd852,32'd856,32'd860,32'd864,32'd868,32'd872,32'd876,32'd880,32'd884,32'd888,32'd892,32'd896,32'd900,32'd904,32'd908,32'd912,32'd916,32'd920,32'd924,32'd928,32'd932,32'd936,32'd940,32'd944,32'd948,32'd952,32'd956,32'd960,32'd964,32'd968,32'd972,32'd976,32'd980,32'd984,32'd988,32'd992,32'd996,32'd1000,32'd1004,32'd1008,32'd1012,32'd1016,32'd1020,32'd1024,32'd1028,32'd1032,32'd1036,32'd1040,32'd1044,32'd1048,32'd1052,32'd1056,32'd1060,32'd1064,32'd1068,32'd1072,32'd1076,32'd1080,32'd1084,32'd1088,32'd1092,32'd1096,32'd1100,32'd1104,32'd1108,32'd1112,32'd1116,32'd1120,32'd1124,32'd1128,32'd1132,32'd1136,32'd1140,32'd1144,32'd1148,32'd1152,32'd1156,32'd1160,32'd1164,32'd1168,32'd1172,32'd1176,32'd1180,32'd1184,32'd1188,32'd1192,32'd1196,32'd1200,32'd1204,32'd1208,32'd1212,32'd1216,32'd1220,32'd1224,32'd1228,32'd1232,32'd1236,32'd1240,32'd1244,32'd1248,32'd1252,32'd1256,32'd1260,32'd1264,32'd1268,32'd1272,32'd1276,32'd1280,32'd1284,32'd1288,32'd1292,32'd1296,32'd1300,32'd1304,32'd1308,32'd1312,32'd1316,32'd1320,32'd1324,32'd1328,32'd1332,32'd1336,32'd1340,32'd1344,32'd1348,32'd1352,32'd1356,32'd1360,32'd1364,32'd1368,32'd1372,32'd1376,32'd1380,32'd1384,32'd1388,32'd1392,32'd1396,32'd1400,32'd1404,32'd1408,32'd1412,32'd1416,32'd1420,32'd1424,32'd1428,32'd1432,32'd1436,32'd1440,32'd1444,32'd1448,32'd1452,32'd1456,32'd1460,32'd1464,32'd1468,32'd1472,32'd1476,32'd1480,32'd1484,32'd1488,32'd1492,32'd1496,32'd1500,32'd1504,32'd1508,32'd1512,32'd1516,32'd1520,32'd1524,32'd1528,32'd1532,32'd1536,32'd1540,32'd1544,32'd1548,32'd1552,32'd1556,32'd1560,32'd1564,32'd1568,32'd1572,32'd1576,32'd1580,32'd1584,32'd1588,32'd1592,32'd1596 };matrix[3]='{32'd0,32'd3,32'd6,32'd9,32'd12,32'd15,32'd18,32'd21,32'd24,32'd27,32'd30,32'd33,32'd36,32'd39,32'd42,32'd45,32'd48,32'd51,32'd54,32'd57,32'd60,32'd63,32'd66,32'd69,32'd72,32'd75,32'd78,32'd81,32'd84,32'd87,32'd90,32'd93,32'd96,32'd99,32'd102,32'd105,32'd108,32'd111,32'd114,32'd117,32'd120,32'd123,32'd126,32'd129,32'd132,32'd135,32'd138,32'd141,32'd144,32'd147,32'd150,32'd153,32'd156,32'd159,32'd162,32'd165,32'd168,32'd171,32'd174,32'd177,32'd180,32'd183,32'd186,32'd189,32'd192,32'd195,32'd198,32'd201,32'd204,32'd207,32'd210,32'd213,32'd216,32'd219,32'd222,32'd225,32'd228,32'd231,32'd234,32'd237,32'd240,32'd243,32'd246,32'd249,32'd252,32'd255,32'd258,32'd261,32'd264,32'd267,32'd270,32'd273,32'd276,32'd279,32'd282,32'd285,32'd288,32'd291,32'd294,32'd297,32'd300,32'd303,32'd306,32'd309,32'd312,32'd315,32'd318,32'd321,32'd324,32'd327,32'd330,32'd333,32'd336,32'd339,32'd342,32'd345,32'd348,32'd351,32'd354,32'd357,32'd360,32'd363,32'd366,32'd369,32'd372,32'd375,32'd378,32'd381,32'd384,32'd387,32'd390,32'd393,32'd396,32'd399,32'd402,32'd405,32'd408,32'd411,32'd414,32'd417,32'd420,32'd423,32'd426,32'd429,32'd432,32'd435,32'd438,32'd441,32'd444,32'd447,32'd450,32'd453,32'd456,32'd459,32'd462,32'd465,32'd468,32'd471,32'd474,32'd477,32'd480,32'd483,32'd486,32'd489,32'd492,32'd495,32'd498,32'd501,32'd504,32'd507,32'd510,32'd513,32'd516,32'd519,32'd522,32'd525,32'd528,32'd531,32'd534,32'd537,32'd540,32'd543,32'd546,32'd549,32'd552,32'd555,32'd558,32'd561,32'd564,32'd567,32'd570,32'd573,32'd576,32'd579,32'd582,32'd585,32'd588,32'd591,32'd594,32'd597,32'd600,32'd603,32'd606,32'd609,32'd612,32'd615,32'd618,32'd621,32'd624,32'd627,32'd630,32'd633,32'd636,32'd639,32'd642,32'd645,32'd648,32'd651,32'd654,32'd657,32'd660,32'd663,32'd666,32'd669,32'd672,32'd675,32'd678,32'd681,32'd684,32'd687,32'd690,32'd693,32'd696,32'd699,32'd702,32'd705,32'd708,32'd711,32'd714,32'd717,32'd720,32'd723,32'd726,32'd729,32'd732,32'd735,32'd738,32'd741,32'd744,32'd747,32'd750,32'd753,32'd756,32'd759,32'd762,32'd765,32'd768,32'd771,32'd774,32'd777,32'd780,32'd783,32'd786,32'd789,32'd792,32'd795,32'd798,32'd801,32'd804,32'd807,32'd810,32'd813,32'd816,32'd819,32'd822,32'd825,32'd828,32'd831,32'd834,32'd837,32'd840,32'd843,32'd846,32'd849,32'd852,32'd855,32'd858,32'd861,32'd864,32'd867,32'd870,32'd873,32'd876,32'd879,32'd882,32'd885,32'd888,32'd891,32'd894,32'd897,32'd900,32'd903,32'd906,32'd909,32'd912,32'd915,32'd918,32'd921,32'd924,32'd927,32'd930,32'd933,32'd936,32'd939,32'd942,32'd945,32'd948,32'd951,32'd954,32'd957,32'd960,32'd963,32'd966,32'd969,32'd972,32'd975,32'd978,32'd981,32'd984,32'd987,32'd990,32'd993,32'd996,32'd999,32'd1002,32'd1005,32'd1008,32'd1011,32'd1014,32'd1017,32'd1020,32'd1023,32'd1026,32'd1029,32'd1032,32'd1035,32'd1038,32'd1041,32'd1044,32'd1047,32'd1050,32'd1053,32'd1056,32'd1059,32'd1062,32'd1065,32'd1068,32'd1071,32'd1074,32'd1077,32'd1080,32'd1083,32'd1086,32'd1089,32'd1092,32'd1095,32'd1098,32'd1101,32'd1104,32'd1107,32'd1110,32'd1113,32'd1116,32'd1119,32'd1122,32'd1125,32'd1128,32'd1131,32'd1134,32'd1137,32'd1140,32'd1143,32'd1146,32'd1149,32'd1152,32'd1155,32'd1158,32'd1161,32'd1164,32'd1167,32'd1170,32'd1173,32'd1176,32'd1179,32'd1182,32'd1185,32'd1188,32'd1191,32'd1194,32'd1197 };matrix[6]='{32'd0,32'd6,32'd12,32'd18,32'd24,32'd30,32'd36,32'd42,32'd48,32'd54,32'd60,32'd66,32'd72,32'd78,32'd84,32'd90,32'd96,32'd102,32'd108,32'd114,32'd120,32'd126,32'd132,32'd138,32'd144,32'd150,32'd156,32'd162,32'd168,32'd174,32'd180,32'd186,32'd192,32'd198,32'd204,32'd210,32'd216,32'd222,32'd228,32'd234,32'd240,32'd246,32'd252,32'd258,32'd264,32'd270,32'd276,32'd282,32'd288,32'd294,32'd300,32'd306,32'd312,32'd318,32'd324,32'd330,32'd336,32'd342,32'd348,32'd354,32'd360,32'd366,32'd372,32'd378,32'd384,32'd390,32'd396,32'd402,32'd408,32'd414,32'd420,32'd426,32'd432,32'd438,32'd444,32'd450,32'd456,32'd462,32'd468,32'd474,32'd480,32'd486,32'd492,32'd498,32'd504,32'd510,32'd516,32'd522,32'd528,32'd534,32'd540,32'd546,32'd552,32'd558,32'd564,32'd570,32'd576,32'd582,32'd588,32'd594,32'd600,32'd606,32'd612,32'd618,32'd624,32'd630,32'd636,32'd642,32'd648,32'd654,32'd660,32'd666,32'd672,32'd678,32'd684,32'd690,32'd696,32'd702,32'd708,32'd714,32'd720,32'd726,32'd732,32'd738,32'd744,32'd750,32'd756,32'd762,32'd768,32'd774,32'd780,32'd786,32'd792,32'd798,32'd804,32'd810,32'd816,32'd822,32'd828,32'd834,32'd840,32'd846,32'd852,32'd858,32'd864,32'd870,32'd876,32'd882,32'd888,32'd894,32'd900,32'd906,32'd912,32'd918,32'd924,32'd930,32'd936,32'd942,32'd948,32'd954,32'd960,32'd966,32'd972,32'd978,32'd984,32'd990,32'd996,32'd1002,32'd1008,32'd1014,32'd1020,32'd1026,32'd1032,32'd1038,32'd1044,32'd1050,32'd1056,32'd1062,32'd1068,32'd1074,32'd1080,32'd1086,32'd1092,32'd1098,32'd1104,32'd1110,32'd1116,32'd1122,32'd1128,32'd1134,32'd1140,32'd1146,32'd1152,32'd1158,32'd1164,32'd1170,32'd1176,32'd1182,32'd1188,32'd1194,32'd1200,32'd1206,32'd1212,32'd1218,32'd1224,32'd1230,32'd1236,32'd1242,32'd1248,32'd1254,32'd1260,32'd1266,32'd1272,32'd1278,32'd1284,32'd1290,32'd1296,32'd1302,32'd1308,32'd1314,32'd1320,32'd1326,32'd1332,32'd1338,32'd1344,32'd1350,32'd1356,32'd1362,32'd1368,32'd1374,32'd1380,32'd1386,32'd1392,32'd1398,32'd1404,32'd1410,32'd1416,32'd1422,32'd1428,32'd1434,32'd1440,32'd1446,32'd1452,32'd1458,32'd1464,32'd1470,32'd1476,32'd1482,32'd1488,32'd1494,32'd1500,32'd1506,32'd1512,32'd1518,32'd1524,32'd1530,32'd1536,32'd1542,32'd1548,32'd1554,32'd1560,32'd1566,32'd1572,32'd1578,32'd1584,32'd1590,32'd1596,32'd1602,32'd1608,32'd1614,32'd1620,32'd1626,32'd1632,32'd1638,32'd1644,32'd1650,32'd1656,32'd1662,32'd1668,32'd1674,32'd1680,32'd1686,32'd1692,32'd1698,32'd1704,32'd1710,32'd1716,32'd1722,32'd1728,32'd1734,32'd1740,32'd1746,32'd1752,32'd1758,32'd1764,32'd1770,32'd1776,32'd1782,32'd1788,32'd1794,32'd1800,32'd1806,32'd1812,32'd1818,32'd1824,32'd1830,32'd1836,32'd1842,32'd1848,32'd1854,32'd1860,32'd1866,32'd1872,32'd1878,32'd1884,32'd1890,32'd1896,32'd1902,32'd1908,32'd1914,32'd1920,32'd1926,32'd1932,32'd1938,32'd1944,32'd1950,32'd1956,32'd1962,32'd1968,32'd1974,32'd1980,32'd1986,32'd1992,32'd1998,32'd2004,32'd2010,32'd2016,32'd2022,32'd2028,32'd2034,32'd2040,32'd2046,32'd2052,32'd2058,32'd2064,32'd2070,32'd2076,32'd2082,32'd2088,32'd2094,32'd2100,32'd2106,32'd2112,32'd2118,32'd2124,32'd2130,32'd2136,32'd2142,32'd2148,32'd2154,32'd2160,32'd2166,32'd2172,32'd2178,32'd2184,32'd2190,32'd2196,32'd2202,32'd2208,32'd2214,32'd2220,32'd2226,32'd2232,32'd2238,32'd2244,32'd2250,32'd2256,32'd2262,32'd2268,32'd2274,32'd2280,32'd2286,32'd2292,32'd2298,32'd2304,32'd2310,32'd2316,32'd2322,32'd2328,32'd2334,32'd2340,32'd2346,32'd2352,32'd2358,32'd2364,32'd2370,32'd2376,32'd2382,32'd2388,32'd2394 };matrix[7]='{32'd0,32'd7,32'd14,32'd21,32'd28,32'd35,32'd42,32'd49,32'd56,32'd63,32'd70,32'd77,32'd84,32'd91,32'd98,32'd105,32'd112,32'd119,32'd126,32'd133,32'd140,32'd147,32'd154,32'd161,32'd168,32'd175,32'd182,32'd189,32'd196,32'd203,32'd210,32'd217,32'd224,32'd231,32'd238,32'd245,32'd252,32'd259,32'd266,32'd273,32'd280,32'd287,32'd294,32'd301,32'd308,32'd315,32'd322,32'd329,32'd336,32'd343,32'd350,32'd357,32'd364,32'd371,32'd378,32'd385,32'd392,32'd399,32'd406,32'd413,32'd420,32'd427,32'd434,32'd441,32'd448,32'd455,32'd462,32'd469,32'd476,32'd483,32'd490,32'd497,32'd504,32'd511,32'd518,32'd525,32'd532,32'd539,32'd546,32'd553,32'd560,32'd567,32'd574,32'd581,32'd588,32'd595,32'd602,32'd609,32'd616,32'd623,32'd630,32'd637,32'd644,32'd651,32'd658,32'd665,32'd672,32'd679,32'd686,32'd693,32'd700,32'd707,32'd714,32'd721,32'd728,32'd735,32'd742,32'd749,32'd756,32'd763,32'd770,32'd777,32'd784,32'd791,32'd798,32'd805,32'd812,32'd819,32'd826,32'd833,32'd840,32'd847,32'd854,32'd861,32'd868,32'd875,32'd882,32'd889,32'd896,32'd903,32'd910,32'd917,32'd924,32'd931,32'd938,32'd945,32'd952,32'd959,32'd966,32'd973,32'd980,32'd987,32'd994,32'd1001,32'd1008,32'd1015,32'd1022,32'd1029,32'd1036,32'd1043,32'd1050,32'd1057,32'd1064,32'd1071,32'd1078,32'd1085,32'd1092,32'd1099,32'd1106,32'd1113,32'd1120,32'd1127,32'd1134,32'd1141,32'd1148,32'd1155,32'd1162,32'd1169,32'd1176,32'd1183,32'd1190,32'd1197,32'd1204,32'd1211,32'd1218,32'd1225,32'd1232,32'd1239,32'd1246,32'd1253,32'd1260,32'd1267,32'd1274,32'd1281,32'd1288,32'd1295,32'd1302,32'd1309,32'd1316,32'd1323,32'd1330,32'd1337,32'd1344,32'd1351,32'd1358,32'd1365,32'd1372,32'd1379,32'd1386,32'd1393,32'd1400,32'd1407,32'd1414,32'd1421,32'd1428,32'd1435,32'd1442,32'd1449,32'd1456,32'd1463,32'd1470,32'd1477,32'd1484,32'd1491,32'd1498,32'd1505,32'd1512,32'd1519,32'd1526,32'd1533,32'd1540,32'd1547,32'd1554,32'd1561,32'd1568,32'd1575,32'd1582,32'd1589,32'd1596,32'd1603,32'd1610,32'd1617,32'd1624,32'd1631,32'd1638,32'd1645,32'd1652,32'd1659,32'd1666,32'd1673,32'd1680,32'd1687,32'd1694,32'd1701,32'd1708,32'd1715,32'd1722,32'd1729,32'd1736,32'd1743,32'd1750,32'd1757,32'd1764,32'd1771,32'd1778,32'd1785,32'd1792,32'd1799,32'd1806,32'd1813,32'd1820,32'd1827,32'd1834,32'd1841,32'd1848,32'd1855,32'd1862,32'd1869,32'd1876,32'd1883,32'd1890,32'd1897,32'd1904,32'd1911,32'd1918,32'd1925,32'd1932,32'd1939,32'd1946,32'd1953,32'd1960,32'd1967,32'd1974,32'd1981,32'd1988,32'd1995,32'd2002,32'd2009,32'd2016,32'd2023,32'd2030,32'd2037,32'd2044,32'd2051,32'd2058,32'd2065,32'd2072,32'd2079,32'd2086,32'd2093,32'd2100,32'd2107,32'd2114,32'd2121,32'd2128,32'd2135,32'd2142,32'd2149,32'd2156,32'd2163,32'd2170,32'd2177,32'd2184,32'd2191,32'd2198,32'd2205,32'd2212,32'd2219,32'd2226,32'd2233,32'd2240,32'd2247,32'd2254,32'd2261,32'd2268,32'd2275,32'd2282,32'd2289,32'd2296,32'd2303,32'd2310,32'd2317,32'd2324,32'd2331,32'd2338,32'd2345,32'd2352,32'd2359,32'd2366,32'd2373,32'd2380,32'd2387,32'd2394,32'd2401,32'd2408,32'd2415,32'd2422,32'd2429,32'd2436,32'd2443,32'd2450,32'd2457,32'd2464,32'd2471,32'd2478,32'd2485,32'd2492,32'd2499,32'd2506,32'd2513,32'd2520,32'd2527,32'd2534,32'd2541,32'd2548,32'd2555,32'd2562,32'd2569,32'd2576,32'd2583,32'd2590,32'd2597,32'd2604,32'd2611,32'd2618,32'd2625,32'd2632,32'd2639,32'd2646,32'd2653,32'd2660,32'd2667,32'd2674,32'd2681,32'd2688,32'd2695,32'd2702,32'd2709,32'd2716,32'd2723,32'd2730,32'd2737,32'd2744,32'd2751,32'd2758,32'd2765,32'd2772,32'd2779,32'd2786,32'd2793 };matrix[8]='{32'd0,32'd8,32'd16,32'd24,32'd32,32'd40,32'd48,32'd56,32'd64,32'd72,32'd80,32'd88,32'd96,32'd104,32'd112,32'd120,32'd128,32'd136,32'd144,32'd152,32'd160,32'd168,32'd176,32'd184,32'd192,32'd200,32'd208,32'd216,32'd224,32'd232,32'd240,32'd248,32'd256,32'd264,32'd272,32'd280,32'd288,32'd296,32'd304,32'd312,32'd320,32'd328,32'd336,32'd344,32'd352,32'd360,32'd368,32'd376,32'd384,32'd392,32'd400,32'd408,32'd416,32'd424,32'd432,32'd440,32'd448,32'd456,32'd464,32'd472,32'd480,32'd488,32'd496,32'd504,32'd512,32'd520,32'd528,32'd536,32'd544,32'd552,32'd560,32'd568,32'd576,32'd584,32'd592,32'd600,32'd608,32'd616,32'd624,32'd632,32'd640,32'd648,32'd656,32'd664,32'd672,32'd680,32'd688,32'd696,32'd704,32'd712,32'd720,32'd728,32'd736,32'd744,32'd752,32'd760,32'd768,32'd776,32'd784,32'd792,32'd800,32'd808,32'd816,32'd824,32'd832,32'd840,32'd848,32'd856,32'd864,32'd872,32'd880,32'd888,32'd896,32'd904,32'd912,32'd920,32'd928,32'd936,32'd944,32'd952,32'd960,32'd968,32'd976,32'd984,32'd992,32'd1000,32'd1008,32'd1016,32'd1024,32'd1032,32'd1040,32'd1048,32'd1056,32'd1064,32'd1072,32'd1080,32'd1088,32'd1096,32'd1104,32'd1112,32'd1120,32'd1128,32'd1136,32'd1144,32'd1152,32'd1160,32'd1168,32'd1176,32'd1184,32'd1192,32'd1200,32'd1208,32'd1216,32'd1224,32'd1232,32'd1240,32'd1248,32'd1256,32'd1264,32'd1272,32'd1280,32'd1288,32'd1296,32'd1304,32'd1312,32'd1320,32'd1328,32'd1336,32'd1344,32'd1352,32'd1360,32'd1368,32'd1376,32'd1384,32'd1392,32'd1400,32'd1408,32'd1416,32'd1424,32'd1432,32'd1440,32'd1448,32'd1456,32'd1464,32'd1472,32'd1480,32'd1488,32'd1496,32'd1504,32'd1512,32'd1520,32'd1528,32'd1536,32'd1544,32'd1552,32'd1560,32'd1568,32'd1576,32'd1584,32'd1592,32'd1600,32'd1608,32'd1616,32'd1624,32'd1632,32'd1640,32'd1648,32'd1656,32'd1664,32'd1672,32'd1680,32'd1688,32'd1696,32'd1704,32'd1712,32'd1720,32'd1728,32'd1736,32'd1744,32'd1752,32'd1760,32'd1768,32'd1776,32'd1784,32'd1792,32'd1800,32'd1808,32'd1816,32'd1824,32'd1832,32'd1840,32'd1848,32'd1856,32'd1864,32'd1872,32'd1880,32'd1888,32'd1896,32'd1904,32'd1912,32'd1920,32'd1928,32'd1936,32'd1944,32'd1952,32'd1960,32'd1968,32'd1976,32'd1984,32'd1992,32'd2000,32'd2008,32'd2016,32'd2024,32'd2032,32'd2040,32'd2048,32'd2056,32'd2064,32'd2072,32'd2080,32'd2088,32'd2096,32'd2104,32'd2112,32'd2120,32'd2128,32'd2136,32'd2144,32'd2152,32'd2160,32'd2168,32'd2176,32'd2184,32'd2192,32'd2200,32'd2208,32'd2216,32'd2224,32'd2232,32'd2240,32'd2248,32'd2256,32'd2264,32'd2272,32'd2280,32'd2288,32'd2296,32'd2304,32'd2312,32'd2320,32'd2328,32'd2336,32'd2344,32'd2352,32'd2360,32'd2368,32'd2376,32'd2384,32'd2392,32'd2400,32'd2408,32'd2416,32'd2424,32'd2432,32'd2440,32'd2448,32'd2456,32'd2464,32'd2472,32'd2480,32'd2488,32'd2496,32'd2504,32'd2512,32'd2520,32'd2528,32'd2536,32'd2544,32'd2552,32'd2560,32'd2568,32'd2576,32'd2584,32'd2592,32'd2600,32'd2608,32'd2616,32'd2624,32'd2632,32'd2640,32'd2648,32'd2656,32'd2664,32'd2672,32'd2680,32'd2688,32'd2696,32'd2704,32'd2712,32'd2720,32'd2728,32'd2736,32'd2744,32'd2752,32'd2760,32'd2768,32'd2776,32'd2784,32'd2792,32'd2800,32'd2808,32'd2816,32'd2824,32'd2832,32'd2840,32'd2848,32'd2856,32'd2864,32'd2872,32'd2880,32'd2888,32'd2896,32'd2904,32'd2912,32'd2920,32'd2928,32'd2936,32'd2944,32'd2952,32'd2960,32'd2968,32'd2976,32'd2984,32'd2992,32'd3000,32'd3008,32'd3016,32'd3024,32'd3032,32'd3040,32'd3048,32'd3056,32'd3064,32'd3072,32'd3080,32'd3088,32'd3096,32'd3104,32'd3112,32'd3120,32'd3128,32'd3136,32'd3144,32'd3152,32'd3160,32'd3168,32'd3176,32'd3184,32'd3192 };matrix[9]='{32'd0,32'd9,32'd18,32'd27,32'd36,32'd45,32'd54,32'd63,32'd72,32'd81,32'd90,32'd99,32'd108,32'd117,32'd126,32'd135,32'd144,32'd153,32'd162,32'd171,32'd180,32'd189,32'd198,32'd207,32'd216,32'd225,32'd234,32'd243,32'd252,32'd261,32'd270,32'd279,32'd288,32'd297,32'd306,32'd315,32'd324,32'd333,32'd342,32'd351,32'd360,32'd369,32'd378,32'd387,32'd396,32'd405,32'd414,32'd423,32'd432,32'd441,32'd450,32'd459,32'd468,32'd477,32'd486,32'd495,32'd504,32'd513,32'd522,32'd531,32'd540,32'd549,32'd558,32'd567,32'd576,32'd585,32'd594,32'd603,32'd612,32'd621,32'd630,32'd639,32'd648,32'd657,32'd666,32'd675,32'd684,32'd693,32'd702,32'd711,32'd720,32'd729,32'd738,32'd747,32'd756,32'd765,32'd774,32'd783,32'd792,32'd801,32'd810,32'd819,32'd828,32'd837,32'd846,32'd855,32'd864,32'd873,32'd882,32'd891,32'd900,32'd909,32'd918,32'd927,32'd936,32'd945,32'd954,32'd963,32'd972,32'd981,32'd990,32'd999,32'd1008,32'd1017,32'd1026,32'd1035,32'd1044,32'd1053,32'd1062,32'd1071,32'd1080,32'd1089,32'd1098,32'd1107,32'd1116,32'd1125,32'd1134,32'd1143,32'd1152,32'd1161,32'd1170,32'd1179,32'd1188,32'd1197,32'd1206,32'd1215,32'd1224,32'd1233,32'd1242,32'd1251,32'd1260,32'd1269,32'd1278,32'd1287,32'd1296,32'd1305,32'd1314,32'd1323,32'd1332,32'd1341,32'd1350,32'd1359,32'd1368,32'd1377,32'd1386,32'd1395,32'd1404,32'd1413,32'd1422,32'd1431,32'd1440,32'd1449,32'd1458,32'd1467,32'd1476,32'd1485,32'd1494,32'd1503,32'd1512,32'd1521,32'd1530,32'd1539,32'd1548,32'd1557,32'd1566,32'd1575,32'd1584,32'd1593,32'd1602,32'd1611,32'd1620,32'd1629,32'd1638,32'd1647,32'd1656,32'd1665,32'd1674,32'd1683,32'd1692,32'd1701,32'd1710,32'd1719,32'd1728,32'd1737,32'd1746,32'd1755,32'd1764,32'd1773,32'd1782,32'd1791,32'd1800,32'd1809,32'd1818,32'd1827,32'd1836,32'd1845,32'd1854,32'd1863,32'd1872,32'd1881,32'd1890,32'd1899,32'd1908,32'd1917,32'd1926,32'd1935,32'd1944,32'd1953,32'd1962,32'd1971,32'd1980,32'd1989,32'd1998,32'd2007,32'd2016,32'd2025,32'd2034,32'd2043,32'd2052,32'd2061,32'd2070,32'd2079,32'd2088,32'd2097,32'd2106,32'd2115,32'd2124,32'd2133,32'd2142,32'd2151,32'd2160,32'd2169,32'd2178,32'd2187,32'd2196,32'd2205,32'd2214,32'd2223,32'd2232,32'd2241,32'd2250,32'd2259,32'd2268,32'd2277,32'd2286,32'd2295,32'd2304,32'd2313,32'd2322,32'd2331,32'd2340,32'd2349,32'd2358,32'd2367,32'd2376,32'd2385,32'd2394,32'd2403,32'd2412,32'd2421,32'd2430,32'd2439,32'd2448,32'd2457,32'd2466,32'd2475,32'd2484,32'd2493,32'd2502,32'd2511,32'd2520,32'd2529,32'd2538,32'd2547,32'd2556,32'd2565,32'd2574,32'd2583,32'd2592,32'd2601,32'd2610,32'd2619,32'd2628,32'd2637,32'd2646,32'd2655,32'd2664,32'd2673,32'd2682,32'd2691,32'd2700,32'd2709,32'd2718,32'd2727,32'd2736,32'd2745,32'd2754,32'd2763,32'd2772,32'd2781,32'd2790,32'd2799,32'd2808,32'd2817,32'd2826,32'd2835,32'd2844,32'd2853,32'd2862,32'd2871,32'd2880,32'd2889,32'd2898,32'd2907,32'd2916,32'd2925,32'd2934,32'd2943,32'd2952,32'd2961,32'd2970,32'd2979,32'd2988,32'd2997,32'd3006,32'd3015,32'd3024,32'd3033,32'd3042,32'd3051,32'd3060,32'd3069,32'd3078,32'd3087,32'd3096,32'd3105,32'd3114,32'd3123,32'd3132,32'd3141,32'd3150,32'd3159,32'd3168,32'd3177,32'd3186,32'd3195,32'd3204,32'd3213,32'd3222,32'd3231,32'd3240,32'd3249,32'd3258,32'd3267,32'd3276,32'd3285,32'd3294,32'd3303,32'd3312,32'd3321,32'd3330,32'd3339,32'd3348,32'd3357,32'd3366,32'd3375,32'd3384,32'd3393,32'd3402,32'd3411,32'd3420,32'd3429,32'd3438,32'd3447,32'd3456,32'd3465,32'd3474,32'd3483,32'd3492,32'd3501,32'd3510,32'd3519,32'd3528,32'd3537,32'd3546,32'd3555,32'd3564,32'd3573,32'd3582,32'd3591 };matrix[11]='{32'd0,32'd11,32'd22,32'd33,32'd44,32'd55,32'd66,32'd77,32'd88,32'd99,32'd110,32'd121,32'd132,32'd143,32'd154,32'd165,32'd176,32'd187,32'd198,32'd209,32'd220,32'd231,32'd242,32'd253,32'd264,32'd275,32'd286,32'd297,32'd308,32'd319,32'd330,32'd341,32'd352,32'd363,32'd374,32'd385,32'd396,32'd407,32'd418,32'd429,32'd440,32'd451,32'd462,32'd473,32'd484,32'd495,32'd506,32'd517,32'd528,32'd539,32'd550,32'd561,32'd572,32'd583,32'd594,32'd605,32'd616,32'd627,32'd638,32'd649,32'd660,32'd671,32'd682,32'd693,32'd704,32'd715,32'd726,32'd737,32'd748,32'd759,32'd770,32'd781,32'd792,32'd803,32'd814,32'd825,32'd836,32'd847,32'd858,32'd869,32'd880,32'd891,32'd902,32'd913,32'd924,32'd935,32'd946,32'd957,32'd968,32'd979,32'd990,32'd1001,32'd1012,32'd1023,32'd1034,32'd1045,32'd1056,32'd1067,32'd1078,32'd1089,32'd1100,32'd1111,32'd1122,32'd1133,32'd1144,32'd1155,32'd1166,32'd1177,32'd1188,32'd1199,32'd1210,32'd1221,32'd1232,32'd1243,32'd1254,32'd1265,32'd1276,32'd1287,32'd1298,32'd1309,32'd1320,32'd1331,32'd1342,32'd1353,32'd1364,32'd1375,32'd1386,32'd1397,32'd1408,32'd1419,32'd1430,32'd1441,32'd1452,32'd1463,32'd1474,32'd1485,32'd1496,32'd1507,32'd1518,32'd1529,32'd1540,32'd1551,32'd1562,32'd1573,32'd1584,32'd1595,32'd1606,32'd1617,32'd1628,32'd1639,32'd1650,32'd1661,32'd1672,32'd1683,32'd1694,32'd1705,32'd1716,32'd1727,32'd1738,32'd1749,32'd1760,32'd1771,32'd1782,32'd1793,32'd1804,32'd1815,32'd1826,32'd1837,32'd1848,32'd1859,32'd1870,32'd1881,32'd1892,32'd1903,32'd1914,32'd1925,32'd1936,32'd1947,32'd1958,32'd1969,32'd1980,32'd1991,32'd2002,32'd2013,32'd2024,32'd2035,32'd2046,32'd2057,32'd2068,32'd2079,32'd2090,32'd2101,32'd2112,32'd2123,32'd2134,32'd2145,32'd2156,32'd2167,32'd2178,32'd2189,32'd2200,32'd2211,32'd2222,32'd2233,32'd2244,32'd2255,32'd2266,32'd2277,32'd2288,32'd2299,32'd2310,32'd2321,32'd2332,32'd2343,32'd2354,32'd2365,32'd2376,32'd2387,32'd2398,32'd2409,32'd2420,32'd2431,32'd2442,32'd2453,32'd2464,32'd2475,32'd2486,32'd2497,32'd2508,32'd2519,32'd2530,32'd2541,32'd2552,32'd2563,32'd2574,32'd2585,32'd2596,32'd2607,32'd2618,32'd2629,32'd2640,32'd2651,32'd2662,32'd2673,32'd2684,32'd2695,32'd2706,32'd2717,32'd2728,32'd2739,32'd2750,32'd2761,32'd2772,32'd2783,32'd2794,32'd2805,32'd2816,32'd2827,32'd2838,32'd2849,32'd2860,32'd2871,32'd2882,32'd2893,32'd2904,32'd2915,32'd2926,32'd2937,32'd2948,32'd2959,32'd2970,32'd2981,32'd2992,32'd3003,32'd3014,32'd3025,32'd3036,32'd3047,32'd3058,32'd3069,32'd3080,32'd3091,32'd3102,32'd3113,32'd3124,32'd3135,32'd3146,32'd3157,32'd3168,32'd3179,32'd3190,32'd3201,32'd3212,32'd3223,32'd3234,32'd3245,32'd3256,32'd3267,32'd3278,32'd3289,32'd3300,32'd3311,32'd3322,32'd3333,32'd3344,32'd3355,32'd3366,32'd3377,32'd3388,32'd3399,32'd3410,32'd3421,32'd3432,32'd3443,32'd3454,32'd3465,32'd3476,32'd3487,32'd3498,32'd3509,32'd3520,32'd3531,32'd3542,32'd3553,32'd3564,32'd3575,32'd3586,32'd3597,32'd3608,32'd3619,32'd3630,32'd3641,32'd3652,32'd3663,32'd3674,32'd3685,32'd3696,32'd3707,32'd3718,32'd3729,32'd3740,32'd3751,32'd3762,32'd3773,32'd3784,32'd3795,32'd3806,32'd3817,32'd3828,32'd3839,32'd3850,32'd3861,32'd3872,32'd3883,32'd3894,32'd3905,32'd3916,32'd3927,32'd3938,32'd3949,32'd3960,32'd3971,32'd3982,32'd3993,32'd4004,32'd4015,32'd4026,32'd4037,32'd4048,32'd4059,32'd4070,32'd4081,32'd4092,32'd4103,32'd4114,32'd4125,32'd4136,32'd4147,32'd4158,32'd4169,32'd4180,32'd4191,32'd4202,32'd4213,32'd4224,32'd4235,32'd4246,32'd4257,32'd4268,32'd4279,32'd4290,32'd4301,32'd4312,32'd4323,32'd4334,32'd4345,32'd4356,32'd4367,32'd4378,32'd4389 };matrix[10]='{32'd0,32'd10,32'd20,32'd30,32'd40,32'd50,32'd60,32'd70,32'd80,32'd90,32'd100,32'd110,32'd120,32'd130,32'd140,32'd150,32'd160,32'd170,32'd180,32'd190,32'd200,32'd210,32'd220,32'd230,32'd240,32'd250,32'd260,32'd270,32'd280,32'd290,32'd300,32'd310,32'd320,32'd330,32'd340,32'd350,32'd360,32'd370,32'd380,32'd390,32'd400,32'd410,32'd420,32'd430,32'd440,32'd450,32'd460,32'd470,32'd480,32'd490,32'd500,32'd510,32'd520,32'd530,32'd540,32'd550,32'd560,32'd570,32'd580,32'd590,32'd600,32'd610,32'd620,32'd630,32'd640,32'd650,32'd660,32'd670,32'd680,32'd690,32'd700,32'd710,32'd720,32'd730,32'd740,32'd750,32'd760,32'd770,32'd780,32'd790,32'd800,32'd810,32'd820,32'd830,32'd840,32'd850,32'd860,32'd870,32'd880,32'd890,32'd900,32'd910,32'd920,32'd930,32'd940,32'd950,32'd960,32'd970,32'd980,32'd990,32'd1000,32'd1010,32'd1020,32'd1030,32'd1040,32'd1050,32'd1060,32'd1070,32'd1080,32'd1090,32'd1100,32'd1110,32'd1120,32'd1130,32'd1140,32'd1150,32'd1160,32'd1170,32'd1180,32'd1190,32'd1200,32'd1210,32'd1220,32'd1230,32'd1240,32'd1250,32'd1260,32'd1270,32'd1280,32'd1290,32'd1300,32'd1310,32'd1320,32'd1330,32'd1340,32'd1350,32'd1360,32'd1370,32'd1380,32'd1390,32'd1400,32'd1410,32'd1420,32'd1430,32'd1440,32'd1450,32'd1460,32'd1470,32'd1480,32'd1490,32'd1500,32'd1510,32'd1520,32'd1530,32'd1540,32'd1550,32'd1560,32'd1570,32'd1580,32'd1590,32'd1600,32'd1610,32'd1620,32'd1630,32'd1640,32'd1650,32'd1660,32'd1670,32'd1680,32'd1690,32'd1700,32'd1710,32'd1720,32'd1730,32'd1740,32'd1750,32'd1760,32'd1770,32'd1780,32'd1790,32'd1800,32'd1810,32'd1820,32'd1830,32'd1840,32'd1850,32'd1860,32'd1870,32'd1880,32'd1890,32'd1900,32'd1910,32'd1920,32'd1930,32'd1940,32'd1950,32'd1960,32'd1970,32'd1980,32'd1990,32'd2000,32'd2010,32'd2020,32'd2030,32'd2040,32'd2050,32'd2060,32'd2070,32'd2080,32'd2090,32'd2100,32'd2110,32'd2120,32'd2130,32'd2140,32'd2150,32'd2160,32'd2170,32'd2180,32'd2190,32'd2200,32'd2210,32'd2220,32'd2230,32'd2240,32'd2250,32'd2260,32'd2270,32'd2280,32'd2290,32'd2300,32'd2310,32'd2320,32'd2330,32'd2340,32'd2350,32'd2360,32'd2370,32'd2380,32'd2390,32'd2400,32'd2410,32'd2420,32'd2430,32'd2440,32'd2450,32'd2460,32'd2470,32'd2480,32'd2490,32'd2500,32'd2510,32'd2520,32'd2530,32'd2540,32'd2550,32'd2560,32'd2570,32'd2580,32'd2590,32'd2600,32'd2610,32'd2620,32'd2630,32'd2640,32'd2650,32'd2660,32'd2670,32'd2680,32'd2690,32'd2700,32'd2710,32'd2720,32'd2730,32'd2740,32'd2750,32'd2760,32'd2770,32'd2780,32'd2790,32'd2800,32'd2810,32'd2820,32'd2830,32'd2840,32'd2850,32'd2860,32'd2870,32'd2880,32'd2890,32'd2900,32'd2910,32'd2920,32'd2930,32'd2940,32'd2950,32'd2960,32'd2970,32'd2980,32'd2990,32'd3000,32'd3010,32'd3020,32'd3030,32'd3040,32'd3050,32'd3060,32'd3070,32'd3080,32'd3090,32'd3100,32'd3110,32'd3120,32'd3130,32'd3140,32'd3150,32'd3160,32'd3170,32'd3180,32'd3190,32'd3200,32'd3210,32'd3220,32'd3230,32'd3240,32'd3250,32'd3260,32'd3270,32'd3280,32'd3290,32'd3300,32'd3310,32'd3320,32'd3330,32'd3340,32'd3350,32'd3360,32'd3370,32'd3380,32'd3390,32'd3400,32'd3410,32'd3420,32'd3430,32'd3440,32'd3450,32'd3460,32'd3470,32'd3480,32'd3490,32'd3500,32'd3510,32'd3520,32'd3530,32'd3540,32'd3550,32'd3560,32'd3570,32'd3580,32'd3590,32'd3600,32'd3610,32'd3620,32'd3630,32'd3640,32'd3650,32'd3660,32'd3670,32'd3680,32'd3690,32'd3700,32'd3710,32'd3720,32'd3730,32'd3740,32'd3750,32'd3760,32'd3770,32'd3780,32'd3790,32'd3800,32'd3810,32'd3820,32'd3830,32'd3840,32'd3850,32'd3860,32'd3870,32'd3880,32'd3890,32'd3900,32'd3910,32'd3920,32'd3930,32'd3940,32'd3950,32'd3960,32'd3970,32'd3980,32'd3990 };matrix[12]='{32'd0,32'd12,32'd24,32'd36,32'd48,32'd60,32'd72,32'd84,32'd96,32'd108,32'd120,32'd132,32'd144,32'd156,32'd168,32'd180,32'd192,32'd204,32'd216,32'd228,32'd240,32'd252,32'd264,32'd276,32'd288,32'd300,32'd312,32'd324,32'd336,32'd348,32'd360,32'd372,32'd384,32'd396,32'd408,32'd420,32'd432,32'd444,32'd456,32'd468,32'd480,32'd492,32'd504,32'd516,32'd528,32'd540,32'd552,32'd564,32'd576,32'd588,32'd600,32'd612,32'd624,32'd636,32'd648,32'd660,32'd672,32'd684,32'd696,32'd708,32'd720,32'd732,32'd744,32'd756,32'd768,32'd780,32'd792,32'd804,32'd816,32'd828,32'd840,32'd852,32'd864,32'd876,32'd888,32'd900,32'd912,32'd924,32'd936,32'd948,32'd960,32'd972,32'd984,32'd996,32'd1008,32'd1020,32'd1032,32'd1044,32'd1056,32'd1068,32'd1080,32'd1092,32'd1104,32'd1116,32'd1128,32'd1140,32'd1152,32'd1164,32'd1176,32'd1188,32'd1200,32'd1212,32'd1224,32'd1236,32'd1248,32'd1260,32'd1272,32'd1284,32'd1296,32'd1308,32'd1320,32'd1332,32'd1344,32'd1356,32'd1368,32'd1380,32'd1392,32'd1404,32'd1416,32'd1428,32'd1440,32'd1452,32'd1464,32'd1476,32'd1488,32'd1500,32'd1512,32'd1524,32'd1536,32'd1548,32'd1560,32'd1572,32'd1584,32'd1596,32'd1608,32'd1620,32'd1632,32'd1644,32'd1656,32'd1668,32'd1680,32'd1692,32'd1704,32'd1716,32'd1728,32'd1740,32'd1752,32'd1764,32'd1776,32'd1788,32'd1800,32'd1812,32'd1824,32'd1836,32'd1848,32'd1860,32'd1872,32'd1884,32'd1896,32'd1908,32'd1920,32'd1932,32'd1944,32'd1956,32'd1968,32'd1980,32'd1992,32'd2004,32'd2016,32'd2028,32'd2040,32'd2052,32'd2064,32'd2076,32'd2088,32'd2100,32'd2112,32'd2124,32'd2136,32'd2148,32'd2160,32'd2172,32'd2184,32'd2196,32'd2208,32'd2220,32'd2232,32'd2244,32'd2256,32'd2268,32'd2280,32'd2292,32'd2304,32'd2316,32'd2328,32'd2340,32'd2352,32'd2364,32'd2376,32'd2388,32'd2400,32'd2412,32'd2424,32'd2436,32'd2448,32'd2460,32'd2472,32'd2484,32'd2496,32'd2508,32'd2520,32'd2532,32'd2544,32'd2556,32'd2568,32'd2580,32'd2592,32'd2604,32'd2616,32'd2628,32'd2640,32'd2652,32'd2664,32'd2676,32'd2688,32'd2700,32'd2712,32'd2724,32'd2736,32'd2748,32'd2760,32'd2772,32'd2784,32'd2796,32'd2808,32'd2820,32'd2832,32'd2844,32'd2856,32'd2868,32'd2880,32'd2892,32'd2904,32'd2916,32'd2928,32'd2940,32'd2952,32'd2964,32'd2976,32'd2988,32'd3000,32'd3012,32'd3024,32'd3036,32'd3048,32'd3060,32'd3072,32'd3084,32'd3096,32'd3108,32'd3120,32'd3132,32'd3144,32'd3156,32'd3168,32'd3180,32'd3192,32'd3204,32'd3216,32'd3228,32'd3240,32'd3252,32'd3264,32'd3276,32'd3288,32'd3300,32'd3312,32'd3324,32'd3336,32'd3348,32'd3360,32'd3372,32'd3384,32'd3396,32'd3408,32'd3420,32'd3432,32'd3444,32'd3456,32'd3468,32'd3480,32'd3492,32'd3504,32'd3516,32'd3528,32'd3540,32'd3552,32'd3564,32'd3576,32'd3588,32'd3600,32'd3612,32'd3624,32'd3636,32'd3648,32'd3660,32'd3672,32'd3684,32'd3696,32'd3708,32'd3720,32'd3732,32'd3744,32'd3756,32'd3768,32'd3780,32'd3792,32'd3804,32'd3816,32'd3828,32'd3840,32'd3852,32'd3864,32'd3876,32'd3888,32'd3900,32'd3912,32'd3924,32'd3936,32'd3948,32'd3960,32'd3972,32'd3984,32'd3996,32'd4008,32'd4020,32'd4032,32'd4044,32'd4056,32'd4068,32'd4080,32'd4092,32'd4104,32'd4116,32'd4128,32'd4140,32'd4152,32'd4164,32'd4176,32'd4188,32'd4200,32'd4212,32'd4224,32'd4236,32'd4248,32'd4260,32'd4272,32'd4284,32'd4296,32'd4308,32'd4320,32'd4332,32'd4344,32'd4356,32'd4368,32'd4380,32'd4392,32'd4404,32'd4416,32'd4428,32'd4440,32'd4452,32'd4464,32'd4476,32'd4488,32'd4500,32'd4512,32'd4524,32'd4536,32'd4548,32'd4560,32'd4572,32'd4584,32'd4596,32'd4608,32'd4620,32'd4632,32'd4644,32'd4656,32'd4668,32'd4680,32'd4692,32'd4704,32'd4716,32'd4728,32'd4740,32'd4752,32'd4764,32'd4776,32'd4788 };matrix[13]='{32'd0,32'd13,32'd26,32'd39,32'd52,32'd65,32'd78,32'd91,32'd104,32'd117,32'd130,32'd143,32'd156,32'd169,32'd182,32'd195,32'd208,32'd221,32'd234,32'd247,32'd260,32'd273,32'd286,32'd299,32'd312,32'd325,32'd338,32'd351,32'd364,32'd377,32'd390,32'd403,32'd416,32'd429,32'd442,32'd455,32'd468,32'd481,32'd494,32'd507,32'd520,32'd533,32'd546,32'd559,32'd572,32'd585,32'd598,32'd611,32'd624,32'd637,32'd650,32'd663,32'd676,32'd689,32'd702,32'd715,32'd728,32'd741,32'd754,32'd767,32'd780,32'd793,32'd806,32'd819,32'd832,32'd845,32'd858,32'd871,32'd884,32'd897,32'd910,32'd923,32'd936,32'd949,32'd962,32'd975,32'd988,32'd1001,32'd1014,32'd1027,32'd1040,32'd1053,32'd1066,32'd1079,32'd1092,32'd1105,32'd1118,32'd1131,32'd1144,32'd1157,32'd1170,32'd1183,32'd1196,32'd1209,32'd1222,32'd1235,32'd1248,32'd1261,32'd1274,32'd1287,32'd1300,32'd1313,32'd1326,32'd1339,32'd1352,32'd1365,32'd1378,32'd1391,32'd1404,32'd1417,32'd1430,32'd1443,32'd1456,32'd1469,32'd1482,32'd1495,32'd1508,32'd1521,32'd1534,32'd1547,32'd1560,32'd1573,32'd1586,32'd1599,32'd1612,32'd1625,32'd1638,32'd1651,32'd1664,32'd1677,32'd1690,32'd1703,32'd1716,32'd1729,32'd1742,32'd1755,32'd1768,32'd1781,32'd1794,32'd1807,32'd1820,32'd1833,32'd1846,32'd1859,32'd1872,32'd1885,32'd1898,32'd1911,32'd1924,32'd1937,32'd1950,32'd1963,32'd1976,32'd1989,32'd2002,32'd2015,32'd2028,32'd2041,32'd2054,32'd2067,32'd2080,32'd2093,32'd2106,32'd2119,32'd2132,32'd2145,32'd2158,32'd2171,32'd2184,32'd2197,32'd2210,32'd2223,32'd2236,32'd2249,32'd2262,32'd2275,32'd2288,32'd2301,32'd2314,32'd2327,32'd2340,32'd2353,32'd2366,32'd2379,32'd2392,32'd2405,32'd2418,32'd2431,32'd2444,32'd2457,32'd2470,32'd2483,32'd2496,32'd2509,32'd2522,32'd2535,32'd2548,32'd2561,32'd2574,32'd2587,32'd2600,32'd2613,32'd2626,32'd2639,32'd2652,32'd2665,32'd2678,32'd2691,32'd2704,32'd2717,32'd2730,32'd2743,32'd2756,32'd2769,32'd2782,32'd2795,32'd2808,32'd2821,32'd2834,32'd2847,32'd2860,32'd2873,32'd2886,32'd2899,32'd2912,32'd2925,32'd2938,32'd2951,32'd2964,32'd2977,32'd2990,32'd3003,32'd3016,32'd3029,32'd3042,32'd3055,32'd3068,32'd3081,32'd3094,32'd3107,32'd3120,32'd3133,32'd3146,32'd3159,32'd3172,32'd3185,32'd3198,32'd3211,32'd3224,32'd3237,32'd3250,32'd3263,32'd3276,32'd3289,32'd3302,32'd3315,32'd3328,32'd3341,32'd3354,32'd3367,32'd3380,32'd3393,32'd3406,32'd3419,32'd3432,32'd3445,32'd3458,32'd3471,32'd3484,32'd3497,32'd3510,32'd3523,32'd3536,32'd3549,32'd3562,32'd3575,32'd3588,32'd3601,32'd3614,32'd3627,32'd3640,32'd3653,32'd3666,32'd3679,32'd3692,32'd3705,32'd3718,32'd3731,32'd3744,32'd3757,32'd3770,32'd3783,32'd3796,32'd3809,32'd3822,32'd3835,32'd3848,32'd3861,32'd3874,32'd3887,32'd3900,32'd3913,32'd3926,32'd3939,32'd3952,32'd3965,32'd3978,32'd3991,32'd4004,32'd4017,32'd4030,32'd4043,32'd4056,32'd4069,32'd4082,32'd4095,32'd4108,32'd4121,32'd4134,32'd4147,32'd4160,32'd4173,32'd4186,32'd4199,32'd4212,32'd4225,32'd4238,32'd4251,32'd4264,32'd4277,32'd4290,32'd4303,32'd4316,32'd4329,32'd4342,32'd4355,32'd4368,32'd4381,32'd4394,32'd4407,32'd4420,32'd4433,32'd4446,32'd4459,32'd4472,32'd4485,32'd4498,32'd4511,32'd4524,32'd4537,32'd4550,32'd4563,32'd4576,32'd4589,32'd4602,32'd4615,32'd4628,32'd4641,32'd4654,32'd4667,32'd4680,32'd4693,32'd4706,32'd4719,32'd4732,32'd4745,32'd4758,32'd4771,32'd4784,32'd4797,32'd4810,32'd4823,32'd4836,32'd4849,32'd4862,32'd4875,32'd4888,32'd4901,32'd4914,32'd4927,32'd4940,32'd4953,32'd4966,32'd4979,32'd4992,32'd5005,32'd5018,32'd5031,32'd5044,32'd5057,32'd5070,32'd5083,32'd5096,32'd5109,32'd5122,32'd5135,32'd5148,32'd5161,32'd5174,32'd5187 };matrix[14]='{32'd0,32'd14,32'd28,32'd42,32'd56,32'd70,32'd84,32'd98,32'd112,32'd126,32'd140,32'd154,32'd168,32'd182,32'd196,32'd210,32'd224,32'd238,32'd252,32'd266,32'd280,32'd294,32'd308,32'd322,32'd336,32'd350,32'd364,32'd378,32'd392,32'd406,32'd420,32'd434,32'd448,32'd462,32'd476,32'd490,32'd504,32'd518,32'd532,32'd546,32'd560,32'd574,32'd588,32'd602,32'd616,32'd630,32'd644,32'd658,32'd672,32'd686,32'd700,32'd714,32'd728,32'd742,32'd756,32'd770,32'd784,32'd798,32'd812,32'd826,32'd840,32'd854,32'd868,32'd882,32'd896,32'd910,32'd924,32'd938,32'd952,32'd966,32'd980,32'd994,32'd1008,32'd1022,32'd1036,32'd1050,32'd1064,32'd1078,32'd1092,32'd1106,32'd1120,32'd1134,32'd1148,32'd1162,32'd1176,32'd1190,32'd1204,32'd1218,32'd1232,32'd1246,32'd1260,32'd1274,32'd1288,32'd1302,32'd1316,32'd1330,32'd1344,32'd1358,32'd1372,32'd1386,32'd1400,32'd1414,32'd1428,32'd1442,32'd1456,32'd1470,32'd1484,32'd1498,32'd1512,32'd1526,32'd1540,32'd1554,32'd1568,32'd1582,32'd1596,32'd1610,32'd1624,32'd1638,32'd1652,32'd1666,32'd1680,32'd1694,32'd1708,32'd1722,32'd1736,32'd1750,32'd1764,32'd1778,32'd1792,32'd1806,32'd1820,32'd1834,32'd1848,32'd1862,32'd1876,32'd1890,32'd1904,32'd1918,32'd1932,32'd1946,32'd1960,32'd1974,32'd1988,32'd2002,32'd2016,32'd2030,32'd2044,32'd2058,32'd2072,32'd2086,32'd2100,32'd2114,32'd2128,32'd2142,32'd2156,32'd2170,32'd2184,32'd2198,32'd2212,32'd2226,32'd2240,32'd2254,32'd2268,32'd2282,32'd2296,32'd2310,32'd2324,32'd2338,32'd2352,32'd2366,32'd2380,32'd2394,32'd2408,32'd2422,32'd2436,32'd2450,32'd2464,32'd2478,32'd2492,32'd2506,32'd2520,32'd2534,32'd2548,32'd2562,32'd2576,32'd2590,32'd2604,32'd2618,32'd2632,32'd2646,32'd2660,32'd2674,32'd2688,32'd2702,32'd2716,32'd2730,32'd2744,32'd2758,32'd2772,32'd2786,32'd2800,32'd2814,32'd2828,32'd2842,32'd2856,32'd2870,32'd2884,32'd2898,32'd2912,32'd2926,32'd2940,32'd2954,32'd2968,32'd2982,32'd2996,32'd3010,32'd3024,32'd3038,32'd3052,32'd3066,32'd3080,32'd3094,32'd3108,32'd3122,32'd3136,32'd3150,32'd3164,32'd3178,32'd3192,32'd3206,32'd3220,32'd3234,32'd3248,32'd3262,32'd3276,32'd3290,32'd3304,32'd3318,32'd3332,32'd3346,32'd3360,32'd3374,32'd3388,32'd3402,32'd3416,32'd3430,32'd3444,32'd3458,32'd3472,32'd3486,32'd3500,32'd3514,32'd3528,32'd3542,32'd3556,32'd3570,32'd3584,32'd3598,32'd3612,32'd3626,32'd3640,32'd3654,32'd3668,32'd3682,32'd3696,32'd3710,32'd3724,32'd3738,32'd3752,32'd3766,32'd3780,32'd3794,32'd3808,32'd3822,32'd3836,32'd3850,32'd3864,32'd3878,32'd3892,32'd3906,32'd3920,32'd3934,32'd3948,32'd3962,32'd3976,32'd3990,32'd4004,32'd4018,32'd4032,32'd4046,32'd4060,32'd4074,32'd4088,32'd4102,32'd4116,32'd4130,32'd4144,32'd4158,32'd4172,32'd4186,32'd4200,32'd4214,32'd4228,32'd4242,32'd4256,32'd4270,32'd4284,32'd4298,32'd4312,32'd4326,32'd4340,32'd4354,32'd4368,32'd4382,32'd4396,32'd4410,32'd4424,32'd4438,32'd4452,32'd4466,32'd4480,32'd4494,32'd4508,32'd4522,32'd4536,32'd4550,32'd4564,32'd4578,32'd4592,32'd4606,32'd4620,32'd4634,32'd4648,32'd4662,32'd4676,32'd4690,32'd4704,32'd4718,32'd4732,32'd4746,32'd4760,32'd4774,32'd4788,32'd4802,32'd4816,32'd4830,32'd4844,32'd4858,32'd4872,32'd4886,32'd4900,32'd4914,32'd4928,32'd4942,32'd4956,32'd4970,32'd4984,32'd4998,32'd5012,32'd5026,32'd5040,32'd5054,32'd5068,32'd5082,32'd5096,32'd5110,32'd5124,32'd5138,32'd5152,32'd5166,32'd5180,32'd5194,32'd5208,32'd5222,32'd5236,32'd5250,32'd5264,32'd5278,32'd5292,32'd5306,32'd5320,32'd5334,32'd5348,32'd5362,32'd5376,32'd5390,32'd5404,32'd5418,32'd5432,32'd5446,32'd5460,32'd5474,32'd5488,32'd5502,32'd5516,32'd5530,32'd5544,32'd5558,32'd5572,32'd5586 };matrix[15]='{32'd0,32'd15,32'd30,32'd45,32'd60,32'd75,32'd90,32'd105,32'd120,32'd135,32'd150,32'd165,32'd180,32'd195,32'd210,32'd225,32'd240,32'd255,32'd270,32'd285,32'd300,32'd315,32'd330,32'd345,32'd360,32'd375,32'd390,32'd405,32'd420,32'd435,32'd450,32'd465,32'd480,32'd495,32'd510,32'd525,32'd540,32'd555,32'd570,32'd585,32'd600,32'd615,32'd630,32'd645,32'd660,32'd675,32'd690,32'd705,32'd720,32'd735,32'd750,32'd765,32'd780,32'd795,32'd810,32'd825,32'd840,32'd855,32'd870,32'd885,32'd900,32'd915,32'd930,32'd945,32'd960,32'd975,32'd990,32'd1005,32'd1020,32'd1035,32'd1050,32'd1065,32'd1080,32'd1095,32'd1110,32'd1125,32'd1140,32'd1155,32'd1170,32'd1185,32'd1200,32'd1215,32'd1230,32'd1245,32'd1260,32'd1275,32'd1290,32'd1305,32'd1320,32'd1335,32'd1350,32'd1365,32'd1380,32'd1395,32'd1410,32'd1425,32'd1440,32'd1455,32'd1470,32'd1485,32'd1500,32'd1515,32'd1530,32'd1545,32'd1560,32'd1575,32'd1590,32'd1605,32'd1620,32'd1635,32'd1650,32'd1665,32'd1680,32'd1695,32'd1710,32'd1725,32'd1740,32'd1755,32'd1770,32'd1785,32'd1800,32'd1815,32'd1830,32'd1845,32'd1860,32'd1875,32'd1890,32'd1905,32'd1920,32'd1935,32'd1950,32'd1965,32'd1980,32'd1995,32'd2010,32'd2025,32'd2040,32'd2055,32'd2070,32'd2085,32'd2100,32'd2115,32'd2130,32'd2145,32'd2160,32'd2175,32'd2190,32'd2205,32'd2220,32'd2235,32'd2250,32'd2265,32'd2280,32'd2295,32'd2310,32'd2325,32'd2340,32'd2355,32'd2370,32'd2385,32'd2400,32'd2415,32'd2430,32'd2445,32'd2460,32'd2475,32'd2490,32'd2505,32'd2520,32'd2535,32'd2550,32'd2565,32'd2580,32'd2595,32'd2610,32'd2625,32'd2640,32'd2655,32'd2670,32'd2685,32'd2700,32'd2715,32'd2730,32'd2745,32'd2760,32'd2775,32'd2790,32'd2805,32'd2820,32'd2835,32'd2850,32'd2865,32'd2880,32'd2895,32'd2910,32'd2925,32'd2940,32'd2955,32'd2970,32'd2985,32'd3000,32'd3015,32'd3030,32'd3045,32'd3060,32'd3075,32'd3090,32'd3105,32'd3120,32'd3135,32'd3150,32'd3165,32'd3180,32'd3195,32'd3210,32'd3225,32'd3240,32'd3255,32'd3270,32'd3285,32'd3300,32'd3315,32'd3330,32'd3345,32'd3360,32'd3375,32'd3390,32'd3405,32'd3420,32'd3435,32'd3450,32'd3465,32'd3480,32'd3495,32'd3510,32'd3525,32'd3540,32'd3555,32'd3570,32'd3585,32'd3600,32'd3615,32'd3630,32'd3645,32'd3660,32'd3675,32'd3690,32'd3705,32'd3720,32'd3735,32'd3750,32'd3765,32'd3780,32'd3795,32'd3810,32'd3825,32'd3840,32'd3855,32'd3870,32'd3885,32'd3900,32'd3915,32'd3930,32'd3945,32'd3960,32'd3975,32'd3990,32'd4005,32'd4020,32'd4035,32'd4050,32'd4065,32'd4080,32'd4095,32'd4110,32'd4125,32'd4140,32'd4155,32'd4170,32'd4185,32'd4200,32'd4215,32'd4230,32'd4245,32'd4260,32'd4275,32'd4290,32'd4305,32'd4320,32'd4335,32'd4350,32'd4365,32'd4380,32'd4395,32'd4410,32'd4425,32'd4440,32'd4455,32'd4470,32'd4485,32'd4500,32'd4515,32'd4530,32'd4545,32'd4560,32'd4575,32'd4590,32'd4605,32'd4620,32'd4635,32'd4650,32'd4665,32'd4680,32'd4695,32'd4710,32'd4725,32'd4740,32'd4755,32'd4770,32'd4785,32'd4800,32'd4815,32'd4830,32'd4845,32'd4860,32'd4875,32'd4890,32'd4905,32'd4920,32'd4935,32'd4950,32'd4965,32'd4980,32'd4995,32'd5010,32'd5025,32'd5040,32'd5055,32'd5070,32'd5085,32'd5100,32'd5115,32'd5130,32'd5145,32'd5160,32'd5175,32'd5190,32'd5205,32'd5220,32'd5235,32'd5250,32'd5265,32'd5280,32'd5295,32'd5310,32'd5325,32'd5340,32'd5355,32'd5370,32'd5385,32'd5400,32'd5415,32'd5430,32'd5445,32'd5460,32'd5475,32'd5490,32'd5505,32'd5520,32'd5535,32'd5550,32'd5565,32'd5580,32'd5595,32'd5610,32'd5625,32'd5640,32'd5655,32'd5670,32'd5685,32'd5700,32'd5715,32'd5730,32'd5745,32'd5760,32'd5775,32'd5790,32'd5805,32'd5820,32'd5835,32'd5850,32'd5865,32'd5880,32'd5895,32'd5910,32'd5925,32'd5940,32'd5955,32'd5970,32'd5985 };matrix[16]='{32'd0,32'd16,32'd32,32'd48,32'd64,32'd80,32'd96,32'd112,32'd128,32'd144,32'd160,32'd176,32'd192,32'd208,32'd224,32'd240,32'd256,32'd272,32'd288,32'd304,32'd320,32'd336,32'd352,32'd368,32'd384,32'd400,32'd416,32'd432,32'd448,32'd464,32'd480,32'd496,32'd512,32'd528,32'd544,32'd560,32'd576,32'd592,32'd608,32'd624,32'd640,32'd656,32'd672,32'd688,32'd704,32'd720,32'd736,32'd752,32'd768,32'd784,32'd800,32'd816,32'd832,32'd848,32'd864,32'd880,32'd896,32'd912,32'd928,32'd944,32'd960,32'd976,32'd992,32'd1008,32'd1024,32'd1040,32'd1056,32'd1072,32'd1088,32'd1104,32'd1120,32'd1136,32'd1152,32'd1168,32'd1184,32'd1200,32'd1216,32'd1232,32'd1248,32'd1264,32'd1280,32'd1296,32'd1312,32'd1328,32'd1344,32'd1360,32'd1376,32'd1392,32'd1408,32'd1424,32'd1440,32'd1456,32'd1472,32'd1488,32'd1504,32'd1520,32'd1536,32'd1552,32'd1568,32'd1584,32'd1600,32'd1616,32'd1632,32'd1648,32'd1664,32'd1680,32'd1696,32'd1712,32'd1728,32'd1744,32'd1760,32'd1776,32'd1792,32'd1808,32'd1824,32'd1840,32'd1856,32'd1872,32'd1888,32'd1904,32'd1920,32'd1936,32'd1952,32'd1968,32'd1984,32'd2000,32'd2016,32'd2032,32'd2048,32'd2064,32'd2080,32'd2096,32'd2112,32'd2128,32'd2144,32'd2160,32'd2176,32'd2192,32'd2208,32'd2224,32'd2240,32'd2256,32'd2272,32'd2288,32'd2304,32'd2320,32'd2336,32'd2352,32'd2368,32'd2384,32'd2400,32'd2416,32'd2432,32'd2448,32'd2464,32'd2480,32'd2496,32'd2512,32'd2528,32'd2544,32'd2560,32'd2576,32'd2592,32'd2608,32'd2624,32'd2640,32'd2656,32'd2672,32'd2688,32'd2704,32'd2720,32'd2736,32'd2752,32'd2768,32'd2784,32'd2800,32'd2816,32'd2832,32'd2848,32'd2864,32'd2880,32'd2896,32'd2912,32'd2928,32'd2944,32'd2960,32'd2976,32'd2992,32'd3008,32'd3024,32'd3040,32'd3056,32'd3072,32'd3088,32'd3104,32'd3120,32'd3136,32'd3152,32'd3168,32'd3184,32'd3200,32'd3216,32'd3232,32'd3248,32'd3264,32'd3280,32'd3296,32'd3312,32'd3328,32'd3344,32'd3360,32'd3376,32'd3392,32'd3408,32'd3424,32'd3440,32'd3456,32'd3472,32'd3488,32'd3504,32'd3520,32'd3536,32'd3552,32'd3568,32'd3584,32'd3600,32'd3616,32'd3632,32'd3648,32'd3664,32'd3680,32'd3696,32'd3712,32'd3728,32'd3744,32'd3760,32'd3776,32'd3792,32'd3808,32'd3824,32'd3840,32'd3856,32'd3872,32'd3888,32'd3904,32'd3920,32'd3936,32'd3952,32'd3968,32'd3984,32'd4000,32'd4016,32'd4032,32'd4048,32'd4064,32'd4080,32'd4096,32'd4112,32'd4128,32'd4144,32'd4160,32'd4176,32'd4192,32'd4208,32'd4224,32'd4240,32'd4256,32'd4272,32'd4288,32'd4304,32'd4320,32'd4336,32'd4352,32'd4368,32'd4384,32'd4400,32'd4416,32'd4432,32'd4448,32'd4464,32'd4480,32'd4496,32'd4512,32'd4528,32'd4544,32'd4560,32'd4576,32'd4592,32'd4608,32'd4624,32'd4640,32'd4656,32'd4672,32'd4688,32'd4704,32'd4720,32'd4736,32'd4752,32'd4768,32'd4784,32'd4800,32'd4816,32'd4832,32'd4848,32'd4864,32'd4880,32'd4896,32'd4912,32'd4928,32'd4944,32'd4960,32'd4976,32'd4992,32'd5008,32'd5024,32'd5040,32'd5056,32'd5072,32'd5088,32'd5104,32'd5120,32'd5136,32'd5152,32'd5168,32'd5184,32'd5200,32'd5216,32'd5232,32'd5248,32'd5264,32'd5280,32'd5296,32'd5312,32'd5328,32'd5344,32'd5360,32'd5376,32'd5392,32'd5408,32'd5424,32'd5440,32'd5456,32'd5472,32'd5488,32'd5504,32'd5520,32'd5536,32'd5552,32'd5568,32'd5584,32'd5600,32'd5616,32'd5632,32'd5648,32'd5664,32'd5680,32'd5696,32'd5712,32'd5728,32'd5744,32'd5760,32'd5776,32'd5792,32'd5808,32'd5824,32'd5840,32'd5856,32'd5872,32'd5888,32'd5904,32'd5920,32'd5936,32'd5952,32'd5968,32'd5984,32'd6000,32'd6016,32'd6032,32'd6048,32'd6064,32'd6080,32'd6096,32'd6112,32'd6128,32'd6144,32'd6160,32'd6176,32'd6192,32'd6208,32'd6224,32'd6240,32'd6256,32'd6272,32'd6288,32'd6304,32'd6320,32'd6336,32'd6352,32'd6368,32'd6384 };matrix[17]='{32'd0,32'd17,32'd34,32'd51,32'd68,32'd85,32'd102,32'd119,32'd136,32'd153,32'd170,32'd187,32'd204,32'd221,32'd238,32'd255,32'd272,32'd289,32'd306,32'd323,32'd340,32'd357,32'd374,32'd391,32'd408,32'd425,32'd442,32'd459,32'd476,32'd493,32'd510,32'd527,32'd544,32'd561,32'd578,32'd595,32'd612,32'd629,32'd646,32'd663,32'd680,32'd697,32'd714,32'd731,32'd748,32'd765,32'd782,32'd799,32'd816,32'd833,32'd850,32'd867,32'd884,32'd901,32'd918,32'd935,32'd952,32'd969,32'd986,32'd1003,32'd1020,32'd1037,32'd1054,32'd1071,32'd1088,32'd1105,32'd1122,32'd1139,32'd1156,32'd1173,32'd1190,32'd1207,32'd1224,32'd1241,32'd1258,32'd1275,32'd1292,32'd1309,32'd1326,32'd1343,32'd1360,32'd1377,32'd1394,32'd1411,32'd1428,32'd1445,32'd1462,32'd1479,32'd1496,32'd1513,32'd1530,32'd1547,32'd1564,32'd1581,32'd1598,32'd1615,32'd1632,32'd1649,32'd1666,32'd1683,32'd1700,32'd1717,32'd1734,32'd1751,32'd1768,32'd1785,32'd1802,32'd1819,32'd1836,32'd1853,32'd1870,32'd1887,32'd1904,32'd1921,32'd1938,32'd1955,32'd1972,32'd1989,32'd2006,32'd2023,32'd2040,32'd2057,32'd2074,32'd2091,32'd2108,32'd2125,32'd2142,32'd2159,32'd2176,32'd2193,32'd2210,32'd2227,32'd2244,32'd2261,32'd2278,32'd2295,32'd2312,32'd2329,32'd2346,32'd2363,32'd2380,32'd2397,32'd2414,32'd2431,32'd2448,32'd2465,32'd2482,32'd2499,32'd2516,32'd2533,32'd2550,32'd2567,32'd2584,32'd2601,32'd2618,32'd2635,32'd2652,32'd2669,32'd2686,32'd2703,32'd2720,32'd2737,32'd2754,32'd2771,32'd2788,32'd2805,32'd2822,32'd2839,32'd2856,32'd2873,32'd2890,32'd2907,32'd2924,32'd2941,32'd2958,32'd2975,32'd2992,32'd3009,32'd3026,32'd3043,32'd3060,32'd3077,32'd3094,32'd3111,32'd3128,32'd3145,32'd3162,32'd3179,32'd3196,32'd3213,32'd3230,32'd3247,32'd3264,32'd3281,32'd3298,32'd3315,32'd3332,32'd3349,32'd3366,32'd3383,32'd3400,32'd3417,32'd3434,32'd3451,32'd3468,32'd3485,32'd3502,32'd3519,32'd3536,32'd3553,32'd3570,32'd3587,32'd3604,32'd3621,32'd3638,32'd3655,32'd3672,32'd3689,32'd3706,32'd3723,32'd3740,32'd3757,32'd3774,32'd3791,32'd3808,32'd3825,32'd3842,32'd3859,32'd3876,32'd3893,32'd3910,32'd3927,32'd3944,32'd3961,32'd3978,32'd3995,32'd4012,32'd4029,32'd4046,32'd4063,32'd4080,32'd4097,32'd4114,32'd4131,32'd4148,32'd4165,32'd4182,32'd4199,32'd4216,32'd4233,32'd4250,32'd4267,32'd4284,32'd4301,32'd4318,32'd4335,32'd4352,32'd4369,32'd4386,32'd4403,32'd4420,32'd4437,32'd4454,32'd4471,32'd4488,32'd4505,32'd4522,32'd4539,32'd4556,32'd4573,32'd4590,32'd4607,32'd4624,32'd4641,32'd4658,32'd4675,32'd4692,32'd4709,32'd4726,32'd4743,32'd4760,32'd4777,32'd4794,32'd4811,32'd4828,32'd4845,32'd4862,32'd4879,32'd4896,32'd4913,32'd4930,32'd4947,32'd4964,32'd4981,32'd4998,32'd5015,32'd5032,32'd5049,32'd5066,32'd5083,32'd5100,32'd5117,32'd5134,32'd5151,32'd5168,32'd5185,32'd5202,32'd5219,32'd5236,32'd5253,32'd5270,32'd5287,32'd5304,32'd5321,32'd5338,32'd5355,32'd5372,32'd5389,32'd5406,32'd5423,32'd5440,32'd5457,32'd5474,32'd5491,32'd5508,32'd5525,32'd5542,32'd5559,32'd5576,32'd5593,32'd5610,32'd5627,32'd5644,32'd5661,32'd5678,32'd5695,32'd5712,32'd5729,32'd5746,32'd5763,32'd5780,32'd5797,32'd5814,32'd5831,32'd5848,32'd5865,32'd5882,32'd5899,32'd5916,32'd5933,32'd5950,32'd5967,32'd5984,32'd6001,32'd6018,32'd6035,32'd6052,32'd6069,32'd6086,32'd6103,32'd6120,32'd6137,32'd6154,32'd6171,32'd6188,32'd6205,32'd6222,32'd6239,32'd6256,32'd6273,32'd6290,32'd6307,32'd6324,32'd6341,32'd6358,32'd6375,32'd6392,32'd6409,32'd6426,32'd6443,32'd6460,32'd6477,32'd6494,32'd6511,32'd6528,32'd6545,32'd6562,32'd6579,32'd6596,32'd6613,32'd6630,32'd6647,32'd6664,32'd6681,32'd6698,32'd6715,32'd6732,32'd6749,32'd6766,32'd6783 };matrix[18]='{32'd0,32'd18,32'd36,32'd54,32'd72,32'd90,32'd108,32'd126,32'd144,32'd162,32'd180,32'd198,32'd216,32'd234,32'd252,32'd270,32'd288,32'd306,32'd324,32'd342,32'd360,32'd378,32'd396,32'd414,32'd432,32'd450,32'd468,32'd486,32'd504,32'd522,32'd540,32'd558,32'd576,32'd594,32'd612,32'd630,32'd648,32'd666,32'd684,32'd702,32'd720,32'd738,32'd756,32'd774,32'd792,32'd810,32'd828,32'd846,32'd864,32'd882,32'd900,32'd918,32'd936,32'd954,32'd972,32'd990,32'd1008,32'd1026,32'd1044,32'd1062,32'd1080,32'd1098,32'd1116,32'd1134,32'd1152,32'd1170,32'd1188,32'd1206,32'd1224,32'd1242,32'd1260,32'd1278,32'd1296,32'd1314,32'd1332,32'd1350,32'd1368,32'd1386,32'd1404,32'd1422,32'd1440,32'd1458,32'd1476,32'd1494,32'd1512,32'd1530,32'd1548,32'd1566,32'd1584,32'd1602,32'd1620,32'd1638,32'd1656,32'd1674,32'd1692,32'd1710,32'd1728,32'd1746,32'd1764,32'd1782,32'd1800,32'd1818,32'd1836,32'd1854,32'd1872,32'd1890,32'd1908,32'd1926,32'd1944,32'd1962,32'd1980,32'd1998,32'd2016,32'd2034,32'd2052,32'd2070,32'd2088,32'd2106,32'd2124,32'd2142,32'd2160,32'd2178,32'd2196,32'd2214,32'd2232,32'd2250,32'd2268,32'd2286,32'd2304,32'd2322,32'd2340,32'd2358,32'd2376,32'd2394,32'd2412,32'd2430,32'd2448,32'd2466,32'd2484,32'd2502,32'd2520,32'd2538,32'd2556,32'd2574,32'd2592,32'd2610,32'd2628,32'd2646,32'd2664,32'd2682,32'd2700,32'd2718,32'd2736,32'd2754,32'd2772,32'd2790,32'd2808,32'd2826,32'd2844,32'd2862,32'd2880,32'd2898,32'd2916,32'd2934,32'd2952,32'd2970,32'd2988,32'd3006,32'd3024,32'd3042,32'd3060,32'd3078,32'd3096,32'd3114,32'd3132,32'd3150,32'd3168,32'd3186,32'd3204,32'd3222,32'd3240,32'd3258,32'd3276,32'd3294,32'd3312,32'd3330,32'd3348,32'd3366,32'd3384,32'd3402,32'd3420,32'd3438,32'd3456,32'd3474,32'd3492,32'd3510,32'd3528,32'd3546,32'd3564,32'd3582,32'd3600,32'd3618,32'd3636,32'd3654,32'd3672,32'd3690,32'd3708,32'd3726,32'd3744,32'd3762,32'd3780,32'd3798,32'd3816,32'd3834,32'd3852,32'd3870,32'd3888,32'd3906,32'd3924,32'd3942,32'd3960,32'd3978,32'd3996,32'd4014,32'd4032,32'd4050,32'd4068,32'd4086,32'd4104,32'd4122,32'd4140,32'd4158,32'd4176,32'd4194,32'd4212,32'd4230,32'd4248,32'd4266,32'd4284,32'd4302,32'd4320,32'd4338,32'd4356,32'd4374,32'd4392,32'd4410,32'd4428,32'd4446,32'd4464,32'd4482,32'd4500,32'd4518,32'd4536,32'd4554,32'd4572,32'd4590,32'd4608,32'd4626,32'd4644,32'd4662,32'd4680,32'd4698,32'd4716,32'd4734,32'd4752,32'd4770,32'd4788,32'd4806,32'd4824,32'd4842,32'd4860,32'd4878,32'd4896,32'd4914,32'd4932,32'd4950,32'd4968,32'd4986,32'd5004,32'd5022,32'd5040,32'd5058,32'd5076,32'd5094,32'd5112,32'd5130,32'd5148,32'd5166,32'd5184,32'd5202,32'd5220,32'd5238,32'd5256,32'd5274,32'd5292,32'd5310,32'd5328,32'd5346,32'd5364,32'd5382,32'd5400,32'd5418,32'd5436,32'd5454,32'd5472,32'd5490,32'd5508,32'd5526,32'd5544,32'd5562,32'd5580,32'd5598,32'd5616,32'd5634,32'd5652,32'd5670,32'd5688,32'd5706,32'd5724,32'd5742,32'd5760,32'd5778,32'd5796,32'd5814,32'd5832,32'd5850,32'd5868,32'd5886,32'd5904,32'd5922,32'd5940,32'd5958,32'd5976,32'd5994,32'd6012,32'd6030,32'd6048,32'd6066,32'd6084,32'd6102,32'd6120,32'd6138,32'd6156,32'd6174,32'd6192,32'd6210,32'd6228,32'd6246,32'd6264,32'd6282,32'd6300,32'd6318,32'd6336,32'd6354,32'd6372,32'd6390,32'd6408,32'd6426,32'd6444,32'd6462,32'd6480,32'd6498,32'd6516,32'd6534,32'd6552,32'd6570,32'd6588,32'd6606,32'd6624,32'd6642,32'd6660,32'd6678,32'd6696,32'd6714,32'd6732,32'd6750,32'd6768,32'd6786,32'd6804,32'd6822,32'd6840,32'd6858,32'd6876,32'd6894,32'd6912,32'd6930,32'd6948,32'd6966,32'd6984,32'd7002,32'd7020,32'd7038,32'd7056,32'd7074,32'd7092,32'd7110,32'd7128,32'd7146,32'd7164,32'd7182 };matrix[19]='{32'd0,32'd19,32'd38,32'd57,32'd76,32'd95,32'd114,32'd133,32'd152,32'd171,32'd190,32'd209,32'd228,32'd247,32'd266,32'd285,32'd304,32'd323,32'd342,32'd361,32'd380,32'd399,32'd418,32'd437,32'd456,32'd475,32'd494,32'd513,32'd532,32'd551,32'd570,32'd589,32'd608,32'd627,32'd646,32'd665,32'd684,32'd703,32'd722,32'd741,32'd760,32'd779,32'd798,32'd817,32'd836,32'd855,32'd874,32'd893,32'd912,32'd931,32'd950,32'd969,32'd988,32'd1007,32'd1026,32'd1045,32'd1064,32'd1083,32'd1102,32'd1121,32'd1140,32'd1159,32'd1178,32'd1197,32'd1216,32'd1235,32'd1254,32'd1273,32'd1292,32'd1311,32'd1330,32'd1349,32'd1368,32'd1387,32'd1406,32'd1425,32'd1444,32'd1463,32'd1482,32'd1501,32'd1520,32'd1539,32'd1558,32'd1577,32'd1596,32'd1615,32'd1634,32'd1653,32'd1672,32'd1691,32'd1710,32'd1729,32'd1748,32'd1767,32'd1786,32'd1805,32'd1824,32'd1843,32'd1862,32'd1881,32'd1900,32'd1919,32'd1938,32'd1957,32'd1976,32'd1995,32'd2014,32'd2033,32'd2052,32'd2071,32'd2090,32'd2109,32'd2128,32'd2147,32'd2166,32'd2185,32'd2204,32'd2223,32'd2242,32'd2261,32'd2280,32'd2299,32'd2318,32'd2337,32'd2356,32'd2375,32'd2394,32'd2413,32'd2432,32'd2451,32'd2470,32'd2489,32'd2508,32'd2527,32'd2546,32'd2565,32'd2584,32'd2603,32'd2622,32'd2641,32'd2660,32'd2679,32'd2698,32'd2717,32'd2736,32'd2755,32'd2774,32'd2793,32'd2812,32'd2831,32'd2850,32'd2869,32'd2888,32'd2907,32'd2926,32'd2945,32'd2964,32'd2983,32'd3002,32'd3021,32'd3040,32'd3059,32'd3078,32'd3097,32'd3116,32'd3135,32'd3154,32'd3173,32'd3192,32'd3211,32'd3230,32'd3249,32'd3268,32'd3287,32'd3306,32'd3325,32'd3344,32'd3363,32'd3382,32'd3401,32'd3420,32'd3439,32'd3458,32'd3477,32'd3496,32'd3515,32'd3534,32'd3553,32'd3572,32'd3591,32'd3610,32'd3629,32'd3648,32'd3667,32'd3686,32'd3705,32'd3724,32'd3743,32'd3762,32'd3781,32'd3800,32'd3819,32'd3838,32'd3857,32'd3876,32'd3895,32'd3914,32'd3933,32'd3952,32'd3971,32'd3990,32'd4009,32'd4028,32'd4047,32'd4066,32'd4085,32'd4104,32'd4123,32'd4142,32'd4161,32'd4180,32'd4199,32'd4218,32'd4237,32'd4256,32'd4275,32'd4294,32'd4313,32'd4332,32'd4351,32'd4370,32'd4389,32'd4408,32'd4427,32'd4446,32'd4465,32'd4484,32'd4503,32'd4522,32'd4541,32'd4560,32'd4579,32'd4598,32'd4617,32'd4636,32'd4655,32'd4674,32'd4693,32'd4712,32'd4731,32'd4750,32'd4769,32'd4788,32'd4807,32'd4826,32'd4845,32'd4864,32'd4883,32'd4902,32'd4921,32'd4940,32'd4959,32'd4978,32'd4997,32'd5016,32'd5035,32'd5054,32'd5073,32'd5092,32'd5111,32'd5130,32'd5149,32'd5168,32'd5187,32'd5206,32'd5225,32'd5244,32'd5263,32'd5282,32'd5301,32'd5320,32'd5339,32'd5358,32'd5377,32'd5396,32'd5415,32'd5434,32'd5453,32'd5472,32'd5491,32'd5510,32'd5529,32'd5548,32'd5567,32'd5586,32'd5605,32'd5624,32'd5643,32'd5662,32'd5681,32'd5700,32'd5719,32'd5738,32'd5757,32'd5776,32'd5795,32'd5814,32'd5833,32'd5852,32'd5871,32'd5890,32'd5909,32'd5928,32'd5947,32'd5966,32'd5985,32'd6004,32'd6023,32'd6042,32'd6061,32'd6080,32'd6099,32'd6118,32'd6137,32'd6156,32'd6175,32'd6194,32'd6213,32'd6232,32'd6251,32'd6270,32'd6289,32'd6308,32'd6327,32'd6346,32'd6365,32'd6384,32'd6403,32'd6422,32'd6441,32'd6460,32'd6479,32'd6498,32'd6517,32'd6536,32'd6555,32'd6574,32'd6593,32'd6612,32'd6631,32'd6650,32'd6669,32'd6688,32'd6707,32'd6726,32'd6745,32'd6764,32'd6783,32'd6802,32'd6821,32'd6840,32'd6859,32'd6878,32'd6897,32'd6916,32'd6935,32'd6954,32'd6973,32'd6992,32'd7011,32'd7030,32'd7049,32'd7068,32'd7087,32'd7106,32'd7125,32'd7144,32'd7163,32'd7182,32'd7201,32'd7220,32'd7239,32'd7258,32'd7277,32'd7296,32'd7315,32'd7334,32'd7353,32'd7372,32'd7391,32'd7410,32'd7429,32'd7448,32'd7467,32'd7486,32'd7505,32'd7524,32'd7543,32'd7562,32'd7581 };matrix[20]='{32'd0,32'd20,32'd40,32'd60,32'd80,32'd100,32'd120,32'd140,32'd160,32'd180,32'd200,32'd220,32'd240,32'd260,32'd280,32'd300,32'd320,32'd340,32'd360,32'd380,32'd400,32'd420,32'd440,32'd460,32'd480,32'd500,32'd520,32'd540,32'd560,32'd580,32'd600,32'd620,32'd640,32'd660,32'd680,32'd700,32'd720,32'd740,32'd760,32'd780,32'd800,32'd820,32'd840,32'd860,32'd880,32'd900,32'd920,32'd940,32'd960,32'd980,32'd1000,32'd1020,32'd1040,32'd1060,32'd1080,32'd1100,32'd1120,32'd1140,32'd1160,32'd1180,32'd1200,32'd1220,32'd1240,32'd1260,32'd1280,32'd1300,32'd1320,32'd1340,32'd1360,32'd1380,32'd1400,32'd1420,32'd1440,32'd1460,32'd1480,32'd1500,32'd1520,32'd1540,32'd1560,32'd1580,32'd1600,32'd1620,32'd1640,32'd1660,32'd1680,32'd1700,32'd1720,32'd1740,32'd1760,32'd1780,32'd1800,32'd1820,32'd1840,32'd1860,32'd1880,32'd1900,32'd1920,32'd1940,32'd1960,32'd1980,32'd2000,32'd2020,32'd2040,32'd2060,32'd2080,32'd2100,32'd2120,32'd2140,32'd2160,32'd2180,32'd2200,32'd2220,32'd2240,32'd2260,32'd2280,32'd2300,32'd2320,32'd2340,32'd2360,32'd2380,32'd2400,32'd2420,32'd2440,32'd2460,32'd2480,32'd2500,32'd2520,32'd2540,32'd2560,32'd2580,32'd2600,32'd2620,32'd2640,32'd2660,32'd2680,32'd2700,32'd2720,32'd2740,32'd2760,32'd2780,32'd2800,32'd2820,32'd2840,32'd2860,32'd2880,32'd2900,32'd2920,32'd2940,32'd2960,32'd2980,32'd3000,32'd3020,32'd3040,32'd3060,32'd3080,32'd3100,32'd3120,32'd3140,32'd3160,32'd3180,32'd3200,32'd3220,32'd3240,32'd3260,32'd3280,32'd3300,32'd3320,32'd3340,32'd3360,32'd3380,32'd3400,32'd3420,32'd3440,32'd3460,32'd3480,32'd3500,32'd3520,32'd3540,32'd3560,32'd3580,32'd3600,32'd3620,32'd3640,32'd3660,32'd3680,32'd3700,32'd3720,32'd3740,32'd3760,32'd3780,32'd3800,32'd3820,32'd3840,32'd3860,32'd3880,32'd3900,32'd3920,32'd3940,32'd3960,32'd3980,32'd4000,32'd4020,32'd4040,32'd4060,32'd4080,32'd4100,32'd4120,32'd4140,32'd4160,32'd4180,32'd4200,32'd4220,32'd4240,32'd4260,32'd4280,32'd4300,32'd4320,32'd4340,32'd4360,32'd4380,32'd4400,32'd4420,32'd4440,32'd4460,32'd4480,32'd4500,32'd4520,32'd4540,32'd4560,32'd4580,32'd4600,32'd4620,32'd4640,32'd4660,32'd4680,32'd4700,32'd4720,32'd4740,32'd4760,32'd4780,32'd4800,32'd4820,32'd4840,32'd4860,32'd4880,32'd4900,32'd4920,32'd4940,32'd4960,32'd4980,32'd5000,32'd5020,32'd5040,32'd5060,32'd5080,32'd5100,32'd5120,32'd5140,32'd5160,32'd5180,32'd5200,32'd5220,32'd5240,32'd5260,32'd5280,32'd5300,32'd5320,32'd5340,32'd5360,32'd5380,32'd5400,32'd5420,32'd5440,32'd5460,32'd5480,32'd5500,32'd5520,32'd5540,32'd5560,32'd5580,32'd5600,32'd5620,32'd5640,32'd5660,32'd5680,32'd5700,32'd5720,32'd5740,32'd5760,32'd5780,32'd5800,32'd5820,32'd5840,32'd5860,32'd5880,32'd5900,32'd5920,32'd5940,32'd5960,32'd5980,32'd6000,32'd6020,32'd6040,32'd6060,32'd6080,32'd6100,32'd6120,32'd6140,32'd6160,32'd6180,32'd6200,32'd6220,32'd6240,32'd6260,32'd6280,32'd6300,32'd6320,32'd6340,32'd6360,32'd6380,32'd6400,32'd6420,32'd6440,32'd6460,32'd6480,32'd6500,32'd6520,32'd6540,32'd6560,32'd6580,32'd6600,32'd6620,32'd6640,32'd6660,32'd6680,32'd6700,32'd6720,32'd6740,32'd6760,32'd6780,32'd6800,32'd6820,32'd6840,32'd6860,32'd6880,32'd6900,32'd6920,32'd6940,32'd6960,32'd6980,32'd7000,32'd7020,32'd7040,32'd7060,32'd7080,32'd7100,32'd7120,32'd7140,32'd7160,32'd7180,32'd7200,32'd7220,32'd7240,32'd7260,32'd7280,32'd7300,32'd7320,32'd7340,32'd7360,32'd7380,32'd7400,32'd7420,32'd7440,32'd7460,32'd7480,32'd7500,32'd7520,32'd7540,32'd7560,32'd7580,32'd7600,32'd7620,32'd7640,32'd7660,32'd7680,32'd7700,32'd7720,32'd7740,32'd7760,32'd7780,32'd7800,32'd7820,32'd7840,32'd7860,32'd7880,32'd7900,32'd7920,32'd7940,32'd7960,32'd7980 };matrix[21]='{32'd0,32'd21,32'd42,32'd63,32'd84,32'd105,32'd126,32'd147,32'd168,32'd189,32'd210,32'd231,32'd252,32'd273,32'd294,32'd315,32'd336,32'd357,32'd378,32'd399,32'd420,32'd441,32'd462,32'd483,32'd504,32'd525,32'd546,32'd567,32'd588,32'd609,32'd630,32'd651,32'd672,32'd693,32'd714,32'd735,32'd756,32'd777,32'd798,32'd819,32'd840,32'd861,32'd882,32'd903,32'd924,32'd945,32'd966,32'd987,32'd1008,32'd1029,32'd1050,32'd1071,32'd1092,32'd1113,32'd1134,32'd1155,32'd1176,32'd1197,32'd1218,32'd1239,32'd1260,32'd1281,32'd1302,32'd1323,32'd1344,32'd1365,32'd1386,32'd1407,32'd1428,32'd1449,32'd1470,32'd1491,32'd1512,32'd1533,32'd1554,32'd1575,32'd1596,32'd1617,32'd1638,32'd1659,32'd1680,32'd1701,32'd1722,32'd1743,32'd1764,32'd1785,32'd1806,32'd1827,32'd1848,32'd1869,32'd1890,32'd1911,32'd1932,32'd1953,32'd1974,32'd1995,32'd2016,32'd2037,32'd2058,32'd2079,32'd2100,32'd2121,32'd2142,32'd2163,32'd2184,32'd2205,32'd2226,32'd2247,32'd2268,32'd2289,32'd2310,32'd2331,32'd2352,32'd2373,32'd2394,32'd2415,32'd2436,32'd2457,32'd2478,32'd2499,32'd2520,32'd2541,32'd2562,32'd2583,32'd2604,32'd2625,32'd2646,32'd2667,32'd2688,32'd2709,32'd2730,32'd2751,32'd2772,32'd2793,32'd2814,32'd2835,32'd2856,32'd2877,32'd2898,32'd2919,32'd2940,32'd2961,32'd2982,32'd3003,32'd3024,32'd3045,32'd3066,32'd3087,32'd3108,32'd3129,32'd3150,32'd3171,32'd3192,32'd3213,32'd3234,32'd3255,32'd3276,32'd3297,32'd3318,32'd3339,32'd3360,32'd3381,32'd3402,32'd3423,32'd3444,32'd3465,32'd3486,32'd3507,32'd3528,32'd3549,32'd3570,32'd3591,32'd3612,32'd3633,32'd3654,32'd3675,32'd3696,32'd3717,32'd3738,32'd3759,32'd3780,32'd3801,32'd3822,32'd3843,32'd3864,32'd3885,32'd3906,32'd3927,32'd3948,32'd3969,32'd3990,32'd4011,32'd4032,32'd4053,32'd4074,32'd4095,32'd4116,32'd4137,32'd4158,32'd4179,32'd4200,32'd4221,32'd4242,32'd4263,32'd4284,32'd4305,32'd4326,32'd4347,32'd4368,32'd4389,32'd4410,32'd4431,32'd4452,32'd4473,32'd4494,32'd4515,32'd4536,32'd4557,32'd4578,32'd4599,32'd4620,32'd4641,32'd4662,32'd4683,32'd4704,32'd4725,32'd4746,32'd4767,32'd4788,32'd4809,32'd4830,32'd4851,32'd4872,32'd4893,32'd4914,32'd4935,32'd4956,32'd4977,32'd4998,32'd5019,32'd5040,32'd5061,32'd5082,32'd5103,32'd5124,32'd5145,32'd5166,32'd5187,32'd5208,32'd5229,32'd5250,32'd5271,32'd5292,32'd5313,32'd5334,32'd5355,32'd5376,32'd5397,32'd5418,32'd5439,32'd5460,32'd5481,32'd5502,32'd5523,32'd5544,32'd5565,32'd5586,32'd5607,32'd5628,32'd5649,32'd5670,32'd5691,32'd5712,32'd5733,32'd5754,32'd5775,32'd5796,32'd5817,32'd5838,32'd5859,32'd5880,32'd5901,32'd5922,32'd5943,32'd5964,32'd5985,32'd6006,32'd6027,32'd6048,32'd6069,32'd6090,32'd6111,32'd6132,32'd6153,32'd6174,32'd6195,32'd6216,32'd6237,32'd6258,32'd6279,32'd6300,32'd6321,32'd6342,32'd6363,32'd6384,32'd6405,32'd6426,32'd6447,32'd6468,32'd6489,32'd6510,32'd6531,32'd6552,32'd6573,32'd6594,32'd6615,32'd6636,32'd6657,32'd6678,32'd6699,32'd6720,32'd6741,32'd6762,32'd6783,32'd6804,32'd6825,32'd6846,32'd6867,32'd6888,32'd6909,32'd6930,32'd6951,32'd6972,32'd6993,32'd7014,32'd7035,32'd7056,32'd7077,32'd7098,32'd7119,32'd7140,32'd7161,32'd7182,32'd7203,32'd7224,32'd7245,32'd7266,32'd7287,32'd7308,32'd7329,32'd7350,32'd7371,32'd7392,32'd7413,32'd7434,32'd7455,32'd7476,32'd7497,32'd7518,32'd7539,32'd7560,32'd7581,32'd7602,32'd7623,32'd7644,32'd7665,32'd7686,32'd7707,32'd7728,32'd7749,32'd7770,32'd7791,32'd7812,32'd7833,32'd7854,32'd7875,32'd7896,32'd7917,32'd7938,32'd7959,32'd7980,32'd8001,32'd8022,32'd8043,32'd8064,32'd8085,32'd8106,32'd8127,32'd8148,32'd8169,32'd8190,32'd8211,32'd8232,32'd8253,32'd8274,32'd8295,32'd8316,32'd8337,32'd8358,32'd8379 };matrix[22]='{32'd0,32'd22,32'd44,32'd66,32'd88,32'd110,32'd132,32'd154,32'd176,32'd198,32'd220,32'd242,32'd264,32'd286,32'd308,32'd330,32'd352,32'd374,32'd396,32'd418,32'd440,32'd462,32'd484,32'd506,32'd528,32'd550,32'd572,32'd594,32'd616,32'd638,32'd660,32'd682,32'd704,32'd726,32'd748,32'd770,32'd792,32'd814,32'd836,32'd858,32'd880,32'd902,32'd924,32'd946,32'd968,32'd990,32'd1012,32'd1034,32'd1056,32'd1078,32'd1100,32'd1122,32'd1144,32'd1166,32'd1188,32'd1210,32'd1232,32'd1254,32'd1276,32'd1298,32'd1320,32'd1342,32'd1364,32'd1386,32'd1408,32'd1430,32'd1452,32'd1474,32'd1496,32'd1518,32'd1540,32'd1562,32'd1584,32'd1606,32'd1628,32'd1650,32'd1672,32'd1694,32'd1716,32'd1738,32'd1760,32'd1782,32'd1804,32'd1826,32'd1848,32'd1870,32'd1892,32'd1914,32'd1936,32'd1958,32'd1980,32'd2002,32'd2024,32'd2046,32'd2068,32'd2090,32'd2112,32'd2134,32'd2156,32'd2178,32'd2200,32'd2222,32'd2244,32'd2266,32'd2288,32'd2310,32'd2332,32'd2354,32'd2376,32'd2398,32'd2420,32'd2442,32'd2464,32'd2486,32'd2508,32'd2530,32'd2552,32'd2574,32'd2596,32'd2618,32'd2640,32'd2662,32'd2684,32'd2706,32'd2728,32'd2750,32'd2772,32'd2794,32'd2816,32'd2838,32'd2860,32'd2882,32'd2904,32'd2926,32'd2948,32'd2970,32'd2992,32'd3014,32'd3036,32'd3058,32'd3080,32'd3102,32'd3124,32'd3146,32'd3168,32'd3190,32'd3212,32'd3234,32'd3256,32'd3278,32'd3300,32'd3322,32'd3344,32'd3366,32'd3388,32'd3410,32'd3432,32'd3454,32'd3476,32'd3498,32'd3520,32'd3542,32'd3564,32'd3586,32'd3608,32'd3630,32'd3652,32'd3674,32'd3696,32'd3718,32'd3740,32'd3762,32'd3784,32'd3806,32'd3828,32'd3850,32'd3872,32'd3894,32'd3916,32'd3938,32'd3960,32'd3982,32'd4004,32'd4026,32'd4048,32'd4070,32'd4092,32'd4114,32'd4136,32'd4158,32'd4180,32'd4202,32'd4224,32'd4246,32'd4268,32'd4290,32'd4312,32'd4334,32'd4356,32'd4378,32'd4400,32'd4422,32'd4444,32'd4466,32'd4488,32'd4510,32'd4532,32'd4554,32'd4576,32'd4598,32'd4620,32'd4642,32'd4664,32'd4686,32'd4708,32'd4730,32'd4752,32'd4774,32'd4796,32'd4818,32'd4840,32'd4862,32'd4884,32'd4906,32'd4928,32'd4950,32'd4972,32'd4994,32'd5016,32'd5038,32'd5060,32'd5082,32'd5104,32'd5126,32'd5148,32'd5170,32'd5192,32'd5214,32'd5236,32'd5258,32'd5280,32'd5302,32'd5324,32'd5346,32'd5368,32'd5390,32'd5412,32'd5434,32'd5456,32'd5478,32'd5500,32'd5522,32'd5544,32'd5566,32'd5588,32'd5610,32'd5632,32'd5654,32'd5676,32'd5698,32'd5720,32'd5742,32'd5764,32'd5786,32'd5808,32'd5830,32'd5852,32'd5874,32'd5896,32'd5918,32'd5940,32'd5962,32'd5984,32'd6006,32'd6028,32'd6050,32'd6072,32'd6094,32'd6116,32'd6138,32'd6160,32'd6182,32'd6204,32'd6226,32'd6248,32'd6270,32'd6292,32'd6314,32'd6336,32'd6358,32'd6380,32'd6402,32'd6424,32'd6446,32'd6468,32'd6490,32'd6512,32'd6534,32'd6556,32'd6578,32'd6600,32'd6622,32'd6644,32'd6666,32'd6688,32'd6710,32'd6732,32'd6754,32'd6776,32'd6798,32'd6820,32'd6842,32'd6864,32'd6886,32'd6908,32'd6930,32'd6952,32'd6974,32'd6996,32'd7018,32'd7040,32'd7062,32'd7084,32'd7106,32'd7128,32'd7150,32'd7172,32'd7194,32'd7216,32'd7238,32'd7260,32'd7282,32'd7304,32'd7326,32'd7348,32'd7370,32'd7392,32'd7414,32'd7436,32'd7458,32'd7480,32'd7502,32'd7524,32'd7546,32'd7568,32'd7590,32'd7612,32'd7634,32'd7656,32'd7678,32'd7700,32'd7722,32'd7744,32'd7766,32'd7788,32'd7810,32'd7832,32'd7854,32'd7876,32'd7898,32'd7920,32'd7942,32'd7964,32'd7986,32'd8008,32'd8030,32'd8052,32'd8074,32'd8096,32'd8118,32'd8140,32'd8162,32'd8184,32'd8206,32'd8228,32'd8250,32'd8272,32'd8294,32'd8316,32'd8338,32'd8360,32'd8382,32'd8404,32'd8426,32'd8448,32'd8470,32'd8492,32'd8514,32'd8536,32'd8558,32'd8580,32'd8602,32'd8624,32'd8646,32'd8668,32'd8690,32'd8712,32'd8734,32'd8756,32'd8778 };matrix[23]='{32'd0,32'd23,32'd46,32'd69,32'd92,32'd115,32'd138,32'd161,32'd184,32'd207,32'd230,32'd253,32'd276,32'd299,32'd322,32'd345,32'd368,32'd391,32'd414,32'd437,32'd460,32'd483,32'd506,32'd529,32'd552,32'd575,32'd598,32'd621,32'd644,32'd667,32'd690,32'd713,32'd736,32'd759,32'd782,32'd805,32'd828,32'd851,32'd874,32'd897,32'd920,32'd943,32'd966,32'd989,32'd1012,32'd1035,32'd1058,32'd1081,32'd1104,32'd1127,32'd1150,32'd1173,32'd1196,32'd1219,32'd1242,32'd1265,32'd1288,32'd1311,32'd1334,32'd1357,32'd1380,32'd1403,32'd1426,32'd1449,32'd1472,32'd1495,32'd1518,32'd1541,32'd1564,32'd1587,32'd1610,32'd1633,32'd1656,32'd1679,32'd1702,32'd1725,32'd1748,32'd1771,32'd1794,32'd1817,32'd1840,32'd1863,32'd1886,32'd1909,32'd1932,32'd1955,32'd1978,32'd2001,32'd2024,32'd2047,32'd2070,32'd2093,32'd2116,32'd2139,32'd2162,32'd2185,32'd2208,32'd2231,32'd2254,32'd2277,32'd2300,32'd2323,32'd2346,32'd2369,32'd2392,32'd2415,32'd2438,32'd2461,32'd2484,32'd2507,32'd2530,32'd2553,32'd2576,32'd2599,32'd2622,32'd2645,32'd2668,32'd2691,32'd2714,32'd2737,32'd2760,32'd2783,32'd2806,32'd2829,32'd2852,32'd2875,32'd2898,32'd2921,32'd2944,32'd2967,32'd2990,32'd3013,32'd3036,32'd3059,32'd3082,32'd3105,32'd3128,32'd3151,32'd3174,32'd3197,32'd3220,32'd3243,32'd3266,32'd3289,32'd3312,32'd3335,32'd3358,32'd3381,32'd3404,32'd3427,32'd3450,32'd3473,32'd3496,32'd3519,32'd3542,32'd3565,32'd3588,32'd3611,32'd3634,32'd3657,32'd3680,32'd3703,32'd3726,32'd3749,32'd3772,32'd3795,32'd3818,32'd3841,32'd3864,32'd3887,32'd3910,32'd3933,32'd3956,32'd3979,32'd4002,32'd4025,32'd4048,32'd4071,32'd4094,32'd4117,32'd4140,32'd4163,32'd4186,32'd4209,32'd4232,32'd4255,32'd4278,32'd4301,32'd4324,32'd4347,32'd4370,32'd4393,32'd4416,32'd4439,32'd4462,32'd4485,32'd4508,32'd4531,32'd4554,32'd4577,32'd4600,32'd4623,32'd4646,32'd4669,32'd4692,32'd4715,32'd4738,32'd4761,32'd4784,32'd4807,32'd4830,32'd4853,32'd4876,32'd4899,32'd4922,32'd4945,32'd4968,32'd4991,32'd5014,32'd5037,32'd5060,32'd5083,32'd5106,32'd5129,32'd5152,32'd5175,32'd5198,32'd5221,32'd5244,32'd5267,32'd5290,32'd5313,32'd5336,32'd5359,32'd5382,32'd5405,32'd5428,32'd5451,32'd5474,32'd5497,32'd5520,32'd5543,32'd5566,32'd5589,32'd5612,32'd5635,32'd5658,32'd5681,32'd5704,32'd5727,32'd5750,32'd5773,32'd5796,32'd5819,32'd5842,32'd5865,32'd5888,32'd5911,32'd5934,32'd5957,32'd5980,32'd6003,32'd6026,32'd6049,32'd6072,32'd6095,32'd6118,32'd6141,32'd6164,32'd6187,32'd6210,32'd6233,32'd6256,32'd6279,32'd6302,32'd6325,32'd6348,32'd6371,32'd6394,32'd6417,32'd6440,32'd6463,32'd6486,32'd6509,32'd6532,32'd6555,32'd6578,32'd6601,32'd6624,32'd6647,32'd6670,32'd6693,32'd6716,32'd6739,32'd6762,32'd6785,32'd6808,32'd6831,32'd6854,32'd6877,32'd6900,32'd6923,32'd6946,32'd6969,32'd6992,32'd7015,32'd7038,32'd7061,32'd7084,32'd7107,32'd7130,32'd7153,32'd7176,32'd7199,32'd7222,32'd7245,32'd7268,32'd7291,32'd7314,32'd7337,32'd7360,32'd7383,32'd7406,32'd7429,32'd7452,32'd7475,32'd7498,32'd7521,32'd7544,32'd7567,32'd7590,32'd7613,32'd7636,32'd7659,32'd7682,32'd7705,32'd7728,32'd7751,32'd7774,32'd7797,32'd7820,32'd7843,32'd7866,32'd7889,32'd7912,32'd7935,32'd7958,32'd7981,32'd8004,32'd8027,32'd8050,32'd8073,32'd8096,32'd8119,32'd8142,32'd8165,32'd8188,32'd8211,32'd8234,32'd8257,32'd8280,32'd8303,32'd8326,32'd8349,32'd8372,32'd8395,32'd8418,32'd8441,32'd8464,32'd8487,32'd8510,32'd8533,32'd8556,32'd8579,32'd8602,32'd8625,32'd8648,32'd8671,32'd8694,32'd8717,32'd8740,32'd8763,32'd8786,32'd8809,32'd8832,32'd8855,32'd8878,32'd8901,32'd8924,32'd8947,32'd8970,32'd8993,32'd9016,32'd9039,32'd9062,32'd9085,32'd9108,32'd9131,32'd9154,32'd9177 };matrix[24]='{32'd0,32'd24,32'd48,32'd72,32'd96,32'd120,32'd144,32'd168,32'd192,32'd216,32'd240,32'd264,32'd288,32'd312,32'd336,32'd360,32'd384,32'd408,32'd432,32'd456,32'd480,32'd504,32'd528,32'd552,32'd576,32'd600,32'd624,32'd648,32'd672,32'd696,32'd720,32'd744,32'd768,32'd792,32'd816,32'd840,32'd864,32'd888,32'd912,32'd936,32'd960,32'd984,32'd1008,32'd1032,32'd1056,32'd1080,32'd1104,32'd1128,32'd1152,32'd1176,32'd1200,32'd1224,32'd1248,32'd1272,32'd1296,32'd1320,32'd1344,32'd1368,32'd1392,32'd1416,32'd1440,32'd1464,32'd1488,32'd1512,32'd1536,32'd1560,32'd1584,32'd1608,32'd1632,32'd1656,32'd1680,32'd1704,32'd1728,32'd1752,32'd1776,32'd1800,32'd1824,32'd1848,32'd1872,32'd1896,32'd1920,32'd1944,32'd1968,32'd1992,32'd2016,32'd2040,32'd2064,32'd2088,32'd2112,32'd2136,32'd2160,32'd2184,32'd2208,32'd2232,32'd2256,32'd2280,32'd2304,32'd2328,32'd2352,32'd2376,32'd2400,32'd2424,32'd2448,32'd2472,32'd2496,32'd2520,32'd2544,32'd2568,32'd2592,32'd2616,32'd2640,32'd2664,32'd2688,32'd2712,32'd2736,32'd2760,32'd2784,32'd2808,32'd2832,32'd2856,32'd2880,32'd2904,32'd2928,32'd2952,32'd2976,32'd3000,32'd3024,32'd3048,32'd3072,32'd3096,32'd3120,32'd3144,32'd3168,32'd3192,32'd3216,32'd3240,32'd3264,32'd3288,32'd3312,32'd3336,32'd3360,32'd3384,32'd3408,32'd3432,32'd3456,32'd3480,32'd3504,32'd3528,32'd3552,32'd3576,32'd3600,32'd3624,32'd3648,32'd3672,32'd3696,32'd3720,32'd3744,32'd3768,32'd3792,32'd3816,32'd3840,32'd3864,32'd3888,32'd3912,32'd3936,32'd3960,32'd3984,32'd4008,32'd4032,32'd4056,32'd4080,32'd4104,32'd4128,32'd4152,32'd4176,32'd4200,32'd4224,32'd4248,32'd4272,32'd4296,32'd4320,32'd4344,32'd4368,32'd4392,32'd4416,32'd4440,32'd4464,32'd4488,32'd4512,32'd4536,32'd4560,32'd4584,32'd4608,32'd4632,32'd4656,32'd4680,32'd4704,32'd4728,32'd4752,32'd4776,32'd4800,32'd4824,32'd4848,32'd4872,32'd4896,32'd4920,32'd4944,32'd4968,32'd4992,32'd5016,32'd5040,32'd5064,32'd5088,32'd5112,32'd5136,32'd5160,32'd5184,32'd5208,32'd5232,32'd5256,32'd5280,32'd5304,32'd5328,32'd5352,32'd5376,32'd5400,32'd5424,32'd5448,32'd5472,32'd5496,32'd5520,32'd5544,32'd5568,32'd5592,32'd5616,32'd5640,32'd5664,32'd5688,32'd5712,32'd5736,32'd5760,32'd5784,32'd5808,32'd5832,32'd5856,32'd5880,32'd5904,32'd5928,32'd5952,32'd5976,32'd6000,32'd6024,32'd6048,32'd6072,32'd6096,32'd6120,32'd6144,32'd6168,32'd6192,32'd6216,32'd6240,32'd6264,32'd6288,32'd6312,32'd6336,32'd6360,32'd6384,32'd6408,32'd6432,32'd6456,32'd6480,32'd6504,32'd6528,32'd6552,32'd6576,32'd6600,32'd6624,32'd6648,32'd6672,32'd6696,32'd6720,32'd6744,32'd6768,32'd6792,32'd6816,32'd6840,32'd6864,32'd6888,32'd6912,32'd6936,32'd6960,32'd6984,32'd7008,32'd7032,32'd7056,32'd7080,32'd7104,32'd7128,32'd7152,32'd7176,32'd7200,32'd7224,32'd7248,32'd7272,32'd7296,32'd7320,32'd7344,32'd7368,32'd7392,32'd7416,32'd7440,32'd7464,32'd7488,32'd7512,32'd7536,32'd7560,32'd7584,32'd7608,32'd7632,32'd7656,32'd7680,32'd7704,32'd7728,32'd7752,32'd7776,32'd7800,32'd7824,32'd7848,32'd7872,32'd7896,32'd7920,32'd7944,32'd7968,32'd7992,32'd8016,32'd8040,32'd8064,32'd8088,32'd8112,32'd8136,32'd8160,32'd8184,32'd8208,32'd8232,32'd8256,32'd8280,32'd8304,32'd8328,32'd8352,32'd8376,32'd8400,32'd8424,32'd8448,32'd8472,32'd8496,32'd8520,32'd8544,32'd8568,32'd8592,32'd8616,32'd8640,32'd8664,32'd8688,32'd8712,32'd8736,32'd8760,32'd8784,32'd8808,32'd8832,32'd8856,32'd8880,32'd8904,32'd8928,32'd8952,32'd8976,32'd9000,32'd9024,32'd9048,32'd9072,32'd9096,32'd9120,32'd9144,32'd9168,32'd9192,32'd9216,32'd9240,32'd9264,32'd9288,32'd9312,32'd9336,32'd9360,32'd9384,32'd9408,32'd9432,32'd9456,32'd9480,32'd9504,32'd9528,32'd9552,32'd9576 };matrix[25]='{32'd0,32'd25,32'd50,32'd75,32'd100,32'd125,32'd150,32'd175,32'd200,32'd225,32'd250,32'd275,32'd300,32'd325,32'd350,32'd375,32'd400,32'd425,32'd450,32'd475,32'd500,32'd525,32'd550,32'd575,32'd600,32'd625,32'd650,32'd675,32'd700,32'd725,32'd750,32'd775,32'd800,32'd825,32'd850,32'd875,32'd900,32'd925,32'd950,32'd975,32'd1000,32'd1025,32'd1050,32'd1075,32'd1100,32'd1125,32'd1150,32'd1175,32'd1200,32'd1225,32'd1250,32'd1275,32'd1300,32'd1325,32'd1350,32'd1375,32'd1400,32'd1425,32'd1450,32'd1475,32'd1500,32'd1525,32'd1550,32'd1575,32'd1600,32'd1625,32'd1650,32'd1675,32'd1700,32'd1725,32'd1750,32'd1775,32'd1800,32'd1825,32'd1850,32'd1875,32'd1900,32'd1925,32'd1950,32'd1975,32'd2000,32'd2025,32'd2050,32'd2075,32'd2100,32'd2125,32'd2150,32'd2175,32'd2200,32'd2225,32'd2250,32'd2275,32'd2300,32'd2325,32'd2350,32'd2375,32'd2400,32'd2425,32'd2450,32'd2475,32'd2500,32'd2525,32'd2550,32'd2575,32'd2600,32'd2625,32'd2650,32'd2675,32'd2700,32'd2725,32'd2750,32'd2775,32'd2800,32'd2825,32'd2850,32'd2875,32'd2900,32'd2925,32'd2950,32'd2975,32'd3000,32'd3025,32'd3050,32'd3075,32'd3100,32'd3125,32'd3150,32'd3175,32'd3200,32'd3225,32'd3250,32'd3275,32'd3300,32'd3325,32'd3350,32'd3375,32'd3400,32'd3425,32'd3450,32'd3475,32'd3500,32'd3525,32'd3550,32'd3575,32'd3600,32'd3625,32'd3650,32'd3675,32'd3700,32'd3725,32'd3750,32'd3775,32'd3800,32'd3825,32'd3850,32'd3875,32'd3900,32'd3925,32'd3950,32'd3975,32'd4000,32'd4025,32'd4050,32'd4075,32'd4100,32'd4125,32'd4150,32'd4175,32'd4200,32'd4225,32'd4250,32'd4275,32'd4300,32'd4325,32'd4350,32'd4375,32'd4400,32'd4425,32'd4450,32'd4475,32'd4500,32'd4525,32'd4550,32'd4575,32'd4600,32'd4625,32'd4650,32'd4675,32'd4700,32'd4725,32'd4750,32'd4775,32'd4800,32'd4825,32'd4850,32'd4875,32'd4900,32'd4925,32'd4950,32'd4975,32'd5000,32'd5025,32'd5050,32'd5075,32'd5100,32'd5125,32'd5150,32'd5175,32'd5200,32'd5225,32'd5250,32'd5275,32'd5300,32'd5325,32'd5350,32'd5375,32'd5400,32'd5425,32'd5450,32'd5475,32'd5500,32'd5525,32'd5550,32'd5575,32'd5600,32'd5625,32'd5650,32'd5675,32'd5700,32'd5725,32'd5750,32'd5775,32'd5800,32'd5825,32'd5850,32'd5875,32'd5900,32'd5925,32'd5950,32'd5975,32'd6000,32'd6025,32'd6050,32'd6075,32'd6100,32'd6125,32'd6150,32'd6175,32'd6200,32'd6225,32'd6250,32'd6275,32'd6300,32'd6325,32'd6350,32'd6375,32'd6400,32'd6425,32'd6450,32'd6475,32'd6500,32'd6525,32'd6550,32'd6575,32'd6600,32'd6625,32'd6650,32'd6675,32'd6700,32'd6725,32'd6750,32'd6775,32'd6800,32'd6825,32'd6850,32'd6875,32'd6900,32'd6925,32'd6950,32'd6975,32'd7000,32'd7025,32'd7050,32'd7075,32'd7100,32'd7125,32'd7150,32'd7175,32'd7200,32'd7225,32'd7250,32'd7275,32'd7300,32'd7325,32'd7350,32'd7375,32'd7400,32'd7425,32'd7450,32'd7475,32'd7500,32'd7525,32'd7550,32'd7575,32'd7600,32'd7625,32'd7650,32'd7675,32'd7700,32'd7725,32'd7750,32'd7775,32'd7800,32'd7825,32'd7850,32'd7875,32'd7900,32'd7925,32'd7950,32'd7975,32'd8000,32'd8025,32'd8050,32'd8075,32'd8100,32'd8125,32'd8150,32'd8175,32'd8200,32'd8225,32'd8250,32'd8275,32'd8300,32'd8325,32'd8350,32'd8375,32'd8400,32'd8425,32'd8450,32'd8475,32'd8500,32'd8525,32'd8550,32'd8575,32'd8600,32'd8625,32'd8650,32'd8675,32'd8700,32'd8725,32'd8750,32'd8775,32'd8800,32'd8825,32'd8850,32'd8875,32'd8900,32'd8925,32'd8950,32'd8975,32'd9000,32'd9025,32'd9050,32'd9075,32'd9100,32'd9125,32'd9150,32'd9175,32'd9200,32'd9225,32'd9250,32'd9275,32'd9300,32'd9325,32'd9350,32'd9375,32'd9400,32'd9425,32'd9450,32'd9475,32'd9500,32'd9525,32'd9550,32'd9575,32'd9600,32'd9625,32'd9650,32'd9675,32'd9700,32'd9725,32'd9750,32'd9775,32'd9800,32'd9825,32'd9850,32'd9875,32'd9900,32'd9925,32'd9950,32'd9975 };matrix[26]='{32'd0,32'd26,32'd52,32'd78,32'd104,32'd130,32'd156,32'd182,32'd208,32'd234,32'd260,32'd286,32'd312,32'd338,32'd364,32'd390,32'd416,32'd442,32'd468,32'd494,32'd520,32'd546,32'd572,32'd598,32'd624,32'd650,32'd676,32'd702,32'd728,32'd754,32'd780,32'd806,32'd832,32'd858,32'd884,32'd910,32'd936,32'd962,32'd988,32'd1014,32'd1040,32'd1066,32'd1092,32'd1118,32'd1144,32'd1170,32'd1196,32'd1222,32'd1248,32'd1274,32'd1300,32'd1326,32'd1352,32'd1378,32'd1404,32'd1430,32'd1456,32'd1482,32'd1508,32'd1534,32'd1560,32'd1586,32'd1612,32'd1638,32'd1664,32'd1690,32'd1716,32'd1742,32'd1768,32'd1794,32'd1820,32'd1846,32'd1872,32'd1898,32'd1924,32'd1950,32'd1976,32'd2002,32'd2028,32'd2054,32'd2080,32'd2106,32'd2132,32'd2158,32'd2184,32'd2210,32'd2236,32'd2262,32'd2288,32'd2314,32'd2340,32'd2366,32'd2392,32'd2418,32'd2444,32'd2470,32'd2496,32'd2522,32'd2548,32'd2574,32'd2600,32'd2626,32'd2652,32'd2678,32'd2704,32'd2730,32'd2756,32'd2782,32'd2808,32'd2834,32'd2860,32'd2886,32'd2912,32'd2938,32'd2964,32'd2990,32'd3016,32'd3042,32'd3068,32'd3094,32'd3120,32'd3146,32'd3172,32'd3198,32'd3224,32'd3250,32'd3276,32'd3302,32'd3328,32'd3354,32'd3380,32'd3406,32'd3432,32'd3458,32'd3484,32'd3510,32'd3536,32'd3562,32'd3588,32'd3614,32'd3640,32'd3666,32'd3692,32'd3718,32'd3744,32'd3770,32'd3796,32'd3822,32'd3848,32'd3874,32'd3900,32'd3926,32'd3952,32'd3978,32'd4004,32'd4030,32'd4056,32'd4082,32'd4108,32'd4134,32'd4160,32'd4186,32'd4212,32'd4238,32'd4264,32'd4290,32'd4316,32'd4342,32'd4368,32'd4394,32'd4420,32'd4446,32'd4472,32'd4498,32'd4524,32'd4550,32'd4576,32'd4602,32'd4628,32'd4654,32'd4680,32'd4706,32'd4732,32'd4758,32'd4784,32'd4810,32'd4836,32'd4862,32'd4888,32'd4914,32'd4940,32'd4966,32'd4992,32'd5018,32'd5044,32'd5070,32'd5096,32'd5122,32'd5148,32'd5174,32'd5200,32'd5226,32'd5252,32'd5278,32'd5304,32'd5330,32'd5356,32'd5382,32'd5408,32'd5434,32'd5460,32'd5486,32'd5512,32'd5538,32'd5564,32'd5590,32'd5616,32'd5642,32'd5668,32'd5694,32'd5720,32'd5746,32'd5772,32'd5798,32'd5824,32'd5850,32'd5876,32'd5902,32'd5928,32'd5954,32'd5980,32'd6006,32'd6032,32'd6058,32'd6084,32'd6110,32'd6136,32'd6162,32'd6188,32'd6214,32'd6240,32'd6266,32'd6292,32'd6318,32'd6344,32'd6370,32'd6396,32'd6422,32'd6448,32'd6474,32'd6500,32'd6526,32'd6552,32'd6578,32'd6604,32'd6630,32'd6656,32'd6682,32'd6708,32'd6734,32'd6760,32'd6786,32'd6812,32'd6838,32'd6864,32'd6890,32'd6916,32'd6942,32'd6968,32'd6994,32'd7020,32'd7046,32'd7072,32'd7098,32'd7124,32'd7150,32'd7176,32'd7202,32'd7228,32'd7254,32'd7280,32'd7306,32'd7332,32'd7358,32'd7384,32'd7410,32'd7436,32'd7462,32'd7488,32'd7514,32'd7540,32'd7566,32'd7592,32'd7618,32'd7644,32'd7670,32'd7696,32'd7722,32'd7748,32'd7774,32'd7800,32'd7826,32'd7852,32'd7878,32'd7904,32'd7930,32'd7956,32'd7982,32'd8008,32'd8034,32'd8060,32'd8086,32'd8112,32'd8138,32'd8164,32'd8190,32'd8216,32'd8242,32'd8268,32'd8294,32'd8320,32'd8346,32'd8372,32'd8398,32'd8424,32'd8450,32'd8476,32'd8502,32'd8528,32'd8554,32'd8580,32'd8606,32'd8632,32'd8658,32'd8684,32'd8710,32'd8736,32'd8762,32'd8788,32'd8814,32'd8840,32'd8866,32'd8892,32'd8918,32'd8944,32'd8970,32'd8996,32'd9022,32'd9048,32'd9074,32'd9100,32'd9126,32'd9152,32'd9178,32'd9204,32'd9230,32'd9256,32'd9282,32'd9308,32'd9334,32'd9360,32'd9386,32'd9412,32'd9438,32'd9464,32'd9490,32'd9516,32'd9542,32'd9568,32'd9594,32'd9620,32'd9646,32'd9672,32'd9698,32'd9724,32'd9750,32'd9776,32'd9802,32'd9828,32'd9854,32'd9880,32'd9906,32'd9932,32'd9958,32'd9984,32'd10010,32'd10036,32'd10062,32'd10088,32'd10114,32'd10140,32'd10166,32'd10192,32'd10218,32'd10244,32'd10270,32'd10296,32'd10322,32'd10348,32'd10374 };matrix[27]='{32'd0,32'd27,32'd54,32'd81,32'd108,32'd135,32'd162,32'd189,32'd216,32'd243,32'd270,32'd297,32'd324,32'd351,32'd378,32'd405,32'd432,32'd459,32'd486,32'd513,32'd540,32'd567,32'd594,32'd621,32'd648,32'd675,32'd702,32'd729,32'd756,32'd783,32'd810,32'd837,32'd864,32'd891,32'd918,32'd945,32'd972,32'd999,32'd1026,32'd1053,32'd1080,32'd1107,32'd1134,32'd1161,32'd1188,32'd1215,32'd1242,32'd1269,32'd1296,32'd1323,32'd1350,32'd1377,32'd1404,32'd1431,32'd1458,32'd1485,32'd1512,32'd1539,32'd1566,32'd1593,32'd1620,32'd1647,32'd1674,32'd1701,32'd1728,32'd1755,32'd1782,32'd1809,32'd1836,32'd1863,32'd1890,32'd1917,32'd1944,32'd1971,32'd1998,32'd2025,32'd2052,32'd2079,32'd2106,32'd2133,32'd2160,32'd2187,32'd2214,32'd2241,32'd2268,32'd2295,32'd2322,32'd2349,32'd2376,32'd2403,32'd2430,32'd2457,32'd2484,32'd2511,32'd2538,32'd2565,32'd2592,32'd2619,32'd2646,32'd2673,32'd2700,32'd2727,32'd2754,32'd2781,32'd2808,32'd2835,32'd2862,32'd2889,32'd2916,32'd2943,32'd2970,32'd2997,32'd3024,32'd3051,32'd3078,32'd3105,32'd3132,32'd3159,32'd3186,32'd3213,32'd3240,32'd3267,32'd3294,32'd3321,32'd3348,32'd3375,32'd3402,32'd3429,32'd3456,32'd3483,32'd3510,32'd3537,32'd3564,32'd3591,32'd3618,32'd3645,32'd3672,32'd3699,32'd3726,32'd3753,32'd3780,32'd3807,32'd3834,32'd3861,32'd3888,32'd3915,32'd3942,32'd3969,32'd3996,32'd4023,32'd4050,32'd4077,32'd4104,32'd4131,32'd4158,32'd4185,32'd4212,32'd4239,32'd4266,32'd4293,32'd4320,32'd4347,32'd4374,32'd4401,32'd4428,32'd4455,32'd4482,32'd4509,32'd4536,32'd4563,32'd4590,32'd4617,32'd4644,32'd4671,32'd4698,32'd4725,32'd4752,32'd4779,32'd4806,32'd4833,32'd4860,32'd4887,32'd4914,32'd4941,32'd4968,32'd4995,32'd5022,32'd5049,32'd5076,32'd5103,32'd5130,32'd5157,32'd5184,32'd5211,32'd5238,32'd5265,32'd5292,32'd5319,32'd5346,32'd5373,32'd5400,32'd5427,32'd5454,32'd5481,32'd5508,32'd5535,32'd5562,32'd5589,32'd5616,32'd5643,32'd5670,32'd5697,32'd5724,32'd5751,32'd5778,32'd5805,32'd5832,32'd5859,32'd5886,32'd5913,32'd5940,32'd5967,32'd5994,32'd6021,32'd6048,32'd6075,32'd6102,32'd6129,32'd6156,32'd6183,32'd6210,32'd6237,32'd6264,32'd6291,32'd6318,32'd6345,32'd6372,32'd6399,32'd6426,32'd6453,32'd6480,32'd6507,32'd6534,32'd6561,32'd6588,32'd6615,32'd6642,32'd6669,32'd6696,32'd6723,32'd6750,32'd6777,32'd6804,32'd6831,32'd6858,32'd6885,32'd6912,32'd6939,32'd6966,32'd6993,32'd7020,32'd7047,32'd7074,32'd7101,32'd7128,32'd7155,32'd7182,32'd7209,32'd7236,32'd7263,32'd7290,32'd7317,32'd7344,32'd7371,32'd7398,32'd7425,32'd7452,32'd7479,32'd7506,32'd7533,32'd7560,32'd7587,32'd7614,32'd7641,32'd7668,32'd7695,32'd7722,32'd7749,32'd7776,32'd7803,32'd7830,32'd7857,32'd7884,32'd7911,32'd7938,32'd7965,32'd7992,32'd8019,32'd8046,32'd8073,32'd8100,32'd8127,32'd8154,32'd8181,32'd8208,32'd8235,32'd8262,32'd8289,32'd8316,32'd8343,32'd8370,32'd8397,32'd8424,32'd8451,32'd8478,32'd8505,32'd8532,32'd8559,32'd8586,32'd8613,32'd8640,32'd8667,32'd8694,32'd8721,32'd8748,32'd8775,32'd8802,32'd8829,32'd8856,32'd8883,32'd8910,32'd8937,32'd8964,32'd8991,32'd9018,32'd9045,32'd9072,32'd9099,32'd9126,32'd9153,32'd9180,32'd9207,32'd9234,32'd9261,32'd9288,32'd9315,32'd9342,32'd9369,32'd9396,32'd9423,32'd9450,32'd9477,32'd9504,32'd9531,32'd9558,32'd9585,32'd9612,32'd9639,32'd9666,32'd9693,32'd9720,32'd9747,32'd9774,32'd9801,32'd9828,32'd9855,32'd9882,32'd9909,32'd9936,32'd9963,32'd9990,32'd10017,32'd10044,32'd10071,32'd10098,32'd10125,32'd10152,32'd10179,32'd10206,32'd10233,32'd10260,32'd10287,32'd10314,32'd10341,32'd10368,32'd10395,32'd10422,32'd10449,32'd10476,32'd10503,32'd10530,32'd10557,32'd10584,32'd10611,32'd10638,32'd10665,32'd10692,32'd10719,32'd10746,32'd10773 };matrix[28]='{32'd0,32'd28,32'd56,32'd84,32'd112,32'd140,32'd168,32'd196,32'd224,32'd252,32'd280,32'd308,32'd336,32'd364,32'd392,32'd420,32'd448,32'd476,32'd504,32'd532,32'd560,32'd588,32'd616,32'd644,32'd672,32'd700,32'd728,32'd756,32'd784,32'd812,32'd840,32'd868,32'd896,32'd924,32'd952,32'd980,32'd1008,32'd1036,32'd1064,32'd1092,32'd1120,32'd1148,32'd1176,32'd1204,32'd1232,32'd1260,32'd1288,32'd1316,32'd1344,32'd1372,32'd1400,32'd1428,32'd1456,32'd1484,32'd1512,32'd1540,32'd1568,32'd1596,32'd1624,32'd1652,32'd1680,32'd1708,32'd1736,32'd1764,32'd1792,32'd1820,32'd1848,32'd1876,32'd1904,32'd1932,32'd1960,32'd1988,32'd2016,32'd2044,32'd2072,32'd2100,32'd2128,32'd2156,32'd2184,32'd2212,32'd2240,32'd2268,32'd2296,32'd2324,32'd2352,32'd2380,32'd2408,32'd2436,32'd2464,32'd2492,32'd2520,32'd2548,32'd2576,32'd2604,32'd2632,32'd2660,32'd2688,32'd2716,32'd2744,32'd2772,32'd2800,32'd2828,32'd2856,32'd2884,32'd2912,32'd2940,32'd2968,32'd2996,32'd3024,32'd3052,32'd3080,32'd3108,32'd3136,32'd3164,32'd3192,32'd3220,32'd3248,32'd3276,32'd3304,32'd3332,32'd3360,32'd3388,32'd3416,32'd3444,32'd3472,32'd3500,32'd3528,32'd3556,32'd3584,32'd3612,32'd3640,32'd3668,32'd3696,32'd3724,32'd3752,32'd3780,32'd3808,32'd3836,32'd3864,32'd3892,32'd3920,32'd3948,32'd3976,32'd4004,32'd4032,32'd4060,32'd4088,32'd4116,32'd4144,32'd4172,32'd4200,32'd4228,32'd4256,32'd4284,32'd4312,32'd4340,32'd4368,32'd4396,32'd4424,32'd4452,32'd4480,32'd4508,32'd4536,32'd4564,32'd4592,32'd4620,32'd4648,32'd4676,32'd4704,32'd4732,32'd4760,32'd4788,32'd4816,32'd4844,32'd4872,32'd4900,32'd4928,32'd4956,32'd4984,32'd5012,32'd5040,32'd5068,32'd5096,32'd5124,32'd5152,32'd5180,32'd5208,32'd5236,32'd5264,32'd5292,32'd5320,32'd5348,32'd5376,32'd5404,32'd5432,32'd5460,32'd5488,32'd5516,32'd5544,32'd5572,32'd5600,32'd5628,32'd5656,32'd5684,32'd5712,32'd5740,32'd5768,32'd5796,32'd5824,32'd5852,32'd5880,32'd5908,32'd5936,32'd5964,32'd5992,32'd6020,32'd6048,32'd6076,32'd6104,32'd6132,32'd6160,32'd6188,32'd6216,32'd6244,32'd6272,32'd6300,32'd6328,32'd6356,32'd6384,32'd6412,32'd6440,32'd6468,32'd6496,32'd6524,32'd6552,32'd6580,32'd6608,32'd6636,32'd6664,32'd6692,32'd6720,32'd6748,32'd6776,32'd6804,32'd6832,32'd6860,32'd6888,32'd6916,32'd6944,32'd6972,32'd7000,32'd7028,32'd7056,32'd7084,32'd7112,32'd7140,32'd7168,32'd7196,32'd7224,32'd7252,32'd7280,32'd7308,32'd7336,32'd7364,32'd7392,32'd7420,32'd7448,32'd7476,32'd7504,32'd7532,32'd7560,32'd7588,32'd7616,32'd7644,32'd7672,32'd7700,32'd7728,32'd7756,32'd7784,32'd7812,32'd7840,32'd7868,32'd7896,32'd7924,32'd7952,32'd7980,32'd8008,32'd8036,32'd8064,32'd8092,32'd8120,32'd8148,32'd8176,32'd8204,32'd8232,32'd8260,32'd8288,32'd8316,32'd8344,32'd8372,32'd8400,32'd8428,32'd8456,32'd8484,32'd8512,32'd8540,32'd8568,32'd8596,32'd8624,32'd8652,32'd8680,32'd8708,32'd8736,32'd8764,32'd8792,32'd8820,32'd8848,32'd8876,32'd8904,32'd8932,32'd8960,32'd8988,32'd9016,32'd9044,32'd9072,32'd9100,32'd9128,32'd9156,32'd9184,32'd9212,32'd9240,32'd9268,32'd9296,32'd9324,32'd9352,32'd9380,32'd9408,32'd9436,32'd9464,32'd9492,32'd9520,32'd9548,32'd9576,32'd9604,32'd9632,32'd9660,32'd9688,32'd9716,32'd9744,32'd9772,32'd9800,32'd9828,32'd9856,32'd9884,32'd9912,32'd9940,32'd9968,32'd9996,32'd10024,32'd10052,32'd10080,32'd10108,32'd10136,32'd10164,32'd10192,32'd10220,32'd10248,32'd10276,32'd10304,32'd10332,32'd10360,32'd10388,32'd10416,32'd10444,32'd10472,32'd10500,32'd10528,32'd10556,32'd10584,32'd10612,32'd10640,32'd10668,32'd10696,32'd10724,32'd10752,32'd10780,32'd10808,32'd10836,32'd10864,32'd10892,32'd10920,32'd10948,32'd10976,32'd11004,32'd11032,32'd11060,32'd11088,32'd11116,32'd11144,32'd11172 };matrix[29]='{32'd0,32'd29,32'd58,32'd87,32'd116,32'd145,32'd174,32'd203,32'd232,32'd261,32'd290,32'd319,32'd348,32'd377,32'd406,32'd435,32'd464,32'd493,32'd522,32'd551,32'd580,32'd609,32'd638,32'd667,32'd696,32'd725,32'd754,32'd783,32'd812,32'd841,32'd870,32'd899,32'd928,32'd957,32'd986,32'd1015,32'd1044,32'd1073,32'd1102,32'd1131,32'd1160,32'd1189,32'd1218,32'd1247,32'd1276,32'd1305,32'd1334,32'd1363,32'd1392,32'd1421,32'd1450,32'd1479,32'd1508,32'd1537,32'd1566,32'd1595,32'd1624,32'd1653,32'd1682,32'd1711,32'd1740,32'd1769,32'd1798,32'd1827,32'd1856,32'd1885,32'd1914,32'd1943,32'd1972,32'd2001,32'd2030,32'd2059,32'd2088,32'd2117,32'd2146,32'd2175,32'd2204,32'd2233,32'd2262,32'd2291,32'd2320,32'd2349,32'd2378,32'd2407,32'd2436,32'd2465,32'd2494,32'd2523,32'd2552,32'd2581,32'd2610,32'd2639,32'd2668,32'd2697,32'd2726,32'd2755,32'd2784,32'd2813,32'd2842,32'd2871,32'd2900,32'd2929,32'd2958,32'd2987,32'd3016,32'd3045,32'd3074,32'd3103,32'd3132,32'd3161,32'd3190,32'd3219,32'd3248,32'd3277,32'd3306,32'd3335,32'd3364,32'd3393,32'd3422,32'd3451,32'd3480,32'd3509,32'd3538,32'd3567,32'd3596,32'd3625,32'd3654,32'd3683,32'd3712,32'd3741,32'd3770,32'd3799,32'd3828,32'd3857,32'd3886,32'd3915,32'd3944,32'd3973,32'd4002,32'd4031,32'd4060,32'd4089,32'd4118,32'd4147,32'd4176,32'd4205,32'd4234,32'd4263,32'd4292,32'd4321,32'd4350,32'd4379,32'd4408,32'd4437,32'd4466,32'd4495,32'd4524,32'd4553,32'd4582,32'd4611,32'd4640,32'd4669,32'd4698,32'd4727,32'd4756,32'd4785,32'd4814,32'd4843,32'd4872,32'd4901,32'd4930,32'd4959,32'd4988,32'd5017,32'd5046,32'd5075,32'd5104,32'd5133,32'd5162,32'd5191,32'd5220,32'd5249,32'd5278,32'd5307,32'd5336,32'd5365,32'd5394,32'd5423,32'd5452,32'd5481,32'd5510,32'd5539,32'd5568,32'd5597,32'd5626,32'd5655,32'd5684,32'd5713,32'd5742,32'd5771,32'd5800,32'd5829,32'd5858,32'd5887,32'd5916,32'd5945,32'd5974,32'd6003,32'd6032,32'd6061,32'd6090,32'd6119,32'd6148,32'd6177,32'd6206,32'd6235,32'd6264,32'd6293,32'd6322,32'd6351,32'd6380,32'd6409,32'd6438,32'd6467,32'd6496,32'd6525,32'd6554,32'd6583,32'd6612,32'd6641,32'd6670,32'd6699,32'd6728,32'd6757,32'd6786,32'd6815,32'd6844,32'd6873,32'd6902,32'd6931,32'd6960,32'd6989,32'd7018,32'd7047,32'd7076,32'd7105,32'd7134,32'd7163,32'd7192,32'd7221,32'd7250,32'd7279,32'd7308,32'd7337,32'd7366,32'd7395,32'd7424,32'd7453,32'd7482,32'd7511,32'd7540,32'd7569,32'd7598,32'd7627,32'd7656,32'd7685,32'd7714,32'd7743,32'd7772,32'd7801,32'd7830,32'd7859,32'd7888,32'd7917,32'd7946,32'd7975,32'd8004,32'd8033,32'd8062,32'd8091,32'd8120,32'd8149,32'd8178,32'd8207,32'd8236,32'd8265,32'd8294,32'd8323,32'd8352,32'd8381,32'd8410,32'd8439,32'd8468,32'd8497,32'd8526,32'd8555,32'd8584,32'd8613,32'd8642,32'd8671,32'd8700,32'd8729,32'd8758,32'd8787,32'd8816,32'd8845,32'd8874,32'd8903,32'd8932,32'd8961,32'd8990,32'd9019,32'd9048,32'd9077,32'd9106,32'd9135,32'd9164,32'd9193,32'd9222,32'd9251,32'd9280,32'd9309,32'd9338,32'd9367,32'd9396,32'd9425,32'd9454,32'd9483,32'd9512,32'd9541,32'd9570,32'd9599,32'd9628,32'd9657,32'd9686,32'd9715,32'd9744,32'd9773,32'd9802,32'd9831,32'd9860,32'd9889,32'd9918,32'd9947,32'd9976,32'd10005,32'd10034,32'd10063,32'd10092,32'd10121,32'd10150,32'd10179,32'd10208,32'd10237,32'd10266,32'd10295,32'd10324,32'd10353,32'd10382,32'd10411,32'd10440,32'd10469,32'd10498,32'd10527,32'd10556,32'd10585,32'd10614,32'd10643,32'd10672,32'd10701,32'd10730,32'd10759,32'd10788,32'd10817,32'd10846,32'd10875,32'd10904,32'd10933,32'd10962,32'd10991,32'd11020,32'd11049,32'd11078,32'd11107,32'd11136,32'd11165,32'd11194,32'd11223,32'd11252,32'd11281,32'd11310,32'd11339,32'd11368,32'd11397,32'd11426,32'd11455,32'd11484,32'd11513,32'd11542,32'd11571 };matrix[30]='{32'd0,32'd30,32'd60,32'd90,32'd120,32'd150,32'd180,32'd210,32'd240,32'd270,32'd300,32'd330,32'd360,32'd390,32'd420,32'd450,32'd480,32'd510,32'd540,32'd570,32'd600,32'd630,32'd660,32'd690,32'd720,32'd750,32'd780,32'd810,32'd840,32'd870,32'd900,32'd930,32'd960,32'd990,32'd1020,32'd1050,32'd1080,32'd1110,32'd1140,32'd1170,32'd1200,32'd1230,32'd1260,32'd1290,32'd1320,32'd1350,32'd1380,32'd1410,32'd1440,32'd1470,32'd1500,32'd1530,32'd1560,32'd1590,32'd1620,32'd1650,32'd1680,32'd1710,32'd1740,32'd1770,32'd1800,32'd1830,32'd1860,32'd1890,32'd1920,32'd1950,32'd1980,32'd2010,32'd2040,32'd2070,32'd2100,32'd2130,32'd2160,32'd2190,32'd2220,32'd2250,32'd2280,32'd2310,32'd2340,32'd2370,32'd2400,32'd2430,32'd2460,32'd2490,32'd2520,32'd2550,32'd2580,32'd2610,32'd2640,32'd2670,32'd2700,32'd2730,32'd2760,32'd2790,32'd2820,32'd2850,32'd2880,32'd2910,32'd2940,32'd2970,32'd3000,32'd3030,32'd3060,32'd3090,32'd3120,32'd3150,32'd3180,32'd3210,32'd3240,32'd3270,32'd3300,32'd3330,32'd3360,32'd3390,32'd3420,32'd3450,32'd3480,32'd3510,32'd3540,32'd3570,32'd3600,32'd3630,32'd3660,32'd3690,32'd3720,32'd3750,32'd3780,32'd3810,32'd3840,32'd3870,32'd3900,32'd3930,32'd3960,32'd3990,32'd4020,32'd4050,32'd4080,32'd4110,32'd4140,32'd4170,32'd4200,32'd4230,32'd4260,32'd4290,32'd4320,32'd4350,32'd4380,32'd4410,32'd4440,32'd4470,32'd4500,32'd4530,32'd4560,32'd4590,32'd4620,32'd4650,32'd4680,32'd4710,32'd4740,32'd4770,32'd4800,32'd4830,32'd4860,32'd4890,32'd4920,32'd4950,32'd4980,32'd5010,32'd5040,32'd5070,32'd5100,32'd5130,32'd5160,32'd5190,32'd5220,32'd5250,32'd5280,32'd5310,32'd5340,32'd5370,32'd5400,32'd5430,32'd5460,32'd5490,32'd5520,32'd5550,32'd5580,32'd5610,32'd5640,32'd5670,32'd5700,32'd5730,32'd5760,32'd5790,32'd5820,32'd5850,32'd5880,32'd5910,32'd5940,32'd5970,32'd6000,32'd6030,32'd6060,32'd6090,32'd6120,32'd6150,32'd6180,32'd6210,32'd6240,32'd6270,32'd6300,32'd6330,32'd6360,32'd6390,32'd6420,32'd6450,32'd6480,32'd6510,32'd6540,32'd6570,32'd6600,32'd6630,32'd6660,32'd6690,32'd6720,32'd6750,32'd6780,32'd6810,32'd6840,32'd6870,32'd6900,32'd6930,32'd6960,32'd6990,32'd7020,32'd7050,32'd7080,32'd7110,32'd7140,32'd7170,32'd7200,32'd7230,32'd7260,32'd7290,32'd7320,32'd7350,32'd7380,32'd7410,32'd7440,32'd7470,32'd7500,32'd7530,32'd7560,32'd7590,32'd7620,32'd7650,32'd7680,32'd7710,32'd7740,32'd7770,32'd7800,32'd7830,32'd7860,32'd7890,32'd7920,32'd7950,32'd7980,32'd8010,32'd8040,32'd8070,32'd8100,32'd8130,32'd8160,32'd8190,32'd8220,32'd8250,32'd8280,32'd8310,32'd8340,32'd8370,32'd8400,32'd8430,32'd8460,32'd8490,32'd8520,32'd8550,32'd8580,32'd8610,32'd8640,32'd8670,32'd8700,32'd8730,32'd8760,32'd8790,32'd8820,32'd8850,32'd8880,32'd8910,32'd8940,32'd8970,32'd9000,32'd9030,32'd9060,32'd9090,32'd9120,32'd9150,32'd9180,32'd9210,32'd9240,32'd9270,32'd9300,32'd9330,32'd9360,32'd9390,32'd9420,32'd9450,32'd9480,32'd9510,32'd9540,32'd9570,32'd9600,32'd9630,32'd9660,32'd9690,32'd9720,32'd9750,32'd9780,32'd9810,32'd9840,32'd9870,32'd9900,32'd9930,32'd9960,32'd9990,32'd10020,32'd10050,32'd10080,32'd10110,32'd10140,32'd10170,32'd10200,32'd10230,32'd10260,32'd10290,32'd10320,32'd10350,32'd10380,32'd10410,32'd10440,32'd10470,32'd10500,32'd10530,32'd10560,32'd10590,32'd10620,32'd10650,32'd10680,32'd10710,32'd10740,32'd10770,32'd10800,32'd10830,32'd10860,32'd10890,32'd10920,32'd10950,32'd10980,32'd11010,32'd11040,32'd11070,32'd11100,32'd11130,32'd11160,32'd11190,32'd11220,32'd11250,32'd11280,32'd11310,32'd11340,32'd11370,32'd11400,32'd11430,32'd11460,32'd11490,32'd11520,32'd11550,32'd11580,32'd11610,32'd11640,32'd11670,32'd11700,32'd11730,32'd11760,32'd11790,32'd11820,32'd11850,32'd11880,32'd11910,32'd11940,32'd11970 };matrix[31]='{32'd0,32'd31,32'd62,32'd93,32'd124,32'd155,32'd186,32'd217,32'd248,32'd279,32'd310,32'd341,32'd372,32'd403,32'd434,32'd465,32'd496,32'd527,32'd558,32'd589,32'd620,32'd651,32'd682,32'd713,32'd744,32'd775,32'd806,32'd837,32'd868,32'd899,32'd930,32'd961,32'd992,32'd1023,32'd1054,32'd1085,32'd1116,32'd1147,32'd1178,32'd1209,32'd1240,32'd1271,32'd1302,32'd1333,32'd1364,32'd1395,32'd1426,32'd1457,32'd1488,32'd1519,32'd1550,32'd1581,32'd1612,32'd1643,32'd1674,32'd1705,32'd1736,32'd1767,32'd1798,32'd1829,32'd1860,32'd1891,32'd1922,32'd1953,32'd1984,32'd2015,32'd2046,32'd2077,32'd2108,32'd2139,32'd2170,32'd2201,32'd2232,32'd2263,32'd2294,32'd2325,32'd2356,32'd2387,32'd2418,32'd2449,32'd2480,32'd2511,32'd2542,32'd2573,32'd2604,32'd2635,32'd2666,32'd2697,32'd2728,32'd2759,32'd2790,32'd2821,32'd2852,32'd2883,32'd2914,32'd2945,32'd2976,32'd3007,32'd3038,32'd3069,32'd3100,32'd3131,32'd3162,32'd3193,32'd3224,32'd3255,32'd3286,32'd3317,32'd3348,32'd3379,32'd3410,32'd3441,32'd3472,32'd3503,32'd3534,32'd3565,32'd3596,32'd3627,32'd3658,32'd3689,32'd3720,32'd3751,32'd3782,32'd3813,32'd3844,32'd3875,32'd3906,32'd3937,32'd3968,32'd3999,32'd4030,32'd4061,32'd4092,32'd4123,32'd4154,32'd4185,32'd4216,32'd4247,32'd4278,32'd4309,32'd4340,32'd4371,32'd4402,32'd4433,32'd4464,32'd4495,32'd4526,32'd4557,32'd4588,32'd4619,32'd4650,32'd4681,32'd4712,32'd4743,32'd4774,32'd4805,32'd4836,32'd4867,32'd4898,32'd4929,32'd4960,32'd4991,32'd5022,32'd5053,32'd5084,32'd5115,32'd5146,32'd5177,32'd5208,32'd5239,32'd5270,32'd5301,32'd5332,32'd5363,32'd5394,32'd5425,32'd5456,32'd5487,32'd5518,32'd5549,32'd5580,32'd5611,32'd5642,32'd5673,32'd5704,32'd5735,32'd5766,32'd5797,32'd5828,32'd5859,32'd5890,32'd5921,32'd5952,32'd5983,32'd6014,32'd6045,32'd6076,32'd6107,32'd6138,32'd6169,32'd6200,32'd6231,32'd6262,32'd6293,32'd6324,32'd6355,32'd6386,32'd6417,32'd6448,32'd6479,32'd6510,32'd6541,32'd6572,32'd6603,32'd6634,32'd6665,32'd6696,32'd6727,32'd6758,32'd6789,32'd6820,32'd6851,32'd6882,32'd6913,32'd6944,32'd6975,32'd7006,32'd7037,32'd7068,32'd7099,32'd7130,32'd7161,32'd7192,32'd7223,32'd7254,32'd7285,32'd7316,32'd7347,32'd7378,32'd7409,32'd7440,32'd7471,32'd7502,32'd7533,32'd7564,32'd7595,32'd7626,32'd7657,32'd7688,32'd7719,32'd7750,32'd7781,32'd7812,32'd7843,32'd7874,32'd7905,32'd7936,32'd7967,32'd7998,32'd8029,32'd8060,32'd8091,32'd8122,32'd8153,32'd8184,32'd8215,32'd8246,32'd8277,32'd8308,32'd8339,32'd8370,32'd8401,32'd8432,32'd8463,32'd8494,32'd8525,32'd8556,32'd8587,32'd8618,32'd8649,32'd8680,32'd8711,32'd8742,32'd8773,32'd8804,32'd8835,32'd8866,32'd8897,32'd8928,32'd8959,32'd8990,32'd9021,32'd9052,32'd9083,32'd9114,32'd9145,32'd9176,32'd9207,32'd9238,32'd9269,32'd9300,32'd9331,32'd9362,32'd9393,32'd9424,32'd9455,32'd9486,32'd9517,32'd9548,32'd9579,32'd9610,32'd9641,32'd9672,32'd9703,32'd9734,32'd9765,32'd9796,32'd9827,32'd9858,32'd9889,32'd9920,32'd9951,32'd9982,32'd10013,32'd10044,32'd10075,32'd10106,32'd10137,32'd10168,32'd10199,32'd10230,32'd10261,32'd10292,32'd10323,32'd10354,32'd10385,32'd10416,32'd10447,32'd10478,32'd10509,32'd10540,32'd10571,32'd10602,32'd10633,32'd10664,32'd10695,32'd10726,32'd10757,32'd10788,32'd10819,32'd10850,32'd10881,32'd10912,32'd10943,32'd10974,32'd11005,32'd11036,32'd11067,32'd11098,32'd11129,32'd11160,32'd11191,32'd11222,32'd11253,32'd11284,32'd11315,32'd11346,32'd11377,32'd11408,32'd11439,32'd11470,32'd11501,32'd11532,32'd11563,32'd11594,32'd11625,32'd11656,32'd11687,32'd11718,32'd11749,32'd11780,32'd11811,32'd11842,32'd11873,32'd11904,32'd11935,32'd11966,32'd11997,32'd12028,32'd12059,32'd12090,32'd12121,32'd12152,32'd12183,32'd12214,32'd12245,32'd12276,32'd12307,32'd12338,32'd12369 };matrix[32]='{32'd0,32'd32,32'd64,32'd96,32'd128,32'd160,32'd192,32'd224,32'd256,32'd288,32'd320,32'd352,32'd384,32'd416,32'd448,32'd480,32'd512,32'd544,32'd576,32'd608,32'd640,32'd672,32'd704,32'd736,32'd768,32'd800,32'd832,32'd864,32'd896,32'd928,32'd960,32'd992,32'd1024,32'd1056,32'd1088,32'd1120,32'd1152,32'd1184,32'd1216,32'd1248,32'd1280,32'd1312,32'd1344,32'd1376,32'd1408,32'd1440,32'd1472,32'd1504,32'd1536,32'd1568,32'd1600,32'd1632,32'd1664,32'd1696,32'd1728,32'd1760,32'd1792,32'd1824,32'd1856,32'd1888,32'd1920,32'd1952,32'd1984,32'd2016,32'd2048,32'd2080,32'd2112,32'd2144,32'd2176,32'd2208,32'd2240,32'd2272,32'd2304,32'd2336,32'd2368,32'd2400,32'd2432,32'd2464,32'd2496,32'd2528,32'd2560,32'd2592,32'd2624,32'd2656,32'd2688,32'd2720,32'd2752,32'd2784,32'd2816,32'd2848,32'd2880,32'd2912,32'd2944,32'd2976,32'd3008,32'd3040,32'd3072,32'd3104,32'd3136,32'd3168,32'd3200,32'd3232,32'd3264,32'd3296,32'd3328,32'd3360,32'd3392,32'd3424,32'd3456,32'd3488,32'd3520,32'd3552,32'd3584,32'd3616,32'd3648,32'd3680,32'd3712,32'd3744,32'd3776,32'd3808,32'd3840,32'd3872,32'd3904,32'd3936,32'd3968,32'd4000,32'd4032,32'd4064,32'd4096,32'd4128,32'd4160,32'd4192,32'd4224,32'd4256,32'd4288,32'd4320,32'd4352,32'd4384,32'd4416,32'd4448,32'd4480,32'd4512,32'd4544,32'd4576,32'd4608,32'd4640,32'd4672,32'd4704,32'd4736,32'd4768,32'd4800,32'd4832,32'd4864,32'd4896,32'd4928,32'd4960,32'd4992,32'd5024,32'd5056,32'd5088,32'd5120,32'd5152,32'd5184,32'd5216,32'd5248,32'd5280,32'd5312,32'd5344,32'd5376,32'd5408,32'd5440,32'd5472,32'd5504,32'd5536,32'd5568,32'd5600,32'd5632,32'd5664,32'd5696,32'd5728,32'd5760,32'd5792,32'd5824,32'd5856,32'd5888,32'd5920,32'd5952,32'd5984,32'd6016,32'd6048,32'd6080,32'd6112,32'd6144,32'd6176,32'd6208,32'd6240,32'd6272,32'd6304,32'd6336,32'd6368,32'd6400,32'd6432,32'd6464,32'd6496,32'd6528,32'd6560,32'd6592,32'd6624,32'd6656,32'd6688,32'd6720,32'd6752,32'd6784,32'd6816,32'd6848,32'd6880,32'd6912,32'd6944,32'd6976,32'd7008,32'd7040,32'd7072,32'd7104,32'd7136,32'd7168,32'd7200,32'd7232,32'd7264,32'd7296,32'd7328,32'd7360,32'd7392,32'd7424,32'd7456,32'd7488,32'd7520,32'd7552,32'd7584,32'd7616,32'd7648,32'd7680,32'd7712,32'd7744,32'd7776,32'd7808,32'd7840,32'd7872,32'd7904,32'd7936,32'd7968,32'd8000,32'd8032,32'd8064,32'd8096,32'd8128,32'd8160,32'd8192,32'd8224,32'd8256,32'd8288,32'd8320,32'd8352,32'd8384,32'd8416,32'd8448,32'd8480,32'd8512,32'd8544,32'd8576,32'd8608,32'd8640,32'd8672,32'd8704,32'd8736,32'd8768,32'd8800,32'd8832,32'd8864,32'd8896,32'd8928,32'd8960,32'd8992,32'd9024,32'd9056,32'd9088,32'd9120,32'd9152,32'd9184,32'd9216,32'd9248,32'd9280,32'd9312,32'd9344,32'd9376,32'd9408,32'd9440,32'd9472,32'd9504,32'd9536,32'd9568,32'd9600,32'd9632,32'd9664,32'd9696,32'd9728,32'd9760,32'd9792,32'd9824,32'd9856,32'd9888,32'd9920,32'd9952,32'd9984,32'd10016,32'd10048,32'd10080,32'd10112,32'd10144,32'd10176,32'd10208,32'd10240,32'd10272,32'd10304,32'd10336,32'd10368,32'd10400,32'd10432,32'd10464,32'd10496,32'd10528,32'd10560,32'd10592,32'd10624,32'd10656,32'd10688,32'd10720,32'd10752,32'd10784,32'd10816,32'd10848,32'd10880,32'd10912,32'd10944,32'd10976,32'd11008,32'd11040,32'd11072,32'd11104,32'd11136,32'd11168,32'd11200,32'd11232,32'd11264,32'd11296,32'd11328,32'd11360,32'd11392,32'd11424,32'd11456,32'd11488,32'd11520,32'd11552,32'd11584,32'd11616,32'd11648,32'd11680,32'd11712,32'd11744,32'd11776,32'd11808,32'd11840,32'd11872,32'd11904,32'd11936,32'd11968,32'd12000,32'd12032,32'd12064,32'd12096,32'd12128,32'd12160,32'd12192,32'd12224,32'd12256,32'd12288,32'd12320,32'd12352,32'd12384,32'd12416,32'd12448,32'd12480,32'd12512,32'd12544,32'd12576,32'd12608,32'd12640,32'd12672,32'd12704,32'd12736,32'd12768 };matrix[33]='{32'd0,32'd33,32'd66,32'd99,32'd132,32'd165,32'd198,32'd231,32'd264,32'd297,32'd330,32'd363,32'd396,32'd429,32'd462,32'd495,32'd528,32'd561,32'd594,32'd627,32'd660,32'd693,32'd726,32'd759,32'd792,32'd825,32'd858,32'd891,32'd924,32'd957,32'd990,32'd1023,32'd1056,32'd1089,32'd1122,32'd1155,32'd1188,32'd1221,32'd1254,32'd1287,32'd1320,32'd1353,32'd1386,32'd1419,32'd1452,32'd1485,32'd1518,32'd1551,32'd1584,32'd1617,32'd1650,32'd1683,32'd1716,32'd1749,32'd1782,32'd1815,32'd1848,32'd1881,32'd1914,32'd1947,32'd1980,32'd2013,32'd2046,32'd2079,32'd2112,32'd2145,32'd2178,32'd2211,32'd2244,32'd2277,32'd2310,32'd2343,32'd2376,32'd2409,32'd2442,32'd2475,32'd2508,32'd2541,32'd2574,32'd2607,32'd2640,32'd2673,32'd2706,32'd2739,32'd2772,32'd2805,32'd2838,32'd2871,32'd2904,32'd2937,32'd2970,32'd3003,32'd3036,32'd3069,32'd3102,32'd3135,32'd3168,32'd3201,32'd3234,32'd3267,32'd3300,32'd3333,32'd3366,32'd3399,32'd3432,32'd3465,32'd3498,32'd3531,32'd3564,32'd3597,32'd3630,32'd3663,32'd3696,32'd3729,32'd3762,32'd3795,32'd3828,32'd3861,32'd3894,32'd3927,32'd3960,32'd3993,32'd4026,32'd4059,32'd4092,32'd4125,32'd4158,32'd4191,32'd4224,32'd4257,32'd4290,32'd4323,32'd4356,32'd4389,32'd4422,32'd4455,32'd4488,32'd4521,32'd4554,32'd4587,32'd4620,32'd4653,32'd4686,32'd4719,32'd4752,32'd4785,32'd4818,32'd4851,32'd4884,32'd4917,32'd4950,32'd4983,32'd5016,32'd5049,32'd5082,32'd5115,32'd5148,32'd5181,32'd5214,32'd5247,32'd5280,32'd5313,32'd5346,32'd5379,32'd5412,32'd5445,32'd5478,32'd5511,32'd5544,32'd5577,32'd5610,32'd5643,32'd5676,32'd5709,32'd5742,32'd5775,32'd5808,32'd5841,32'd5874,32'd5907,32'd5940,32'd5973,32'd6006,32'd6039,32'd6072,32'd6105,32'd6138,32'd6171,32'd6204,32'd6237,32'd6270,32'd6303,32'd6336,32'd6369,32'd6402,32'd6435,32'd6468,32'd6501,32'd6534,32'd6567,32'd6600,32'd6633,32'd6666,32'd6699,32'd6732,32'd6765,32'd6798,32'd6831,32'd6864,32'd6897,32'd6930,32'd6963,32'd6996,32'd7029,32'd7062,32'd7095,32'd7128,32'd7161,32'd7194,32'd7227,32'd7260,32'd7293,32'd7326,32'd7359,32'd7392,32'd7425,32'd7458,32'd7491,32'd7524,32'd7557,32'd7590,32'd7623,32'd7656,32'd7689,32'd7722,32'd7755,32'd7788,32'd7821,32'd7854,32'd7887,32'd7920,32'd7953,32'd7986,32'd8019,32'd8052,32'd8085,32'd8118,32'd8151,32'd8184,32'd8217,32'd8250,32'd8283,32'd8316,32'd8349,32'd8382,32'd8415,32'd8448,32'd8481,32'd8514,32'd8547,32'd8580,32'd8613,32'd8646,32'd8679,32'd8712,32'd8745,32'd8778,32'd8811,32'd8844,32'd8877,32'd8910,32'd8943,32'd8976,32'd9009,32'd9042,32'd9075,32'd9108,32'd9141,32'd9174,32'd9207,32'd9240,32'd9273,32'd9306,32'd9339,32'd9372,32'd9405,32'd9438,32'd9471,32'd9504,32'd9537,32'd9570,32'd9603,32'd9636,32'd9669,32'd9702,32'd9735,32'd9768,32'd9801,32'd9834,32'd9867,32'd9900,32'd9933,32'd9966,32'd9999,32'd10032,32'd10065,32'd10098,32'd10131,32'd10164,32'd10197,32'd10230,32'd10263,32'd10296,32'd10329,32'd10362,32'd10395,32'd10428,32'd10461,32'd10494,32'd10527,32'd10560,32'd10593,32'd10626,32'd10659,32'd10692,32'd10725,32'd10758,32'd10791,32'd10824,32'd10857,32'd10890,32'd10923,32'd10956,32'd10989,32'd11022,32'd11055,32'd11088,32'd11121,32'd11154,32'd11187,32'd11220,32'd11253,32'd11286,32'd11319,32'd11352,32'd11385,32'd11418,32'd11451,32'd11484,32'd11517,32'd11550,32'd11583,32'd11616,32'd11649,32'd11682,32'd11715,32'd11748,32'd11781,32'd11814,32'd11847,32'd11880,32'd11913,32'd11946,32'd11979,32'd12012,32'd12045,32'd12078,32'd12111,32'd12144,32'd12177,32'd12210,32'd12243,32'd12276,32'd12309,32'd12342,32'd12375,32'd12408,32'd12441,32'd12474,32'd12507,32'd12540,32'd12573,32'd12606,32'd12639,32'd12672,32'd12705,32'd12738,32'd12771,32'd12804,32'd12837,32'd12870,32'd12903,32'd12936,32'd12969,32'd13002,32'd13035,32'd13068,32'd13101,32'd13134,32'd13167 };matrix[34]='{32'd0,32'd34,32'd68,32'd102,32'd136,32'd170,32'd204,32'd238,32'd272,32'd306,32'd340,32'd374,32'd408,32'd442,32'd476,32'd510,32'd544,32'd578,32'd612,32'd646,32'd680,32'd714,32'd748,32'd782,32'd816,32'd850,32'd884,32'd918,32'd952,32'd986,32'd1020,32'd1054,32'd1088,32'd1122,32'd1156,32'd1190,32'd1224,32'd1258,32'd1292,32'd1326,32'd1360,32'd1394,32'd1428,32'd1462,32'd1496,32'd1530,32'd1564,32'd1598,32'd1632,32'd1666,32'd1700,32'd1734,32'd1768,32'd1802,32'd1836,32'd1870,32'd1904,32'd1938,32'd1972,32'd2006,32'd2040,32'd2074,32'd2108,32'd2142,32'd2176,32'd2210,32'd2244,32'd2278,32'd2312,32'd2346,32'd2380,32'd2414,32'd2448,32'd2482,32'd2516,32'd2550,32'd2584,32'd2618,32'd2652,32'd2686,32'd2720,32'd2754,32'd2788,32'd2822,32'd2856,32'd2890,32'd2924,32'd2958,32'd2992,32'd3026,32'd3060,32'd3094,32'd3128,32'd3162,32'd3196,32'd3230,32'd3264,32'd3298,32'd3332,32'd3366,32'd3400,32'd3434,32'd3468,32'd3502,32'd3536,32'd3570,32'd3604,32'd3638,32'd3672,32'd3706,32'd3740,32'd3774,32'd3808,32'd3842,32'd3876,32'd3910,32'd3944,32'd3978,32'd4012,32'd4046,32'd4080,32'd4114,32'd4148,32'd4182,32'd4216,32'd4250,32'd4284,32'd4318,32'd4352,32'd4386,32'd4420,32'd4454,32'd4488,32'd4522,32'd4556,32'd4590,32'd4624,32'd4658,32'd4692,32'd4726,32'd4760,32'd4794,32'd4828,32'd4862,32'd4896,32'd4930,32'd4964,32'd4998,32'd5032,32'd5066,32'd5100,32'd5134,32'd5168,32'd5202,32'd5236,32'd5270,32'd5304,32'd5338,32'd5372,32'd5406,32'd5440,32'd5474,32'd5508,32'd5542,32'd5576,32'd5610,32'd5644,32'd5678,32'd5712,32'd5746,32'd5780,32'd5814,32'd5848,32'd5882,32'd5916,32'd5950,32'd5984,32'd6018,32'd6052,32'd6086,32'd6120,32'd6154,32'd6188,32'd6222,32'd6256,32'd6290,32'd6324,32'd6358,32'd6392,32'd6426,32'd6460,32'd6494,32'd6528,32'd6562,32'd6596,32'd6630,32'd6664,32'd6698,32'd6732,32'd6766,32'd6800,32'd6834,32'd6868,32'd6902,32'd6936,32'd6970,32'd7004,32'd7038,32'd7072,32'd7106,32'd7140,32'd7174,32'd7208,32'd7242,32'd7276,32'd7310,32'd7344,32'd7378,32'd7412,32'd7446,32'd7480,32'd7514,32'd7548,32'd7582,32'd7616,32'd7650,32'd7684,32'd7718,32'd7752,32'd7786,32'd7820,32'd7854,32'd7888,32'd7922,32'd7956,32'd7990,32'd8024,32'd8058,32'd8092,32'd8126,32'd8160,32'd8194,32'd8228,32'd8262,32'd8296,32'd8330,32'd8364,32'd8398,32'd8432,32'd8466,32'd8500,32'd8534,32'd8568,32'd8602,32'd8636,32'd8670,32'd8704,32'd8738,32'd8772,32'd8806,32'd8840,32'd8874,32'd8908,32'd8942,32'd8976,32'd9010,32'd9044,32'd9078,32'd9112,32'd9146,32'd9180,32'd9214,32'd9248,32'd9282,32'd9316,32'd9350,32'd9384,32'd9418,32'd9452,32'd9486,32'd9520,32'd9554,32'd9588,32'd9622,32'd9656,32'd9690,32'd9724,32'd9758,32'd9792,32'd9826,32'd9860,32'd9894,32'd9928,32'd9962,32'd9996,32'd10030,32'd10064,32'd10098,32'd10132,32'd10166,32'd10200,32'd10234,32'd10268,32'd10302,32'd10336,32'd10370,32'd10404,32'd10438,32'd10472,32'd10506,32'd10540,32'd10574,32'd10608,32'd10642,32'd10676,32'd10710,32'd10744,32'd10778,32'd10812,32'd10846,32'd10880,32'd10914,32'd10948,32'd10982,32'd11016,32'd11050,32'd11084,32'd11118,32'd11152,32'd11186,32'd11220,32'd11254,32'd11288,32'd11322,32'd11356,32'd11390,32'd11424,32'd11458,32'd11492,32'd11526,32'd11560,32'd11594,32'd11628,32'd11662,32'd11696,32'd11730,32'd11764,32'd11798,32'd11832,32'd11866,32'd11900,32'd11934,32'd11968,32'd12002,32'd12036,32'd12070,32'd12104,32'd12138,32'd12172,32'd12206,32'd12240,32'd12274,32'd12308,32'd12342,32'd12376,32'd12410,32'd12444,32'd12478,32'd12512,32'd12546,32'd12580,32'd12614,32'd12648,32'd12682,32'd12716,32'd12750,32'd12784,32'd12818,32'd12852,32'd12886,32'd12920,32'd12954,32'd12988,32'd13022,32'd13056,32'd13090,32'd13124,32'd13158,32'd13192,32'd13226,32'd13260,32'd13294,32'd13328,32'd13362,32'd13396,32'd13430,32'd13464,32'd13498,32'd13532,32'd13566 };matrix[35]='{32'd0,32'd35,32'd70,32'd105,32'd140,32'd175,32'd210,32'd245,32'd280,32'd315,32'd350,32'd385,32'd420,32'd455,32'd490,32'd525,32'd560,32'd595,32'd630,32'd665,32'd700,32'd735,32'd770,32'd805,32'd840,32'd875,32'd910,32'd945,32'd980,32'd1015,32'd1050,32'd1085,32'd1120,32'd1155,32'd1190,32'd1225,32'd1260,32'd1295,32'd1330,32'd1365,32'd1400,32'd1435,32'd1470,32'd1505,32'd1540,32'd1575,32'd1610,32'd1645,32'd1680,32'd1715,32'd1750,32'd1785,32'd1820,32'd1855,32'd1890,32'd1925,32'd1960,32'd1995,32'd2030,32'd2065,32'd2100,32'd2135,32'd2170,32'd2205,32'd2240,32'd2275,32'd2310,32'd2345,32'd2380,32'd2415,32'd2450,32'd2485,32'd2520,32'd2555,32'd2590,32'd2625,32'd2660,32'd2695,32'd2730,32'd2765,32'd2800,32'd2835,32'd2870,32'd2905,32'd2940,32'd2975,32'd3010,32'd3045,32'd3080,32'd3115,32'd3150,32'd3185,32'd3220,32'd3255,32'd3290,32'd3325,32'd3360,32'd3395,32'd3430,32'd3465,32'd3500,32'd3535,32'd3570,32'd3605,32'd3640,32'd3675,32'd3710,32'd3745,32'd3780,32'd3815,32'd3850,32'd3885,32'd3920,32'd3955,32'd3990,32'd4025,32'd4060,32'd4095,32'd4130,32'd4165,32'd4200,32'd4235,32'd4270,32'd4305,32'd4340,32'd4375,32'd4410,32'd4445,32'd4480,32'd4515,32'd4550,32'd4585,32'd4620,32'd4655,32'd4690,32'd4725,32'd4760,32'd4795,32'd4830,32'd4865,32'd4900,32'd4935,32'd4970,32'd5005,32'd5040,32'd5075,32'd5110,32'd5145,32'd5180,32'd5215,32'd5250,32'd5285,32'd5320,32'd5355,32'd5390,32'd5425,32'd5460,32'd5495,32'd5530,32'd5565,32'd5600,32'd5635,32'd5670,32'd5705,32'd5740,32'd5775,32'd5810,32'd5845,32'd5880,32'd5915,32'd5950,32'd5985,32'd6020,32'd6055,32'd6090,32'd6125,32'd6160,32'd6195,32'd6230,32'd6265,32'd6300,32'd6335,32'd6370,32'd6405,32'd6440,32'd6475,32'd6510,32'd6545,32'd6580,32'd6615,32'd6650,32'd6685,32'd6720,32'd6755,32'd6790,32'd6825,32'd6860,32'd6895,32'd6930,32'd6965,32'd7000,32'd7035,32'd7070,32'd7105,32'd7140,32'd7175,32'd7210,32'd7245,32'd7280,32'd7315,32'd7350,32'd7385,32'd7420,32'd7455,32'd7490,32'd7525,32'd7560,32'd7595,32'd7630,32'd7665,32'd7700,32'd7735,32'd7770,32'd7805,32'd7840,32'd7875,32'd7910,32'd7945,32'd7980,32'd8015,32'd8050,32'd8085,32'd8120,32'd8155,32'd8190,32'd8225,32'd8260,32'd8295,32'd8330,32'd8365,32'd8400,32'd8435,32'd8470,32'd8505,32'd8540,32'd8575,32'd8610,32'd8645,32'd8680,32'd8715,32'd8750,32'd8785,32'd8820,32'd8855,32'd8890,32'd8925,32'd8960,32'd8995,32'd9030,32'd9065,32'd9100,32'd9135,32'd9170,32'd9205,32'd9240,32'd9275,32'd9310,32'd9345,32'd9380,32'd9415,32'd9450,32'd9485,32'd9520,32'd9555,32'd9590,32'd9625,32'd9660,32'd9695,32'd9730,32'd9765,32'd9800,32'd9835,32'd9870,32'd9905,32'd9940,32'd9975,32'd10010,32'd10045,32'd10080,32'd10115,32'd10150,32'd10185,32'd10220,32'd10255,32'd10290,32'd10325,32'd10360,32'd10395,32'd10430,32'd10465,32'd10500,32'd10535,32'd10570,32'd10605,32'd10640,32'd10675,32'd10710,32'd10745,32'd10780,32'd10815,32'd10850,32'd10885,32'd10920,32'd10955,32'd10990,32'd11025,32'd11060,32'd11095,32'd11130,32'd11165,32'd11200,32'd11235,32'd11270,32'd11305,32'd11340,32'd11375,32'd11410,32'd11445,32'd11480,32'd11515,32'd11550,32'd11585,32'd11620,32'd11655,32'd11690,32'd11725,32'd11760,32'd11795,32'd11830,32'd11865,32'd11900,32'd11935,32'd11970,32'd12005,32'd12040,32'd12075,32'd12110,32'd12145,32'd12180,32'd12215,32'd12250,32'd12285,32'd12320,32'd12355,32'd12390,32'd12425,32'd12460,32'd12495,32'd12530,32'd12565,32'd12600,32'd12635,32'd12670,32'd12705,32'd12740,32'd12775,32'd12810,32'd12845,32'd12880,32'd12915,32'd12950,32'd12985,32'd13020,32'd13055,32'd13090,32'd13125,32'd13160,32'd13195,32'd13230,32'd13265,32'd13300,32'd13335,32'd13370,32'd13405,32'd13440,32'd13475,32'd13510,32'd13545,32'd13580,32'd13615,32'd13650,32'd13685,32'd13720,32'd13755,32'd13790,32'd13825,32'd13860,32'd13895,32'd13930,32'd13965 };matrix[36]='{32'd0,32'd36,32'd72,32'd108,32'd144,32'd180,32'd216,32'd252,32'd288,32'd324,32'd360,32'd396,32'd432,32'd468,32'd504,32'd540,32'd576,32'd612,32'd648,32'd684,32'd720,32'd756,32'd792,32'd828,32'd864,32'd900,32'd936,32'd972,32'd1008,32'd1044,32'd1080,32'd1116,32'd1152,32'd1188,32'd1224,32'd1260,32'd1296,32'd1332,32'd1368,32'd1404,32'd1440,32'd1476,32'd1512,32'd1548,32'd1584,32'd1620,32'd1656,32'd1692,32'd1728,32'd1764,32'd1800,32'd1836,32'd1872,32'd1908,32'd1944,32'd1980,32'd2016,32'd2052,32'd2088,32'd2124,32'd2160,32'd2196,32'd2232,32'd2268,32'd2304,32'd2340,32'd2376,32'd2412,32'd2448,32'd2484,32'd2520,32'd2556,32'd2592,32'd2628,32'd2664,32'd2700,32'd2736,32'd2772,32'd2808,32'd2844,32'd2880,32'd2916,32'd2952,32'd2988,32'd3024,32'd3060,32'd3096,32'd3132,32'd3168,32'd3204,32'd3240,32'd3276,32'd3312,32'd3348,32'd3384,32'd3420,32'd3456,32'd3492,32'd3528,32'd3564,32'd3600,32'd3636,32'd3672,32'd3708,32'd3744,32'd3780,32'd3816,32'd3852,32'd3888,32'd3924,32'd3960,32'd3996,32'd4032,32'd4068,32'd4104,32'd4140,32'd4176,32'd4212,32'd4248,32'd4284,32'd4320,32'd4356,32'd4392,32'd4428,32'd4464,32'd4500,32'd4536,32'd4572,32'd4608,32'd4644,32'd4680,32'd4716,32'd4752,32'd4788,32'd4824,32'd4860,32'd4896,32'd4932,32'd4968,32'd5004,32'd5040,32'd5076,32'd5112,32'd5148,32'd5184,32'd5220,32'd5256,32'd5292,32'd5328,32'd5364,32'd5400,32'd5436,32'd5472,32'd5508,32'd5544,32'd5580,32'd5616,32'd5652,32'd5688,32'd5724,32'd5760,32'd5796,32'd5832,32'd5868,32'd5904,32'd5940,32'd5976,32'd6012,32'd6048,32'd6084,32'd6120,32'd6156,32'd6192,32'd6228,32'd6264,32'd6300,32'd6336,32'd6372,32'd6408,32'd6444,32'd6480,32'd6516,32'd6552,32'd6588,32'd6624,32'd6660,32'd6696,32'd6732,32'd6768,32'd6804,32'd6840,32'd6876,32'd6912,32'd6948,32'd6984,32'd7020,32'd7056,32'd7092,32'd7128,32'd7164,32'd7200,32'd7236,32'd7272,32'd7308,32'd7344,32'd7380,32'd7416,32'd7452,32'd7488,32'd7524,32'd7560,32'd7596,32'd7632,32'd7668,32'd7704,32'd7740,32'd7776,32'd7812,32'd7848,32'd7884,32'd7920,32'd7956,32'd7992,32'd8028,32'd8064,32'd8100,32'd8136,32'd8172,32'd8208,32'd8244,32'd8280,32'd8316,32'd8352,32'd8388,32'd8424,32'd8460,32'd8496,32'd8532,32'd8568,32'd8604,32'd8640,32'd8676,32'd8712,32'd8748,32'd8784,32'd8820,32'd8856,32'd8892,32'd8928,32'd8964,32'd9000,32'd9036,32'd9072,32'd9108,32'd9144,32'd9180,32'd9216,32'd9252,32'd9288,32'd9324,32'd9360,32'd9396,32'd9432,32'd9468,32'd9504,32'd9540,32'd9576,32'd9612,32'd9648,32'd9684,32'd9720,32'd9756,32'd9792,32'd9828,32'd9864,32'd9900,32'd9936,32'd9972,32'd10008,32'd10044,32'd10080,32'd10116,32'd10152,32'd10188,32'd10224,32'd10260,32'd10296,32'd10332,32'd10368,32'd10404,32'd10440,32'd10476,32'd10512,32'd10548,32'd10584,32'd10620,32'd10656,32'd10692,32'd10728,32'd10764,32'd10800,32'd10836,32'd10872,32'd10908,32'd10944,32'd10980,32'd11016,32'd11052,32'd11088,32'd11124,32'd11160,32'd11196,32'd11232,32'd11268,32'd11304,32'd11340,32'd11376,32'd11412,32'd11448,32'd11484,32'd11520,32'd11556,32'd11592,32'd11628,32'd11664,32'd11700,32'd11736,32'd11772,32'd11808,32'd11844,32'd11880,32'd11916,32'd11952,32'd11988,32'd12024,32'd12060,32'd12096,32'd12132,32'd12168,32'd12204,32'd12240,32'd12276,32'd12312,32'd12348,32'd12384,32'd12420,32'd12456,32'd12492,32'd12528,32'd12564,32'd12600,32'd12636,32'd12672,32'd12708,32'd12744,32'd12780,32'd12816,32'd12852,32'd12888,32'd12924,32'd12960,32'd12996,32'd13032,32'd13068,32'd13104,32'd13140,32'd13176,32'd13212,32'd13248,32'd13284,32'd13320,32'd13356,32'd13392,32'd13428,32'd13464,32'd13500,32'd13536,32'd13572,32'd13608,32'd13644,32'd13680,32'd13716,32'd13752,32'd13788,32'd13824,32'd13860,32'd13896,32'd13932,32'd13968,32'd14004,32'd14040,32'd14076,32'd14112,32'd14148,32'd14184,32'd14220,32'd14256,32'd14292,32'd14328,32'd14364 };matrix[37]='{32'd0,32'd37,32'd74,32'd111,32'd148,32'd185,32'd222,32'd259,32'd296,32'd333,32'd370,32'd407,32'd444,32'd481,32'd518,32'd555,32'd592,32'd629,32'd666,32'd703,32'd740,32'd777,32'd814,32'd851,32'd888,32'd925,32'd962,32'd999,32'd1036,32'd1073,32'd1110,32'd1147,32'd1184,32'd1221,32'd1258,32'd1295,32'd1332,32'd1369,32'd1406,32'd1443,32'd1480,32'd1517,32'd1554,32'd1591,32'd1628,32'd1665,32'd1702,32'd1739,32'd1776,32'd1813,32'd1850,32'd1887,32'd1924,32'd1961,32'd1998,32'd2035,32'd2072,32'd2109,32'd2146,32'd2183,32'd2220,32'd2257,32'd2294,32'd2331,32'd2368,32'd2405,32'd2442,32'd2479,32'd2516,32'd2553,32'd2590,32'd2627,32'd2664,32'd2701,32'd2738,32'd2775,32'd2812,32'd2849,32'd2886,32'd2923,32'd2960,32'd2997,32'd3034,32'd3071,32'd3108,32'd3145,32'd3182,32'd3219,32'd3256,32'd3293,32'd3330,32'd3367,32'd3404,32'd3441,32'd3478,32'd3515,32'd3552,32'd3589,32'd3626,32'd3663,32'd3700,32'd3737,32'd3774,32'd3811,32'd3848,32'd3885,32'd3922,32'd3959,32'd3996,32'd4033,32'd4070,32'd4107,32'd4144,32'd4181,32'd4218,32'd4255,32'd4292,32'd4329,32'd4366,32'd4403,32'd4440,32'd4477,32'd4514,32'd4551,32'd4588,32'd4625,32'd4662,32'd4699,32'd4736,32'd4773,32'd4810,32'd4847,32'd4884,32'd4921,32'd4958,32'd4995,32'd5032,32'd5069,32'd5106,32'd5143,32'd5180,32'd5217,32'd5254,32'd5291,32'd5328,32'd5365,32'd5402,32'd5439,32'd5476,32'd5513,32'd5550,32'd5587,32'd5624,32'd5661,32'd5698,32'd5735,32'd5772,32'd5809,32'd5846,32'd5883,32'd5920,32'd5957,32'd5994,32'd6031,32'd6068,32'd6105,32'd6142,32'd6179,32'd6216,32'd6253,32'd6290,32'd6327,32'd6364,32'd6401,32'd6438,32'd6475,32'd6512,32'd6549,32'd6586,32'd6623,32'd6660,32'd6697,32'd6734,32'd6771,32'd6808,32'd6845,32'd6882,32'd6919,32'd6956,32'd6993,32'd7030,32'd7067,32'd7104,32'd7141,32'd7178,32'd7215,32'd7252,32'd7289,32'd7326,32'd7363,32'd7400,32'd7437,32'd7474,32'd7511,32'd7548,32'd7585,32'd7622,32'd7659,32'd7696,32'd7733,32'd7770,32'd7807,32'd7844,32'd7881,32'd7918,32'd7955,32'd7992,32'd8029,32'd8066,32'd8103,32'd8140,32'd8177,32'd8214,32'd8251,32'd8288,32'd8325,32'd8362,32'd8399,32'd8436,32'd8473,32'd8510,32'd8547,32'd8584,32'd8621,32'd8658,32'd8695,32'd8732,32'd8769,32'd8806,32'd8843,32'd8880,32'd8917,32'd8954,32'd8991,32'd9028,32'd9065,32'd9102,32'd9139,32'd9176,32'd9213,32'd9250,32'd9287,32'd9324,32'd9361,32'd9398,32'd9435,32'd9472,32'd9509,32'd9546,32'd9583,32'd9620,32'd9657,32'd9694,32'd9731,32'd9768,32'd9805,32'd9842,32'd9879,32'd9916,32'd9953,32'd9990,32'd10027,32'd10064,32'd10101,32'd10138,32'd10175,32'd10212,32'd10249,32'd10286,32'd10323,32'd10360,32'd10397,32'd10434,32'd10471,32'd10508,32'd10545,32'd10582,32'd10619,32'd10656,32'd10693,32'd10730,32'd10767,32'd10804,32'd10841,32'd10878,32'd10915,32'd10952,32'd10989,32'd11026,32'd11063,32'd11100,32'd11137,32'd11174,32'd11211,32'd11248,32'd11285,32'd11322,32'd11359,32'd11396,32'd11433,32'd11470,32'd11507,32'd11544,32'd11581,32'd11618,32'd11655,32'd11692,32'd11729,32'd11766,32'd11803,32'd11840,32'd11877,32'd11914,32'd11951,32'd11988,32'd12025,32'd12062,32'd12099,32'd12136,32'd12173,32'd12210,32'd12247,32'd12284,32'd12321,32'd12358,32'd12395,32'd12432,32'd12469,32'd12506,32'd12543,32'd12580,32'd12617,32'd12654,32'd12691,32'd12728,32'd12765,32'd12802,32'd12839,32'd12876,32'd12913,32'd12950,32'd12987,32'd13024,32'd13061,32'd13098,32'd13135,32'd13172,32'd13209,32'd13246,32'd13283,32'd13320,32'd13357,32'd13394,32'd13431,32'd13468,32'd13505,32'd13542,32'd13579,32'd13616,32'd13653,32'd13690,32'd13727,32'd13764,32'd13801,32'd13838,32'd13875,32'd13912,32'd13949,32'd13986,32'd14023,32'd14060,32'd14097,32'd14134,32'd14171,32'd14208,32'd14245,32'd14282,32'd14319,32'd14356,32'd14393,32'd14430,32'd14467,32'd14504,32'd14541,32'd14578,32'd14615,32'd14652,32'd14689,32'd14726,32'd14763 };matrix[38]='{32'd0,32'd38,32'd76,32'd114,32'd152,32'd190,32'd228,32'd266,32'd304,32'd342,32'd380,32'd418,32'd456,32'd494,32'd532,32'd570,32'd608,32'd646,32'd684,32'd722,32'd760,32'd798,32'd836,32'd874,32'd912,32'd950,32'd988,32'd1026,32'd1064,32'd1102,32'd1140,32'd1178,32'd1216,32'd1254,32'd1292,32'd1330,32'd1368,32'd1406,32'd1444,32'd1482,32'd1520,32'd1558,32'd1596,32'd1634,32'd1672,32'd1710,32'd1748,32'd1786,32'd1824,32'd1862,32'd1900,32'd1938,32'd1976,32'd2014,32'd2052,32'd2090,32'd2128,32'd2166,32'd2204,32'd2242,32'd2280,32'd2318,32'd2356,32'd2394,32'd2432,32'd2470,32'd2508,32'd2546,32'd2584,32'd2622,32'd2660,32'd2698,32'd2736,32'd2774,32'd2812,32'd2850,32'd2888,32'd2926,32'd2964,32'd3002,32'd3040,32'd3078,32'd3116,32'd3154,32'd3192,32'd3230,32'd3268,32'd3306,32'd3344,32'd3382,32'd3420,32'd3458,32'd3496,32'd3534,32'd3572,32'd3610,32'd3648,32'd3686,32'd3724,32'd3762,32'd3800,32'd3838,32'd3876,32'd3914,32'd3952,32'd3990,32'd4028,32'd4066,32'd4104,32'd4142,32'd4180,32'd4218,32'd4256,32'd4294,32'd4332,32'd4370,32'd4408,32'd4446,32'd4484,32'd4522,32'd4560,32'd4598,32'd4636,32'd4674,32'd4712,32'd4750,32'd4788,32'd4826,32'd4864,32'd4902,32'd4940,32'd4978,32'd5016,32'd5054,32'd5092,32'd5130,32'd5168,32'd5206,32'd5244,32'd5282,32'd5320,32'd5358,32'd5396,32'd5434,32'd5472,32'd5510,32'd5548,32'd5586,32'd5624,32'd5662,32'd5700,32'd5738,32'd5776,32'd5814,32'd5852,32'd5890,32'd5928,32'd5966,32'd6004,32'd6042,32'd6080,32'd6118,32'd6156,32'd6194,32'd6232,32'd6270,32'd6308,32'd6346,32'd6384,32'd6422,32'd6460,32'd6498,32'd6536,32'd6574,32'd6612,32'd6650,32'd6688,32'd6726,32'd6764,32'd6802,32'd6840,32'd6878,32'd6916,32'd6954,32'd6992,32'd7030,32'd7068,32'd7106,32'd7144,32'd7182,32'd7220,32'd7258,32'd7296,32'd7334,32'd7372,32'd7410,32'd7448,32'd7486,32'd7524,32'd7562,32'd7600,32'd7638,32'd7676,32'd7714,32'd7752,32'd7790,32'd7828,32'd7866,32'd7904,32'd7942,32'd7980,32'd8018,32'd8056,32'd8094,32'd8132,32'd8170,32'd8208,32'd8246,32'd8284,32'd8322,32'd8360,32'd8398,32'd8436,32'd8474,32'd8512,32'd8550,32'd8588,32'd8626,32'd8664,32'd8702,32'd8740,32'd8778,32'd8816,32'd8854,32'd8892,32'd8930,32'd8968,32'd9006,32'd9044,32'd9082,32'd9120,32'd9158,32'd9196,32'd9234,32'd9272,32'd9310,32'd9348,32'd9386,32'd9424,32'd9462,32'd9500,32'd9538,32'd9576,32'd9614,32'd9652,32'd9690,32'd9728,32'd9766,32'd9804,32'd9842,32'd9880,32'd9918,32'd9956,32'd9994,32'd10032,32'd10070,32'd10108,32'd10146,32'd10184,32'd10222,32'd10260,32'd10298,32'd10336,32'd10374,32'd10412,32'd10450,32'd10488,32'd10526,32'd10564,32'd10602,32'd10640,32'd10678,32'd10716,32'd10754,32'd10792,32'd10830,32'd10868,32'd10906,32'd10944,32'd10982,32'd11020,32'd11058,32'd11096,32'd11134,32'd11172,32'd11210,32'd11248,32'd11286,32'd11324,32'd11362,32'd11400,32'd11438,32'd11476,32'd11514,32'd11552,32'd11590,32'd11628,32'd11666,32'd11704,32'd11742,32'd11780,32'd11818,32'd11856,32'd11894,32'd11932,32'd11970,32'd12008,32'd12046,32'd12084,32'd12122,32'd12160,32'd12198,32'd12236,32'd12274,32'd12312,32'd12350,32'd12388,32'd12426,32'd12464,32'd12502,32'd12540,32'd12578,32'd12616,32'd12654,32'd12692,32'd12730,32'd12768,32'd12806,32'd12844,32'd12882,32'd12920,32'd12958,32'd12996,32'd13034,32'd13072,32'd13110,32'd13148,32'd13186,32'd13224,32'd13262,32'd13300,32'd13338,32'd13376,32'd13414,32'd13452,32'd13490,32'd13528,32'd13566,32'd13604,32'd13642,32'd13680,32'd13718,32'd13756,32'd13794,32'd13832,32'd13870,32'd13908,32'd13946,32'd13984,32'd14022,32'd14060,32'd14098,32'd14136,32'd14174,32'd14212,32'd14250,32'd14288,32'd14326,32'd14364,32'd14402,32'd14440,32'd14478,32'd14516,32'd14554,32'd14592,32'd14630,32'd14668,32'd14706,32'd14744,32'd14782,32'd14820,32'd14858,32'd14896,32'd14934,32'd14972,32'd15010,32'd15048,32'd15086,32'd15124,32'd15162 };matrix[39]='{32'd0,32'd39,32'd78,32'd117,32'd156,32'd195,32'd234,32'd273,32'd312,32'd351,32'd390,32'd429,32'd468,32'd507,32'd546,32'd585,32'd624,32'd663,32'd702,32'd741,32'd780,32'd819,32'd858,32'd897,32'd936,32'd975,32'd1014,32'd1053,32'd1092,32'd1131,32'd1170,32'd1209,32'd1248,32'd1287,32'd1326,32'd1365,32'd1404,32'd1443,32'd1482,32'd1521,32'd1560,32'd1599,32'd1638,32'd1677,32'd1716,32'd1755,32'd1794,32'd1833,32'd1872,32'd1911,32'd1950,32'd1989,32'd2028,32'd2067,32'd2106,32'd2145,32'd2184,32'd2223,32'd2262,32'd2301,32'd2340,32'd2379,32'd2418,32'd2457,32'd2496,32'd2535,32'd2574,32'd2613,32'd2652,32'd2691,32'd2730,32'd2769,32'd2808,32'd2847,32'd2886,32'd2925,32'd2964,32'd3003,32'd3042,32'd3081,32'd3120,32'd3159,32'd3198,32'd3237,32'd3276,32'd3315,32'd3354,32'd3393,32'd3432,32'd3471,32'd3510,32'd3549,32'd3588,32'd3627,32'd3666,32'd3705,32'd3744,32'd3783,32'd3822,32'd3861,32'd3900,32'd3939,32'd3978,32'd4017,32'd4056,32'd4095,32'd4134,32'd4173,32'd4212,32'd4251,32'd4290,32'd4329,32'd4368,32'd4407,32'd4446,32'd4485,32'd4524,32'd4563,32'd4602,32'd4641,32'd4680,32'd4719,32'd4758,32'd4797,32'd4836,32'd4875,32'd4914,32'd4953,32'd4992,32'd5031,32'd5070,32'd5109,32'd5148,32'd5187,32'd5226,32'd5265,32'd5304,32'd5343,32'd5382,32'd5421,32'd5460,32'd5499,32'd5538,32'd5577,32'd5616,32'd5655,32'd5694,32'd5733,32'd5772,32'd5811,32'd5850,32'd5889,32'd5928,32'd5967,32'd6006,32'd6045,32'd6084,32'd6123,32'd6162,32'd6201,32'd6240,32'd6279,32'd6318,32'd6357,32'd6396,32'd6435,32'd6474,32'd6513,32'd6552,32'd6591,32'd6630,32'd6669,32'd6708,32'd6747,32'd6786,32'd6825,32'd6864,32'd6903,32'd6942,32'd6981,32'd7020,32'd7059,32'd7098,32'd7137,32'd7176,32'd7215,32'd7254,32'd7293,32'd7332,32'd7371,32'd7410,32'd7449,32'd7488,32'd7527,32'd7566,32'd7605,32'd7644,32'd7683,32'd7722,32'd7761,32'd7800,32'd7839,32'd7878,32'd7917,32'd7956,32'd7995,32'd8034,32'd8073,32'd8112,32'd8151,32'd8190,32'd8229,32'd8268,32'd8307,32'd8346,32'd8385,32'd8424,32'd8463,32'd8502,32'd8541,32'd8580,32'd8619,32'd8658,32'd8697,32'd8736,32'd8775,32'd8814,32'd8853,32'd8892,32'd8931,32'd8970,32'd9009,32'd9048,32'd9087,32'd9126,32'd9165,32'd9204,32'd9243,32'd9282,32'd9321,32'd9360,32'd9399,32'd9438,32'd9477,32'd9516,32'd9555,32'd9594,32'd9633,32'd9672,32'd9711,32'd9750,32'd9789,32'd9828,32'd9867,32'd9906,32'd9945,32'd9984,32'd10023,32'd10062,32'd10101,32'd10140,32'd10179,32'd10218,32'd10257,32'd10296,32'd10335,32'd10374,32'd10413,32'd10452,32'd10491,32'd10530,32'd10569,32'd10608,32'd10647,32'd10686,32'd10725,32'd10764,32'd10803,32'd10842,32'd10881,32'd10920,32'd10959,32'd10998,32'd11037,32'd11076,32'd11115,32'd11154,32'd11193,32'd11232,32'd11271,32'd11310,32'd11349,32'd11388,32'd11427,32'd11466,32'd11505,32'd11544,32'd11583,32'd11622,32'd11661,32'd11700,32'd11739,32'd11778,32'd11817,32'd11856,32'd11895,32'd11934,32'd11973,32'd12012,32'd12051,32'd12090,32'd12129,32'd12168,32'd12207,32'd12246,32'd12285,32'd12324,32'd12363,32'd12402,32'd12441,32'd12480,32'd12519,32'd12558,32'd12597,32'd12636,32'd12675,32'd12714,32'd12753,32'd12792,32'd12831,32'd12870,32'd12909,32'd12948,32'd12987,32'd13026,32'd13065,32'd13104,32'd13143,32'd13182,32'd13221,32'd13260,32'd13299,32'd13338,32'd13377,32'd13416,32'd13455,32'd13494,32'd13533,32'd13572,32'd13611,32'd13650,32'd13689,32'd13728,32'd13767,32'd13806,32'd13845,32'd13884,32'd13923,32'd13962,32'd14001,32'd14040,32'd14079,32'd14118,32'd14157,32'd14196,32'd14235,32'd14274,32'd14313,32'd14352,32'd14391,32'd14430,32'd14469,32'd14508,32'd14547,32'd14586,32'd14625,32'd14664,32'd14703,32'd14742,32'd14781,32'd14820,32'd14859,32'd14898,32'd14937,32'd14976,32'd15015,32'd15054,32'd15093,32'd15132,32'd15171,32'd15210,32'd15249,32'd15288,32'd15327,32'd15366,32'd15405,32'd15444,32'd15483,32'd15522,32'd15561 };matrix[40]='{32'd0,32'd40,32'd80,32'd120,32'd160,32'd200,32'd240,32'd280,32'd320,32'd360,32'd400,32'd440,32'd480,32'd520,32'd560,32'd600,32'd640,32'd680,32'd720,32'd760,32'd800,32'd840,32'd880,32'd920,32'd960,32'd1000,32'd1040,32'd1080,32'd1120,32'd1160,32'd1200,32'd1240,32'd1280,32'd1320,32'd1360,32'd1400,32'd1440,32'd1480,32'd1520,32'd1560,32'd1600,32'd1640,32'd1680,32'd1720,32'd1760,32'd1800,32'd1840,32'd1880,32'd1920,32'd1960,32'd2000,32'd2040,32'd2080,32'd2120,32'd2160,32'd2200,32'd2240,32'd2280,32'd2320,32'd2360,32'd2400,32'd2440,32'd2480,32'd2520,32'd2560,32'd2600,32'd2640,32'd2680,32'd2720,32'd2760,32'd2800,32'd2840,32'd2880,32'd2920,32'd2960,32'd3000,32'd3040,32'd3080,32'd3120,32'd3160,32'd3200,32'd3240,32'd3280,32'd3320,32'd3360,32'd3400,32'd3440,32'd3480,32'd3520,32'd3560,32'd3600,32'd3640,32'd3680,32'd3720,32'd3760,32'd3800,32'd3840,32'd3880,32'd3920,32'd3960,32'd4000,32'd4040,32'd4080,32'd4120,32'd4160,32'd4200,32'd4240,32'd4280,32'd4320,32'd4360,32'd4400,32'd4440,32'd4480,32'd4520,32'd4560,32'd4600,32'd4640,32'd4680,32'd4720,32'd4760,32'd4800,32'd4840,32'd4880,32'd4920,32'd4960,32'd5000,32'd5040,32'd5080,32'd5120,32'd5160,32'd5200,32'd5240,32'd5280,32'd5320,32'd5360,32'd5400,32'd5440,32'd5480,32'd5520,32'd5560,32'd5600,32'd5640,32'd5680,32'd5720,32'd5760,32'd5800,32'd5840,32'd5880,32'd5920,32'd5960,32'd6000,32'd6040,32'd6080,32'd6120,32'd6160,32'd6200,32'd6240,32'd6280,32'd6320,32'd6360,32'd6400,32'd6440,32'd6480,32'd6520,32'd6560,32'd6600,32'd6640,32'd6680,32'd6720,32'd6760,32'd6800,32'd6840,32'd6880,32'd6920,32'd6960,32'd7000,32'd7040,32'd7080,32'd7120,32'd7160,32'd7200,32'd7240,32'd7280,32'd7320,32'd7360,32'd7400,32'd7440,32'd7480,32'd7520,32'd7560,32'd7600,32'd7640,32'd7680,32'd7720,32'd7760,32'd7800,32'd7840,32'd7880,32'd7920,32'd7960,32'd8000,32'd8040,32'd8080,32'd8120,32'd8160,32'd8200,32'd8240,32'd8280,32'd8320,32'd8360,32'd8400,32'd8440,32'd8480,32'd8520,32'd8560,32'd8600,32'd8640,32'd8680,32'd8720,32'd8760,32'd8800,32'd8840,32'd8880,32'd8920,32'd8960,32'd9000,32'd9040,32'd9080,32'd9120,32'd9160,32'd9200,32'd9240,32'd9280,32'd9320,32'd9360,32'd9400,32'd9440,32'd9480,32'd9520,32'd9560,32'd9600,32'd9640,32'd9680,32'd9720,32'd9760,32'd9800,32'd9840,32'd9880,32'd9920,32'd9960,32'd10000,32'd10040,32'd10080,32'd10120,32'd10160,32'd10200,32'd10240,32'd10280,32'd10320,32'd10360,32'd10400,32'd10440,32'd10480,32'd10520,32'd10560,32'd10600,32'd10640,32'd10680,32'd10720,32'd10760,32'd10800,32'd10840,32'd10880,32'd10920,32'd10960,32'd11000,32'd11040,32'd11080,32'd11120,32'd11160,32'd11200,32'd11240,32'd11280,32'd11320,32'd11360,32'd11400,32'd11440,32'd11480,32'd11520,32'd11560,32'd11600,32'd11640,32'd11680,32'd11720,32'd11760,32'd11800,32'd11840,32'd11880,32'd11920,32'd11960,32'd12000,32'd12040,32'd12080,32'd12120,32'd12160,32'd12200,32'd12240,32'd12280,32'd12320,32'd12360,32'd12400,32'd12440,32'd12480,32'd12520,32'd12560,32'd12600,32'd12640,32'd12680,32'd12720,32'd12760,32'd12800,32'd12840,32'd12880,32'd12920,32'd12960,32'd13000,32'd13040,32'd13080,32'd13120,32'd13160,32'd13200,32'd13240,32'd13280,32'd13320,32'd13360,32'd13400,32'd13440,32'd13480,32'd13520,32'd13560,32'd13600,32'd13640,32'd13680,32'd13720,32'd13760,32'd13800,32'd13840,32'd13880,32'd13920,32'd13960,32'd14000,32'd14040,32'd14080,32'd14120,32'd14160,32'd14200,32'd14240,32'd14280,32'd14320,32'd14360,32'd14400,32'd14440,32'd14480,32'd14520,32'd14560,32'd14600,32'd14640,32'd14680,32'd14720,32'd14760,32'd14800,32'd14840,32'd14880,32'd14920,32'd14960,32'd15000,32'd15040,32'd15080,32'd15120,32'd15160,32'd15200,32'd15240,32'd15280,32'd15320,32'd15360,32'd15400,32'd15440,32'd15480,32'd15520,32'd15560,32'd15600,32'd15640,32'd15680,32'd15720,32'd15760,32'd15800,32'd15840,32'd15880,32'd15920,32'd15960 };matrix[41]='{32'd0,32'd41,32'd82,32'd123,32'd164,32'd205,32'd246,32'd287,32'd328,32'd369,32'd410,32'd451,32'd492,32'd533,32'd574,32'd615,32'd656,32'd697,32'd738,32'd779,32'd820,32'd861,32'd902,32'd943,32'd984,32'd1025,32'd1066,32'd1107,32'd1148,32'd1189,32'd1230,32'd1271,32'd1312,32'd1353,32'd1394,32'd1435,32'd1476,32'd1517,32'd1558,32'd1599,32'd1640,32'd1681,32'd1722,32'd1763,32'd1804,32'd1845,32'd1886,32'd1927,32'd1968,32'd2009,32'd2050,32'd2091,32'd2132,32'd2173,32'd2214,32'd2255,32'd2296,32'd2337,32'd2378,32'd2419,32'd2460,32'd2501,32'd2542,32'd2583,32'd2624,32'd2665,32'd2706,32'd2747,32'd2788,32'd2829,32'd2870,32'd2911,32'd2952,32'd2993,32'd3034,32'd3075,32'd3116,32'd3157,32'd3198,32'd3239,32'd3280,32'd3321,32'd3362,32'd3403,32'd3444,32'd3485,32'd3526,32'd3567,32'd3608,32'd3649,32'd3690,32'd3731,32'd3772,32'd3813,32'd3854,32'd3895,32'd3936,32'd3977,32'd4018,32'd4059,32'd4100,32'd4141,32'd4182,32'd4223,32'd4264,32'd4305,32'd4346,32'd4387,32'd4428,32'd4469,32'd4510,32'd4551,32'd4592,32'd4633,32'd4674,32'd4715,32'd4756,32'd4797,32'd4838,32'd4879,32'd4920,32'd4961,32'd5002,32'd5043,32'd5084,32'd5125,32'd5166,32'd5207,32'd5248,32'd5289,32'd5330,32'd5371,32'd5412,32'd5453,32'd5494,32'd5535,32'd5576,32'd5617,32'd5658,32'd5699,32'd5740,32'd5781,32'd5822,32'd5863,32'd5904,32'd5945,32'd5986,32'd6027,32'd6068,32'd6109,32'd6150,32'd6191,32'd6232,32'd6273,32'd6314,32'd6355,32'd6396,32'd6437,32'd6478,32'd6519,32'd6560,32'd6601,32'd6642,32'd6683,32'd6724,32'd6765,32'd6806,32'd6847,32'd6888,32'd6929,32'd6970,32'd7011,32'd7052,32'd7093,32'd7134,32'd7175,32'd7216,32'd7257,32'd7298,32'd7339,32'd7380,32'd7421,32'd7462,32'd7503,32'd7544,32'd7585,32'd7626,32'd7667,32'd7708,32'd7749,32'd7790,32'd7831,32'd7872,32'd7913,32'd7954,32'd7995,32'd8036,32'd8077,32'd8118,32'd8159,32'd8200,32'd8241,32'd8282,32'd8323,32'd8364,32'd8405,32'd8446,32'd8487,32'd8528,32'd8569,32'd8610,32'd8651,32'd8692,32'd8733,32'd8774,32'd8815,32'd8856,32'd8897,32'd8938,32'd8979,32'd9020,32'd9061,32'd9102,32'd9143,32'd9184,32'd9225,32'd9266,32'd9307,32'd9348,32'd9389,32'd9430,32'd9471,32'd9512,32'd9553,32'd9594,32'd9635,32'd9676,32'd9717,32'd9758,32'd9799,32'd9840,32'd9881,32'd9922,32'd9963,32'd10004,32'd10045,32'd10086,32'd10127,32'd10168,32'd10209,32'd10250,32'd10291,32'd10332,32'd10373,32'd10414,32'd10455,32'd10496,32'd10537,32'd10578,32'd10619,32'd10660,32'd10701,32'd10742,32'd10783,32'd10824,32'd10865,32'd10906,32'd10947,32'd10988,32'd11029,32'd11070,32'd11111,32'd11152,32'd11193,32'd11234,32'd11275,32'd11316,32'd11357,32'd11398,32'd11439,32'd11480,32'd11521,32'd11562,32'd11603,32'd11644,32'd11685,32'd11726,32'd11767,32'd11808,32'd11849,32'd11890,32'd11931,32'd11972,32'd12013,32'd12054,32'd12095,32'd12136,32'd12177,32'd12218,32'd12259,32'd12300,32'd12341,32'd12382,32'd12423,32'd12464,32'd12505,32'd12546,32'd12587,32'd12628,32'd12669,32'd12710,32'd12751,32'd12792,32'd12833,32'd12874,32'd12915,32'd12956,32'd12997,32'd13038,32'd13079,32'd13120,32'd13161,32'd13202,32'd13243,32'd13284,32'd13325,32'd13366,32'd13407,32'd13448,32'd13489,32'd13530,32'd13571,32'd13612,32'd13653,32'd13694,32'd13735,32'd13776,32'd13817,32'd13858,32'd13899,32'd13940,32'd13981,32'd14022,32'd14063,32'd14104,32'd14145,32'd14186,32'd14227,32'd14268,32'd14309,32'd14350,32'd14391,32'd14432,32'd14473,32'd14514,32'd14555,32'd14596,32'd14637,32'd14678,32'd14719,32'd14760,32'd14801,32'd14842,32'd14883,32'd14924,32'd14965,32'd15006,32'd15047,32'd15088,32'd15129,32'd15170,32'd15211,32'd15252,32'd15293,32'd15334,32'd15375,32'd15416,32'd15457,32'd15498,32'd15539,32'd15580,32'd15621,32'd15662,32'd15703,32'd15744,32'd15785,32'd15826,32'd15867,32'd15908,32'd15949,32'd15990,32'd16031,32'd16072,32'd16113,32'd16154,32'd16195,32'd16236,32'd16277,32'd16318,32'd16359 };matrix[42]='{32'd0,32'd42,32'd84,32'd126,32'd168,32'd210,32'd252,32'd294,32'd336,32'd378,32'd420,32'd462,32'd504,32'd546,32'd588,32'd630,32'd672,32'd714,32'd756,32'd798,32'd840,32'd882,32'd924,32'd966,32'd1008,32'd1050,32'd1092,32'd1134,32'd1176,32'd1218,32'd1260,32'd1302,32'd1344,32'd1386,32'd1428,32'd1470,32'd1512,32'd1554,32'd1596,32'd1638,32'd1680,32'd1722,32'd1764,32'd1806,32'd1848,32'd1890,32'd1932,32'd1974,32'd2016,32'd2058,32'd2100,32'd2142,32'd2184,32'd2226,32'd2268,32'd2310,32'd2352,32'd2394,32'd2436,32'd2478,32'd2520,32'd2562,32'd2604,32'd2646,32'd2688,32'd2730,32'd2772,32'd2814,32'd2856,32'd2898,32'd2940,32'd2982,32'd3024,32'd3066,32'd3108,32'd3150,32'd3192,32'd3234,32'd3276,32'd3318,32'd3360,32'd3402,32'd3444,32'd3486,32'd3528,32'd3570,32'd3612,32'd3654,32'd3696,32'd3738,32'd3780,32'd3822,32'd3864,32'd3906,32'd3948,32'd3990,32'd4032,32'd4074,32'd4116,32'd4158,32'd4200,32'd4242,32'd4284,32'd4326,32'd4368,32'd4410,32'd4452,32'd4494,32'd4536,32'd4578,32'd4620,32'd4662,32'd4704,32'd4746,32'd4788,32'd4830,32'd4872,32'd4914,32'd4956,32'd4998,32'd5040,32'd5082,32'd5124,32'd5166,32'd5208,32'd5250,32'd5292,32'd5334,32'd5376,32'd5418,32'd5460,32'd5502,32'd5544,32'd5586,32'd5628,32'd5670,32'd5712,32'd5754,32'd5796,32'd5838,32'd5880,32'd5922,32'd5964,32'd6006,32'd6048,32'd6090,32'd6132,32'd6174,32'd6216,32'd6258,32'd6300,32'd6342,32'd6384,32'd6426,32'd6468,32'd6510,32'd6552,32'd6594,32'd6636,32'd6678,32'd6720,32'd6762,32'd6804,32'd6846,32'd6888,32'd6930,32'd6972,32'd7014,32'd7056,32'd7098,32'd7140,32'd7182,32'd7224,32'd7266,32'd7308,32'd7350,32'd7392,32'd7434,32'd7476,32'd7518,32'd7560,32'd7602,32'd7644,32'd7686,32'd7728,32'd7770,32'd7812,32'd7854,32'd7896,32'd7938,32'd7980,32'd8022,32'd8064,32'd8106,32'd8148,32'd8190,32'd8232,32'd8274,32'd8316,32'd8358,32'd8400,32'd8442,32'd8484,32'd8526,32'd8568,32'd8610,32'd8652,32'd8694,32'd8736,32'd8778,32'd8820,32'd8862,32'd8904,32'd8946,32'd8988,32'd9030,32'd9072,32'd9114,32'd9156,32'd9198,32'd9240,32'd9282,32'd9324,32'd9366,32'd9408,32'd9450,32'd9492,32'd9534,32'd9576,32'd9618,32'd9660,32'd9702,32'd9744,32'd9786,32'd9828,32'd9870,32'd9912,32'd9954,32'd9996,32'd10038,32'd10080,32'd10122,32'd10164,32'd10206,32'd10248,32'd10290,32'd10332,32'd10374,32'd10416,32'd10458,32'd10500,32'd10542,32'd10584,32'd10626,32'd10668,32'd10710,32'd10752,32'd10794,32'd10836,32'd10878,32'd10920,32'd10962,32'd11004,32'd11046,32'd11088,32'd11130,32'd11172,32'd11214,32'd11256,32'd11298,32'd11340,32'd11382,32'd11424,32'd11466,32'd11508,32'd11550,32'd11592,32'd11634,32'd11676,32'd11718,32'd11760,32'd11802,32'd11844,32'd11886,32'd11928,32'd11970,32'd12012,32'd12054,32'd12096,32'd12138,32'd12180,32'd12222,32'd12264,32'd12306,32'd12348,32'd12390,32'd12432,32'd12474,32'd12516,32'd12558,32'd12600,32'd12642,32'd12684,32'd12726,32'd12768,32'd12810,32'd12852,32'd12894,32'd12936,32'd12978,32'd13020,32'd13062,32'd13104,32'd13146,32'd13188,32'd13230,32'd13272,32'd13314,32'd13356,32'd13398,32'd13440,32'd13482,32'd13524,32'd13566,32'd13608,32'd13650,32'd13692,32'd13734,32'd13776,32'd13818,32'd13860,32'd13902,32'd13944,32'd13986,32'd14028,32'd14070,32'd14112,32'd14154,32'd14196,32'd14238,32'd14280,32'd14322,32'd14364,32'd14406,32'd14448,32'd14490,32'd14532,32'd14574,32'd14616,32'd14658,32'd14700,32'd14742,32'd14784,32'd14826,32'd14868,32'd14910,32'd14952,32'd14994,32'd15036,32'd15078,32'd15120,32'd15162,32'd15204,32'd15246,32'd15288,32'd15330,32'd15372,32'd15414,32'd15456,32'd15498,32'd15540,32'd15582,32'd15624,32'd15666,32'd15708,32'd15750,32'd15792,32'd15834,32'd15876,32'd15918,32'd15960,32'd16002,32'd16044,32'd16086,32'd16128,32'd16170,32'd16212,32'd16254,32'd16296,32'd16338,32'd16380,32'd16422,32'd16464,32'd16506,32'd16548,32'd16590,32'd16632,32'd16674,32'd16716,32'd16758 };matrix[43]='{32'd0,32'd43,32'd86,32'd129,32'd172,32'd215,32'd258,32'd301,32'd344,32'd387,32'd430,32'd473,32'd516,32'd559,32'd602,32'd645,32'd688,32'd731,32'd774,32'd817,32'd860,32'd903,32'd946,32'd989,32'd1032,32'd1075,32'd1118,32'd1161,32'd1204,32'd1247,32'd1290,32'd1333,32'd1376,32'd1419,32'd1462,32'd1505,32'd1548,32'd1591,32'd1634,32'd1677,32'd1720,32'd1763,32'd1806,32'd1849,32'd1892,32'd1935,32'd1978,32'd2021,32'd2064,32'd2107,32'd2150,32'd2193,32'd2236,32'd2279,32'd2322,32'd2365,32'd2408,32'd2451,32'd2494,32'd2537,32'd2580,32'd2623,32'd2666,32'd2709,32'd2752,32'd2795,32'd2838,32'd2881,32'd2924,32'd2967,32'd3010,32'd3053,32'd3096,32'd3139,32'd3182,32'd3225,32'd3268,32'd3311,32'd3354,32'd3397,32'd3440,32'd3483,32'd3526,32'd3569,32'd3612,32'd3655,32'd3698,32'd3741,32'd3784,32'd3827,32'd3870,32'd3913,32'd3956,32'd3999,32'd4042,32'd4085,32'd4128,32'd4171,32'd4214,32'd4257,32'd4300,32'd4343,32'd4386,32'd4429,32'd4472,32'd4515,32'd4558,32'd4601,32'd4644,32'd4687,32'd4730,32'd4773,32'd4816,32'd4859,32'd4902,32'd4945,32'd4988,32'd5031,32'd5074,32'd5117,32'd5160,32'd5203,32'd5246,32'd5289,32'd5332,32'd5375,32'd5418,32'd5461,32'd5504,32'd5547,32'd5590,32'd5633,32'd5676,32'd5719,32'd5762,32'd5805,32'd5848,32'd5891,32'd5934,32'd5977,32'd6020,32'd6063,32'd6106,32'd6149,32'd6192,32'd6235,32'd6278,32'd6321,32'd6364,32'd6407,32'd6450,32'd6493,32'd6536,32'd6579,32'd6622,32'd6665,32'd6708,32'd6751,32'd6794,32'd6837,32'd6880,32'd6923,32'd6966,32'd7009,32'd7052,32'd7095,32'd7138,32'd7181,32'd7224,32'd7267,32'd7310,32'd7353,32'd7396,32'd7439,32'd7482,32'd7525,32'd7568,32'd7611,32'd7654,32'd7697,32'd7740,32'd7783,32'd7826,32'd7869,32'd7912,32'd7955,32'd7998,32'd8041,32'd8084,32'd8127,32'd8170,32'd8213,32'd8256,32'd8299,32'd8342,32'd8385,32'd8428,32'd8471,32'd8514,32'd8557,32'd8600,32'd8643,32'd8686,32'd8729,32'd8772,32'd8815,32'd8858,32'd8901,32'd8944,32'd8987,32'd9030,32'd9073,32'd9116,32'd9159,32'd9202,32'd9245,32'd9288,32'd9331,32'd9374,32'd9417,32'd9460,32'd9503,32'd9546,32'd9589,32'd9632,32'd9675,32'd9718,32'd9761,32'd9804,32'd9847,32'd9890,32'd9933,32'd9976,32'd10019,32'd10062,32'd10105,32'd10148,32'd10191,32'd10234,32'd10277,32'd10320,32'd10363,32'd10406,32'd10449,32'd10492,32'd10535,32'd10578,32'd10621,32'd10664,32'd10707,32'd10750,32'd10793,32'd10836,32'd10879,32'd10922,32'd10965,32'd11008,32'd11051,32'd11094,32'd11137,32'd11180,32'd11223,32'd11266,32'd11309,32'd11352,32'd11395,32'd11438,32'd11481,32'd11524,32'd11567,32'd11610,32'd11653,32'd11696,32'd11739,32'd11782,32'd11825,32'd11868,32'd11911,32'd11954,32'd11997,32'd12040,32'd12083,32'd12126,32'd12169,32'd12212,32'd12255,32'd12298,32'd12341,32'd12384,32'd12427,32'd12470,32'd12513,32'd12556,32'd12599,32'd12642,32'd12685,32'd12728,32'd12771,32'd12814,32'd12857,32'd12900,32'd12943,32'd12986,32'd13029,32'd13072,32'd13115,32'd13158,32'd13201,32'd13244,32'd13287,32'd13330,32'd13373,32'd13416,32'd13459,32'd13502,32'd13545,32'd13588,32'd13631,32'd13674,32'd13717,32'd13760,32'd13803,32'd13846,32'd13889,32'd13932,32'd13975,32'd14018,32'd14061,32'd14104,32'd14147,32'd14190,32'd14233,32'd14276,32'd14319,32'd14362,32'd14405,32'd14448,32'd14491,32'd14534,32'd14577,32'd14620,32'd14663,32'd14706,32'd14749,32'd14792,32'd14835,32'd14878,32'd14921,32'd14964,32'd15007,32'd15050,32'd15093,32'd15136,32'd15179,32'd15222,32'd15265,32'd15308,32'd15351,32'd15394,32'd15437,32'd15480,32'd15523,32'd15566,32'd15609,32'd15652,32'd15695,32'd15738,32'd15781,32'd15824,32'd15867,32'd15910,32'd15953,32'd15996,32'd16039,32'd16082,32'd16125,32'd16168,32'd16211,32'd16254,32'd16297,32'd16340,32'd16383,32'd16426,32'd16469,32'd16512,32'd16555,32'd16598,32'd16641,32'd16684,32'd16727,32'd16770,32'd16813,32'd16856,32'd16899,32'd16942,32'd16985,32'd17028,32'd17071,32'd17114,32'd17157 };matrix[44]='{32'd0,32'd44,32'd88,32'd132,32'd176,32'd220,32'd264,32'd308,32'd352,32'd396,32'd440,32'd484,32'd528,32'd572,32'd616,32'd660,32'd704,32'd748,32'd792,32'd836,32'd880,32'd924,32'd968,32'd1012,32'd1056,32'd1100,32'd1144,32'd1188,32'd1232,32'd1276,32'd1320,32'd1364,32'd1408,32'd1452,32'd1496,32'd1540,32'd1584,32'd1628,32'd1672,32'd1716,32'd1760,32'd1804,32'd1848,32'd1892,32'd1936,32'd1980,32'd2024,32'd2068,32'd2112,32'd2156,32'd2200,32'd2244,32'd2288,32'd2332,32'd2376,32'd2420,32'd2464,32'd2508,32'd2552,32'd2596,32'd2640,32'd2684,32'd2728,32'd2772,32'd2816,32'd2860,32'd2904,32'd2948,32'd2992,32'd3036,32'd3080,32'd3124,32'd3168,32'd3212,32'd3256,32'd3300,32'd3344,32'd3388,32'd3432,32'd3476,32'd3520,32'd3564,32'd3608,32'd3652,32'd3696,32'd3740,32'd3784,32'd3828,32'd3872,32'd3916,32'd3960,32'd4004,32'd4048,32'd4092,32'd4136,32'd4180,32'd4224,32'd4268,32'd4312,32'd4356,32'd4400,32'd4444,32'd4488,32'd4532,32'd4576,32'd4620,32'd4664,32'd4708,32'd4752,32'd4796,32'd4840,32'd4884,32'd4928,32'd4972,32'd5016,32'd5060,32'd5104,32'd5148,32'd5192,32'd5236,32'd5280,32'd5324,32'd5368,32'd5412,32'd5456,32'd5500,32'd5544,32'd5588,32'd5632,32'd5676,32'd5720,32'd5764,32'd5808,32'd5852,32'd5896,32'd5940,32'd5984,32'd6028,32'd6072,32'd6116,32'd6160,32'd6204,32'd6248,32'd6292,32'd6336,32'd6380,32'd6424,32'd6468,32'd6512,32'd6556,32'd6600,32'd6644,32'd6688,32'd6732,32'd6776,32'd6820,32'd6864,32'd6908,32'd6952,32'd6996,32'd7040,32'd7084,32'd7128,32'd7172,32'd7216,32'd7260,32'd7304,32'd7348,32'd7392,32'd7436,32'd7480,32'd7524,32'd7568,32'd7612,32'd7656,32'd7700,32'd7744,32'd7788,32'd7832,32'd7876,32'd7920,32'd7964,32'd8008,32'd8052,32'd8096,32'd8140,32'd8184,32'd8228,32'd8272,32'd8316,32'd8360,32'd8404,32'd8448,32'd8492,32'd8536,32'd8580,32'd8624,32'd8668,32'd8712,32'd8756,32'd8800,32'd8844,32'd8888,32'd8932,32'd8976,32'd9020,32'd9064,32'd9108,32'd9152,32'd9196,32'd9240,32'd9284,32'd9328,32'd9372,32'd9416,32'd9460,32'd9504,32'd9548,32'd9592,32'd9636,32'd9680,32'd9724,32'd9768,32'd9812,32'd9856,32'd9900,32'd9944,32'd9988,32'd10032,32'd10076,32'd10120,32'd10164,32'd10208,32'd10252,32'd10296,32'd10340,32'd10384,32'd10428,32'd10472,32'd10516,32'd10560,32'd10604,32'd10648,32'd10692,32'd10736,32'd10780,32'd10824,32'd10868,32'd10912,32'd10956,32'd11000,32'd11044,32'd11088,32'd11132,32'd11176,32'd11220,32'd11264,32'd11308,32'd11352,32'd11396,32'd11440,32'd11484,32'd11528,32'd11572,32'd11616,32'd11660,32'd11704,32'd11748,32'd11792,32'd11836,32'd11880,32'd11924,32'd11968,32'd12012,32'd12056,32'd12100,32'd12144,32'd12188,32'd12232,32'd12276,32'd12320,32'd12364,32'd12408,32'd12452,32'd12496,32'd12540,32'd12584,32'd12628,32'd12672,32'd12716,32'd12760,32'd12804,32'd12848,32'd12892,32'd12936,32'd12980,32'd13024,32'd13068,32'd13112,32'd13156,32'd13200,32'd13244,32'd13288,32'd13332,32'd13376,32'd13420,32'd13464,32'd13508,32'd13552,32'd13596,32'd13640,32'd13684,32'd13728,32'd13772,32'd13816,32'd13860,32'd13904,32'd13948,32'd13992,32'd14036,32'd14080,32'd14124,32'd14168,32'd14212,32'd14256,32'd14300,32'd14344,32'd14388,32'd14432,32'd14476,32'd14520,32'd14564,32'd14608,32'd14652,32'd14696,32'd14740,32'd14784,32'd14828,32'd14872,32'd14916,32'd14960,32'd15004,32'd15048,32'd15092,32'd15136,32'd15180,32'd15224,32'd15268,32'd15312,32'd15356,32'd15400,32'd15444,32'd15488,32'd15532,32'd15576,32'd15620,32'd15664,32'd15708,32'd15752,32'd15796,32'd15840,32'd15884,32'd15928,32'd15972,32'd16016,32'd16060,32'd16104,32'd16148,32'd16192,32'd16236,32'd16280,32'd16324,32'd16368,32'd16412,32'd16456,32'd16500,32'd16544,32'd16588,32'd16632,32'd16676,32'd16720,32'd16764,32'd16808,32'd16852,32'd16896,32'd16940,32'd16984,32'd17028,32'd17072,32'd17116,32'd17160,32'd17204,32'd17248,32'd17292,32'd17336,32'd17380,32'd17424,32'd17468,32'd17512,32'd17556 };matrix[45]='{32'd0,32'd45,32'd90,32'd135,32'd180,32'd225,32'd270,32'd315,32'd360,32'd405,32'd450,32'd495,32'd540,32'd585,32'd630,32'd675,32'd720,32'd765,32'd810,32'd855,32'd900,32'd945,32'd990,32'd1035,32'd1080,32'd1125,32'd1170,32'd1215,32'd1260,32'd1305,32'd1350,32'd1395,32'd1440,32'd1485,32'd1530,32'd1575,32'd1620,32'd1665,32'd1710,32'd1755,32'd1800,32'd1845,32'd1890,32'd1935,32'd1980,32'd2025,32'd2070,32'd2115,32'd2160,32'd2205,32'd2250,32'd2295,32'd2340,32'd2385,32'd2430,32'd2475,32'd2520,32'd2565,32'd2610,32'd2655,32'd2700,32'd2745,32'd2790,32'd2835,32'd2880,32'd2925,32'd2970,32'd3015,32'd3060,32'd3105,32'd3150,32'd3195,32'd3240,32'd3285,32'd3330,32'd3375,32'd3420,32'd3465,32'd3510,32'd3555,32'd3600,32'd3645,32'd3690,32'd3735,32'd3780,32'd3825,32'd3870,32'd3915,32'd3960,32'd4005,32'd4050,32'd4095,32'd4140,32'd4185,32'd4230,32'd4275,32'd4320,32'd4365,32'd4410,32'd4455,32'd4500,32'd4545,32'd4590,32'd4635,32'd4680,32'd4725,32'd4770,32'd4815,32'd4860,32'd4905,32'd4950,32'd4995,32'd5040,32'd5085,32'd5130,32'd5175,32'd5220,32'd5265,32'd5310,32'd5355,32'd5400,32'd5445,32'd5490,32'd5535,32'd5580,32'd5625,32'd5670,32'd5715,32'd5760,32'd5805,32'd5850,32'd5895,32'd5940,32'd5985,32'd6030,32'd6075,32'd6120,32'd6165,32'd6210,32'd6255,32'd6300,32'd6345,32'd6390,32'd6435,32'd6480,32'd6525,32'd6570,32'd6615,32'd6660,32'd6705,32'd6750,32'd6795,32'd6840,32'd6885,32'd6930,32'd6975,32'd7020,32'd7065,32'd7110,32'd7155,32'd7200,32'd7245,32'd7290,32'd7335,32'd7380,32'd7425,32'd7470,32'd7515,32'd7560,32'd7605,32'd7650,32'd7695,32'd7740,32'd7785,32'd7830,32'd7875,32'd7920,32'd7965,32'd8010,32'd8055,32'd8100,32'd8145,32'd8190,32'd8235,32'd8280,32'd8325,32'd8370,32'd8415,32'd8460,32'd8505,32'd8550,32'd8595,32'd8640,32'd8685,32'd8730,32'd8775,32'd8820,32'd8865,32'd8910,32'd8955,32'd9000,32'd9045,32'd9090,32'd9135,32'd9180,32'd9225,32'd9270,32'd9315,32'd9360,32'd9405,32'd9450,32'd9495,32'd9540,32'd9585,32'd9630,32'd9675,32'd9720,32'd9765,32'd9810,32'd9855,32'd9900,32'd9945,32'd9990,32'd10035,32'd10080,32'd10125,32'd10170,32'd10215,32'd10260,32'd10305,32'd10350,32'd10395,32'd10440,32'd10485,32'd10530,32'd10575,32'd10620,32'd10665,32'd10710,32'd10755,32'd10800,32'd10845,32'd10890,32'd10935,32'd10980,32'd11025,32'd11070,32'd11115,32'd11160,32'd11205,32'd11250,32'd11295,32'd11340,32'd11385,32'd11430,32'd11475,32'd11520,32'd11565,32'd11610,32'd11655,32'd11700,32'd11745,32'd11790,32'd11835,32'd11880,32'd11925,32'd11970,32'd12015,32'd12060,32'd12105,32'd12150,32'd12195,32'd12240,32'd12285,32'd12330,32'd12375,32'd12420,32'd12465,32'd12510,32'd12555,32'd12600,32'd12645,32'd12690,32'd12735,32'd12780,32'd12825,32'd12870,32'd12915,32'd12960,32'd13005,32'd13050,32'd13095,32'd13140,32'd13185,32'd13230,32'd13275,32'd13320,32'd13365,32'd13410,32'd13455,32'd13500,32'd13545,32'd13590,32'd13635,32'd13680,32'd13725,32'd13770,32'd13815,32'd13860,32'd13905,32'd13950,32'd13995,32'd14040,32'd14085,32'd14130,32'd14175,32'd14220,32'd14265,32'd14310,32'd14355,32'd14400,32'd14445,32'd14490,32'd14535,32'd14580,32'd14625,32'd14670,32'd14715,32'd14760,32'd14805,32'd14850,32'd14895,32'd14940,32'd14985,32'd15030,32'd15075,32'd15120,32'd15165,32'd15210,32'd15255,32'd15300,32'd15345,32'd15390,32'd15435,32'd15480,32'd15525,32'd15570,32'd15615,32'd15660,32'd15705,32'd15750,32'd15795,32'd15840,32'd15885,32'd15930,32'd15975,32'd16020,32'd16065,32'd16110,32'd16155,32'd16200,32'd16245,32'd16290,32'd16335,32'd16380,32'd16425,32'd16470,32'd16515,32'd16560,32'd16605,32'd16650,32'd16695,32'd16740,32'd16785,32'd16830,32'd16875,32'd16920,32'd16965,32'd17010,32'd17055,32'd17100,32'd17145,32'd17190,32'd17235,32'd17280,32'd17325,32'd17370,32'd17415,32'd17460,32'd17505,32'd17550,32'd17595,32'd17640,32'd17685,32'd17730,32'd17775,32'd17820,32'd17865,32'd17910,32'd17955 };matrix[46]='{32'd0,32'd46,32'd92,32'd138,32'd184,32'd230,32'd276,32'd322,32'd368,32'd414,32'd460,32'd506,32'd552,32'd598,32'd644,32'd690,32'd736,32'd782,32'd828,32'd874,32'd920,32'd966,32'd1012,32'd1058,32'd1104,32'd1150,32'd1196,32'd1242,32'd1288,32'd1334,32'd1380,32'd1426,32'd1472,32'd1518,32'd1564,32'd1610,32'd1656,32'd1702,32'd1748,32'd1794,32'd1840,32'd1886,32'd1932,32'd1978,32'd2024,32'd2070,32'd2116,32'd2162,32'd2208,32'd2254,32'd2300,32'd2346,32'd2392,32'd2438,32'd2484,32'd2530,32'd2576,32'd2622,32'd2668,32'd2714,32'd2760,32'd2806,32'd2852,32'd2898,32'd2944,32'd2990,32'd3036,32'd3082,32'd3128,32'd3174,32'd3220,32'd3266,32'd3312,32'd3358,32'd3404,32'd3450,32'd3496,32'd3542,32'd3588,32'd3634,32'd3680,32'd3726,32'd3772,32'd3818,32'd3864,32'd3910,32'd3956,32'd4002,32'd4048,32'd4094,32'd4140,32'd4186,32'd4232,32'd4278,32'd4324,32'd4370,32'd4416,32'd4462,32'd4508,32'd4554,32'd4600,32'd4646,32'd4692,32'd4738,32'd4784,32'd4830,32'd4876,32'd4922,32'd4968,32'd5014,32'd5060,32'd5106,32'd5152,32'd5198,32'd5244,32'd5290,32'd5336,32'd5382,32'd5428,32'd5474,32'd5520,32'd5566,32'd5612,32'd5658,32'd5704,32'd5750,32'd5796,32'd5842,32'd5888,32'd5934,32'd5980,32'd6026,32'd6072,32'd6118,32'd6164,32'd6210,32'd6256,32'd6302,32'd6348,32'd6394,32'd6440,32'd6486,32'd6532,32'd6578,32'd6624,32'd6670,32'd6716,32'd6762,32'd6808,32'd6854,32'd6900,32'd6946,32'd6992,32'd7038,32'd7084,32'd7130,32'd7176,32'd7222,32'd7268,32'd7314,32'd7360,32'd7406,32'd7452,32'd7498,32'd7544,32'd7590,32'd7636,32'd7682,32'd7728,32'd7774,32'd7820,32'd7866,32'd7912,32'd7958,32'd8004,32'd8050,32'd8096,32'd8142,32'd8188,32'd8234,32'd8280,32'd8326,32'd8372,32'd8418,32'd8464,32'd8510,32'd8556,32'd8602,32'd8648,32'd8694,32'd8740,32'd8786,32'd8832,32'd8878,32'd8924,32'd8970,32'd9016,32'd9062,32'd9108,32'd9154,32'd9200,32'd9246,32'd9292,32'd9338,32'd9384,32'd9430,32'd9476,32'd9522,32'd9568,32'd9614,32'd9660,32'd9706,32'd9752,32'd9798,32'd9844,32'd9890,32'd9936,32'd9982,32'd10028,32'd10074,32'd10120,32'd10166,32'd10212,32'd10258,32'd10304,32'd10350,32'd10396,32'd10442,32'd10488,32'd10534,32'd10580,32'd10626,32'd10672,32'd10718,32'd10764,32'd10810,32'd10856,32'd10902,32'd10948,32'd10994,32'd11040,32'd11086,32'd11132,32'd11178,32'd11224,32'd11270,32'd11316,32'd11362,32'd11408,32'd11454,32'd11500,32'd11546,32'd11592,32'd11638,32'd11684,32'd11730,32'd11776,32'd11822,32'd11868,32'd11914,32'd11960,32'd12006,32'd12052,32'd12098,32'd12144,32'd12190,32'd12236,32'd12282,32'd12328,32'd12374,32'd12420,32'd12466,32'd12512,32'd12558,32'd12604,32'd12650,32'd12696,32'd12742,32'd12788,32'd12834,32'd12880,32'd12926,32'd12972,32'd13018,32'd13064,32'd13110,32'd13156,32'd13202,32'd13248,32'd13294,32'd13340,32'd13386,32'd13432,32'd13478,32'd13524,32'd13570,32'd13616,32'd13662,32'd13708,32'd13754,32'd13800,32'd13846,32'd13892,32'd13938,32'd13984,32'd14030,32'd14076,32'd14122,32'd14168,32'd14214,32'd14260,32'd14306,32'd14352,32'd14398,32'd14444,32'd14490,32'd14536,32'd14582,32'd14628,32'd14674,32'd14720,32'd14766,32'd14812,32'd14858,32'd14904,32'd14950,32'd14996,32'd15042,32'd15088,32'd15134,32'd15180,32'd15226,32'd15272,32'd15318,32'd15364,32'd15410,32'd15456,32'd15502,32'd15548,32'd15594,32'd15640,32'd15686,32'd15732,32'd15778,32'd15824,32'd15870,32'd15916,32'd15962,32'd16008,32'd16054,32'd16100,32'd16146,32'd16192,32'd16238,32'd16284,32'd16330,32'd16376,32'd16422,32'd16468,32'd16514,32'd16560,32'd16606,32'd16652,32'd16698,32'd16744,32'd16790,32'd16836,32'd16882,32'd16928,32'd16974,32'd17020,32'd17066,32'd17112,32'd17158,32'd17204,32'd17250,32'd17296,32'd17342,32'd17388,32'd17434,32'd17480,32'd17526,32'd17572,32'd17618,32'd17664,32'd17710,32'd17756,32'd17802,32'd17848,32'd17894,32'd17940,32'd17986,32'd18032,32'd18078,32'd18124,32'd18170,32'd18216,32'd18262,32'd18308,32'd18354 };matrix[47]='{32'd0,32'd47,32'd94,32'd141,32'd188,32'd235,32'd282,32'd329,32'd376,32'd423,32'd470,32'd517,32'd564,32'd611,32'd658,32'd705,32'd752,32'd799,32'd846,32'd893,32'd940,32'd987,32'd1034,32'd1081,32'd1128,32'd1175,32'd1222,32'd1269,32'd1316,32'd1363,32'd1410,32'd1457,32'd1504,32'd1551,32'd1598,32'd1645,32'd1692,32'd1739,32'd1786,32'd1833,32'd1880,32'd1927,32'd1974,32'd2021,32'd2068,32'd2115,32'd2162,32'd2209,32'd2256,32'd2303,32'd2350,32'd2397,32'd2444,32'd2491,32'd2538,32'd2585,32'd2632,32'd2679,32'd2726,32'd2773,32'd2820,32'd2867,32'd2914,32'd2961,32'd3008,32'd3055,32'd3102,32'd3149,32'd3196,32'd3243,32'd3290,32'd3337,32'd3384,32'd3431,32'd3478,32'd3525,32'd3572,32'd3619,32'd3666,32'd3713,32'd3760,32'd3807,32'd3854,32'd3901,32'd3948,32'd3995,32'd4042,32'd4089,32'd4136,32'd4183,32'd4230,32'd4277,32'd4324,32'd4371,32'd4418,32'd4465,32'd4512,32'd4559,32'd4606,32'd4653,32'd4700,32'd4747,32'd4794,32'd4841,32'd4888,32'd4935,32'd4982,32'd5029,32'd5076,32'd5123,32'd5170,32'd5217,32'd5264,32'd5311,32'd5358,32'd5405,32'd5452,32'd5499,32'd5546,32'd5593,32'd5640,32'd5687,32'd5734,32'd5781,32'd5828,32'd5875,32'd5922,32'd5969,32'd6016,32'd6063,32'd6110,32'd6157,32'd6204,32'd6251,32'd6298,32'd6345,32'd6392,32'd6439,32'd6486,32'd6533,32'd6580,32'd6627,32'd6674,32'd6721,32'd6768,32'd6815,32'd6862,32'd6909,32'd6956,32'd7003,32'd7050,32'd7097,32'd7144,32'd7191,32'd7238,32'd7285,32'd7332,32'd7379,32'd7426,32'd7473,32'd7520,32'd7567,32'd7614,32'd7661,32'd7708,32'd7755,32'd7802,32'd7849,32'd7896,32'd7943,32'd7990,32'd8037,32'd8084,32'd8131,32'd8178,32'd8225,32'd8272,32'd8319,32'd8366,32'd8413,32'd8460,32'd8507,32'd8554,32'd8601,32'd8648,32'd8695,32'd8742,32'd8789,32'd8836,32'd8883,32'd8930,32'd8977,32'd9024,32'd9071,32'd9118,32'd9165,32'd9212,32'd9259,32'd9306,32'd9353,32'd9400,32'd9447,32'd9494,32'd9541,32'd9588,32'd9635,32'd9682,32'd9729,32'd9776,32'd9823,32'd9870,32'd9917,32'd9964,32'd10011,32'd10058,32'd10105,32'd10152,32'd10199,32'd10246,32'd10293,32'd10340,32'd10387,32'd10434,32'd10481,32'd10528,32'd10575,32'd10622,32'd10669,32'd10716,32'd10763,32'd10810,32'd10857,32'd10904,32'd10951,32'd10998,32'd11045,32'd11092,32'd11139,32'd11186,32'd11233,32'd11280,32'd11327,32'd11374,32'd11421,32'd11468,32'd11515,32'd11562,32'd11609,32'd11656,32'd11703,32'd11750,32'd11797,32'd11844,32'd11891,32'd11938,32'd11985,32'd12032,32'd12079,32'd12126,32'd12173,32'd12220,32'd12267,32'd12314,32'd12361,32'd12408,32'd12455,32'd12502,32'd12549,32'd12596,32'd12643,32'd12690,32'd12737,32'd12784,32'd12831,32'd12878,32'd12925,32'd12972,32'd13019,32'd13066,32'd13113,32'd13160,32'd13207,32'd13254,32'd13301,32'd13348,32'd13395,32'd13442,32'd13489,32'd13536,32'd13583,32'd13630,32'd13677,32'd13724,32'd13771,32'd13818,32'd13865,32'd13912,32'd13959,32'd14006,32'd14053,32'd14100,32'd14147,32'd14194,32'd14241,32'd14288,32'd14335,32'd14382,32'd14429,32'd14476,32'd14523,32'd14570,32'd14617,32'd14664,32'd14711,32'd14758,32'd14805,32'd14852,32'd14899,32'd14946,32'd14993,32'd15040,32'd15087,32'd15134,32'd15181,32'd15228,32'd15275,32'd15322,32'd15369,32'd15416,32'd15463,32'd15510,32'd15557,32'd15604,32'd15651,32'd15698,32'd15745,32'd15792,32'd15839,32'd15886,32'd15933,32'd15980,32'd16027,32'd16074,32'd16121,32'd16168,32'd16215,32'd16262,32'd16309,32'd16356,32'd16403,32'd16450,32'd16497,32'd16544,32'd16591,32'd16638,32'd16685,32'd16732,32'd16779,32'd16826,32'd16873,32'd16920,32'd16967,32'd17014,32'd17061,32'd17108,32'd17155,32'd17202,32'd17249,32'd17296,32'd17343,32'd17390,32'd17437,32'd17484,32'd17531,32'd17578,32'd17625,32'd17672,32'd17719,32'd17766,32'd17813,32'd17860,32'd17907,32'd17954,32'd18001,32'd18048,32'd18095,32'd18142,32'd18189,32'd18236,32'd18283,32'd18330,32'd18377,32'd18424,32'd18471,32'd18518,32'd18565,32'd18612,32'd18659,32'd18706,32'd18753 };matrix[48]='{32'd0,32'd48,32'd96,32'd144,32'd192,32'd240,32'd288,32'd336,32'd384,32'd432,32'd480,32'd528,32'd576,32'd624,32'd672,32'd720,32'd768,32'd816,32'd864,32'd912,32'd960,32'd1008,32'd1056,32'd1104,32'd1152,32'd1200,32'd1248,32'd1296,32'd1344,32'd1392,32'd1440,32'd1488,32'd1536,32'd1584,32'd1632,32'd1680,32'd1728,32'd1776,32'd1824,32'd1872,32'd1920,32'd1968,32'd2016,32'd2064,32'd2112,32'd2160,32'd2208,32'd2256,32'd2304,32'd2352,32'd2400,32'd2448,32'd2496,32'd2544,32'd2592,32'd2640,32'd2688,32'd2736,32'd2784,32'd2832,32'd2880,32'd2928,32'd2976,32'd3024,32'd3072,32'd3120,32'd3168,32'd3216,32'd3264,32'd3312,32'd3360,32'd3408,32'd3456,32'd3504,32'd3552,32'd3600,32'd3648,32'd3696,32'd3744,32'd3792,32'd3840,32'd3888,32'd3936,32'd3984,32'd4032,32'd4080,32'd4128,32'd4176,32'd4224,32'd4272,32'd4320,32'd4368,32'd4416,32'd4464,32'd4512,32'd4560,32'd4608,32'd4656,32'd4704,32'd4752,32'd4800,32'd4848,32'd4896,32'd4944,32'd4992,32'd5040,32'd5088,32'd5136,32'd5184,32'd5232,32'd5280,32'd5328,32'd5376,32'd5424,32'd5472,32'd5520,32'd5568,32'd5616,32'd5664,32'd5712,32'd5760,32'd5808,32'd5856,32'd5904,32'd5952,32'd6000,32'd6048,32'd6096,32'd6144,32'd6192,32'd6240,32'd6288,32'd6336,32'd6384,32'd6432,32'd6480,32'd6528,32'd6576,32'd6624,32'd6672,32'd6720,32'd6768,32'd6816,32'd6864,32'd6912,32'd6960,32'd7008,32'd7056,32'd7104,32'd7152,32'd7200,32'd7248,32'd7296,32'd7344,32'd7392,32'd7440,32'd7488,32'd7536,32'd7584,32'd7632,32'd7680,32'd7728,32'd7776,32'd7824,32'd7872,32'd7920,32'd7968,32'd8016,32'd8064,32'd8112,32'd8160,32'd8208,32'd8256,32'd8304,32'd8352,32'd8400,32'd8448,32'd8496,32'd8544,32'd8592,32'd8640,32'd8688,32'd8736,32'd8784,32'd8832,32'd8880,32'd8928,32'd8976,32'd9024,32'd9072,32'd9120,32'd9168,32'd9216,32'd9264,32'd9312,32'd9360,32'd9408,32'd9456,32'd9504,32'd9552,32'd9600,32'd9648,32'd9696,32'd9744,32'd9792,32'd9840,32'd9888,32'd9936,32'd9984,32'd10032,32'd10080,32'd10128,32'd10176,32'd10224,32'd10272,32'd10320,32'd10368,32'd10416,32'd10464,32'd10512,32'd10560,32'd10608,32'd10656,32'd10704,32'd10752,32'd10800,32'd10848,32'd10896,32'd10944,32'd10992,32'd11040,32'd11088,32'd11136,32'd11184,32'd11232,32'd11280,32'd11328,32'd11376,32'd11424,32'd11472,32'd11520,32'd11568,32'd11616,32'd11664,32'd11712,32'd11760,32'd11808,32'd11856,32'd11904,32'd11952,32'd12000,32'd12048,32'd12096,32'd12144,32'd12192,32'd12240,32'd12288,32'd12336,32'd12384,32'd12432,32'd12480,32'd12528,32'd12576,32'd12624,32'd12672,32'd12720,32'd12768,32'd12816,32'd12864,32'd12912,32'd12960,32'd13008,32'd13056,32'd13104,32'd13152,32'd13200,32'd13248,32'd13296,32'd13344,32'd13392,32'd13440,32'd13488,32'd13536,32'd13584,32'd13632,32'd13680,32'd13728,32'd13776,32'd13824,32'd13872,32'd13920,32'd13968,32'd14016,32'd14064,32'd14112,32'd14160,32'd14208,32'd14256,32'd14304,32'd14352,32'd14400,32'd14448,32'd14496,32'd14544,32'd14592,32'd14640,32'd14688,32'd14736,32'd14784,32'd14832,32'd14880,32'd14928,32'd14976,32'd15024,32'd15072,32'd15120,32'd15168,32'd15216,32'd15264,32'd15312,32'd15360,32'd15408,32'd15456,32'd15504,32'd15552,32'd15600,32'd15648,32'd15696,32'd15744,32'd15792,32'd15840,32'd15888,32'd15936,32'd15984,32'd16032,32'd16080,32'd16128,32'd16176,32'd16224,32'd16272,32'd16320,32'd16368,32'd16416,32'd16464,32'd16512,32'd16560,32'd16608,32'd16656,32'd16704,32'd16752,32'd16800,32'd16848,32'd16896,32'd16944,32'd16992,32'd17040,32'd17088,32'd17136,32'd17184,32'd17232,32'd17280,32'd17328,32'd17376,32'd17424,32'd17472,32'd17520,32'd17568,32'd17616,32'd17664,32'd17712,32'd17760,32'd17808,32'd17856,32'd17904,32'd17952,32'd18000,32'd18048,32'd18096,32'd18144,32'd18192,32'd18240,32'd18288,32'd18336,32'd18384,32'd18432,32'd18480,32'd18528,32'd18576,32'd18624,32'd18672,32'd18720,32'd18768,32'd18816,32'd18864,32'd18912,32'd18960,32'd19008,32'd19056,32'd19104,32'd19152 };matrix[49]='{32'd0,32'd49,32'd98,32'd147,32'd196,32'd245,32'd294,32'd343,32'd392,32'd441,32'd490,32'd539,32'd588,32'd637,32'd686,32'd735,32'd784,32'd833,32'd882,32'd931,32'd980,32'd1029,32'd1078,32'd1127,32'd1176,32'd1225,32'd1274,32'd1323,32'd1372,32'd1421,32'd1470,32'd1519,32'd1568,32'd1617,32'd1666,32'd1715,32'd1764,32'd1813,32'd1862,32'd1911,32'd1960,32'd2009,32'd2058,32'd2107,32'd2156,32'd2205,32'd2254,32'd2303,32'd2352,32'd2401,32'd2450,32'd2499,32'd2548,32'd2597,32'd2646,32'd2695,32'd2744,32'd2793,32'd2842,32'd2891,32'd2940,32'd2989,32'd3038,32'd3087,32'd3136,32'd3185,32'd3234,32'd3283,32'd3332,32'd3381,32'd3430,32'd3479,32'd3528,32'd3577,32'd3626,32'd3675,32'd3724,32'd3773,32'd3822,32'd3871,32'd3920,32'd3969,32'd4018,32'd4067,32'd4116,32'd4165,32'd4214,32'd4263,32'd4312,32'd4361,32'd4410,32'd4459,32'd4508,32'd4557,32'd4606,32'd4655,32'd4704,32'd4753,32'd4802,32'd4851,32'd4900,32'd4949,32'd4998,32'd5047,32'd5096,32'd5145,32'd5194,32'd5243,32'd5292,32'd5341,32'd5390,32'd5439,32'd5488,32'd5537,32'd5586,32'd5635,32'd5684,32'd5733,32'd5782,32'd5831,32'd5880,32'd5929,32'd5978,32'd6027,32'd6076,32'd6125,32'd6174,32'd6223,32'd6272,32'd6321,32'd6370,32'd6419,32'd6468,32'd6517,32'd6566,32'd6615,32'd6664,32'd6713,32'd6762,32'd6811,32'd6860,32'd6909,32'd6958,32'd7007,32'd7056,32'd7105,32'd7154,32'd7203,32'd7252,32'd7301,32'd7350,32'd7399,32'd7448,32'd7497,32'd7546,32'd7595,32'd7644,32'd7693,32'd7742,32'd7791,32'd7840,32'd7889,32'd7938,32'd7987,32'd8036,32'd8085,32'd8134,32'd8183,32'd8232,32'd8281,32'd8330,32'd8379,32'd8428,32'd8477,32'd8526,32'd8575,32'd8624,32'd8673,32'd8722,32'd8771,32'd8820,32'd8869,32'd8918,32'd8967,32'd9016,32'd9065,32'd9114,32'd9163,32'd9212,32'd9261,32'd9310,32'd9359,32'd9408,32'd9457,32'd9506,32'd9555,32'd9604,32'd9653,32'd9702,32'd9751,32'd9800,32'd9849,32'd9898,32'd9947,32'd9996,32'd10045,32'd10094,32'd10143,32'd10192,32'd10241,32'd10290,32'd10339,32'd10388,32'd10437,32'd10486,32'd10535,32'd10584,32'd10633,32'd10682,32'd10731,32'd10780,32'd10829,32'd10878,32'd10927,32'd10976,32'd11025,32'd11074,32'd11123,32'd11172,32'd11221,32'd11270,32'd11319,32'd11368,32'd11417,32'd11466,32'd11515,32'd11564,32'd11613,32'd11662,32'd11711,32'd11760,32'd11809,32'd11858,32'd11907,32'd11956,32'd12005,32'd12054,32'd12103,32'd12152,32'd12201,32'd12250,32'd12299,32'd12348,32'd12397,32'd12446,32'd12495,32'd12544,32'd12593,32'd12642,32'd12691,32'd12740,32'd12789,32'd12838,32'd12887,32'd12936,32'd12985,32'd13034,32'd13083,32'd13132,32'd13181,32'd13230,32'd13279,32'd13328,32'd13377,32'd13426,32'd13475,32'd13524,32'd13573,32'd13622,32'd13671,32'd13720,32'd13769,32'd13818,32'd13867,32'd13916,32'd13965,32'd14014,32'd14063,32'd14112,32'd14161,32'd14210,32'd14259,32'd14308,32'd14357,32'd14406,32'd14455,32'd14504,32'd14553,32'd14602,32'd14651,32'd14700,32'd14749,32'd14798,32'd14847,32'd14896,32'd14945,32'd14994,32'd15043,32'd15092,32'd15141,32'd15190,32'd15239,32'd15288,32'd15337,32'd15386,32'd15435,32'd15484,32'd15533,32'd15582,32'd15631,32'd15680,32'd15729,32'd15778,32'd15827,32'd15876,32'd15925,32'd15974,32'd16023,32'd16072,32'd16121,32'd16170,32'd16219,32'd16268,32'd16317,32'd16366,32'd16415,32'd16464,32'd16513,32'd16562,32'd16611,32'd16660,32'd16709,32'd16758,32'd16807,32'd16856,32'd16905,32'd16954,32'd17003,32'd17052,32'd17101,32'd17150,32'd17199,32'd17248,32'd17297,32'd17346,32'd17395,32'd17444,32'd17493,32'd17542,32'd17591,32'd17640,32'd17689,32'd17738,32'd17787,32'd17836,32'd17885,32'd17934,32'd17983,32'd18032,32'd18081,32'd18130,32'd18179,32'd18228,32'd18277,32'd18326,32'd18375,32'd18424,32'd18473,32'd18522,32'd18571,32'd18620,32'd18669,32'd18718,32'd18767,32'd18816,32'd18865,32'd18914,32'd18963,32'd19012,32'd19061,32'd19110,32'd19159,32'd19208,32'd19257,32'd19306,32'd19355,32'd19404,32'd19453,32'd19502,32'd19551 };matrix[50]='{32'd0,32'd50,32'd100,32'd150,32'd200,32'd250,32'd300,32'd350,32'd400,32'd450,32'd500,32'd550,32'd600,32'd650,32'd700,32'd750,32'd800,32'd850,32'd900,32'd950,32'd1000,32'd1050,32'd1100,32'd1150,32'd1200,32'd1250,32'd1300,32'd1350,32'd1400,32'd1450,32'd1500,32'd1550,32'd1600,32'd1650,32'd1700,32'd1750,32'd1800,32'd1850,32'd1900,32'd1950,32'd2000,32'd2050,32'd2100,32'd2150,32'd2200,32'd2250,32'd2300,32'd2350,32'd2400,32'd2450,32'd2500,32'd2550,32'd2600,32'd2650,32'd2700,32'd2750,32'd2800,32'd2850,32'd2900,32'd2950,32'd3000,32'd3050,32'd3100,32'd3150,32'd3200,32'd3250,32'd3300,32'd3350,32'd3400,32'd3450,32'd3500,32'd3550,32'd3600,32'd3650,32'd3700,32'd3750,32'd3800,32'd3850,32'd3900,32'd3950,32'd4000,32'd4050,32'd4100,32'd4150,32'd4200,32'd4250,32'd4300,32'd4350,32'd4400,32'd4450,32'd4500,32'd4550,32'd4600,32'd4650,32'd4700,32'd4750,32'd4800,32'd4850,32'd4900,32'd4950,32'd5000,32'd5050,32'd5100,32'd5150,32'd5200,32'd5250,32'd5300,32'd5350,32'd5400,32'd5450,32'd5500,32'd5550,32'd5600,32'd5650,32'd5700,32'd5750,32'd5800,32'd5850,32'd5900,32'd5950,32'd6000,32'd6050,32'd6100,32'd6150,32'd6200,32'd6250,32'd6300,32'd6350,32'd6400,32'd6450,32'd6500,32'd6550,32'd6600,32'd6650,32'd6700,32'd6750,32'd6800,32'd6850,32'd6900,32'd6950,32'd7000,32'd7050,32'd7100,32'd7150,32'd7200,32'd7250,32'd7300,32'd7350,32'd7400,32'd7450,32'd7500,32'd7550,32'd7600,32'd7650,32'd7700,32'd7750,32'd7800,32'd7850,32'd7900,32'd7950,32'd8000,32'd8050,32'd8100,32'd8150,32'd8200,32'd8250,32'd8300,32'd8350,32'd8400,32'd8450,32'd8500,32'd8550,32'd8600,32'd8650,32'd8700,32'd8750,32'd8800,32'd8850,32'd8900,32'd8950,32'd9000,32'd9050,32'd9100,32'd9150,32'd9200,32'd9250,32'd9300,32'd9350,32'd9400,32'd9450,32'd9500,32'd9550,32'd9600,32'd9650,32'd9700,32'd9750,32'd9800,32'd9850,32'd9900,32'd9950,32'd10000,32'd10050,32'd10100,32'd10150,32'd10200,32'd10250,32'd10300,32'd10350,32'd10400,32'd10450,32'd10500,32'd10550,32'd10600,32'd10650,32'd10700,32'd10750,32'd10800,32'd10850,32'd10900,32'd10950,32'd11000,32'd11050,32'd11100,32'd11150,32'd11200,32'd11250,32'd11300,32'd11350,32'd11400,32'd11450,32'd11500,32'd11550,32'd11600,32'd11650,32'd11700,32'd11750,32'd11800,32'd11850,32'd11900,32'd11950,32'd12000,32'd12050,32'd12100,32'd12150,32'd12200,32'd12250,32'd12300,32'd12350,32'd12400,32'd12450,32'd12500,32'd12550,32'd12600,32'd12650,32'd12700,32'd12750,32'd12800,32'd12850,32'd12900,32'd12950,32'd13000,32'd13050,32'd13100,32'd13150,32'd13200,32'd13250,32'd13300,32'd13350,32'd13400,32'd13450,32'd13500,32'd13550,32'd13600,32'd13650,32'd13700,32'd13750,32'd13800,32'd13850,32'd13900,32'd13950,32'd14000,32'd14050,32'd14100,32'd14150,32'd14200,32'd14250,32'd14300,32'd14350,32'd14400,32'd14450,32'd14500,32'd14550,32'd14600,32'd14650,32'd14700,32'd14750,32'd14800,32'd14850,32'd14900,32'd14950,32'd15000,32'd15050,32'd15100,32'd15150,32'd15200,32'd15250,32'd15300,32'd15350,32'd15400,32'd15450,32'd15500,32'd15550,32'd15600,32'd15650,32'd15700,32'd15750,32'd15800,32'd15850,32'd15900,32'd15950,32'd16000,32'd16050,32'd16100,32'd16150,32'd16200,32'd16250,32'd16300,32'd16350,32'd16400,32'd16450,32'd16500,32'd16550,32'd16600,32'd16650,32'd16700,32'd16750,32'd16800,32'd16850,32'd16900,32'd16950,32'd17000,32'd17050,32'd17100,32'd17150,32'd17200,32'd17250,32'd17300,32'd17350,32'd17400,32'd17450,32'd17500,32'd17550,32'd17600,32'd17650,32'd17700,32'd17750,32'd17800,32'd17850,32'd17900,32'd17950,32'd18000,32'd18050,32'd18100,32'd18150,32'd18200,32'd18250,32'd18300,32'd18350,32'd18400,32'd18450,32'd18500,32'd18550,32'd18600,32'd18650,32'd18700,32'd18750,32'd18800,32'd18850,32'd18900,32'd18950,32'd19000,32'd19050,32'd19100,32'd19150,32'd19200,32'd19250,32'd19300,32'd19350,32'd19400,32'd19450,32'd19500,32'd19550,32'd19600,32'd19650,32'd19700,32'd19750,32'd19800,32'd19850,32'd19900,32'd19950 };matrix[51]='{32'd0,32'd51,32'd102,32'd153,32'd204,32'd255,32'd306,32'd357,32'd408,32'd459,32'd510,32'd561,32'd612,32'd663,32'd714,32'd765,32'd816,32'd867,32'd918,32'd969,32'd1020,32'd1071,32'd1122,32'd1173,32'd1224,32'd1275,32'd1326,32'd1377,32'd1428,32'd1479,32'd1530,32'd1581,32'd1632,32'd1683,32'd1734,32'd1785,32'd1836,32'd1887,32'd1938,32'd1989,32'd2040,32'd2091,32'd2142,32'd2193,32'd2244,32'd2295,32'd2346,32'd2397,32'd2448,32'd2499,32'd2550,32'd2601,32'd2652,32'd2703,32'd2754,32'd2805,32'd2856,32'd2907,32'd2958,32'd3009,32'd3060,32'd3111,32'd3162,32'd3213,32'd3264,32'd3315,32'd3366,32'd3417,32'd3468,32'd3519,32'd3570,32'd3621,32'd3672,32'd3723,32'd3774,32'd3825,32'd3876,32'd3927,32'd3978,32'd4029,32'd4080,32'd4131,32'd4182,32'd4233,32'd4284,32'd4335,32'd4386,32'd4437,32'd4488,32'd4539,32'd4590,32'd4641,32'd4692,32'd4743,32'd4794,32'd4845,32'd4896,32'd4947,32'd4998,32'd5049,32'd5100,32'd5151,32'd5202,32'd5253,32'd5304,32'd5355,32'd5406,32'd5457,32'd5508,32'd5559,32'd5610,32'd5661,32'd5712,32'd5763,32'd5814,32'd5865,32'd5916,32'd5967,32'd6018,32'd6069,32'd6120,32'd6171,32'd6222,32'd6273,32'd6324,32'd6375,32'd6426,32'd6477,32'd6528,32'd6579,32'd6630,32'd6681,32'd6732,32'd6783,32'd6834,32'd6885,32'd6936,32'd6987,32'd7038,32'd7089,32'd7140,32'd7191,32'd7242,32'd7293,32'd7344,32'd7395,32'd7446,32'd7497,32'd7548,32'd7599,32'd7650,32'd7701,32'd7752,32'd7803,32'd7854,32'd7905,32'd7956,32'd8007,32'd8058,32'd8109,32'd8160,32'd8211,32'd8262,32'd8313,32'd8364,32'd8415,32'd8466,32'd8517,32'd8568,32'd8619,32'd8670,32'd8721,32'd8772,32'd8823,32'd8874,32'd8925,32'd8976,32'd9027,32'd9078,32'd9129,32'd9180,32'd9231,32'd9282,32'd9333,32'd9384,32'd9435,32'd9486,32'd9537,32'd9588,32'd9639,32'd9690,32'd9741,32'd9792,32'd9843,32'd9894,32'd9945,32'd9996,32'd10047,32'd10098,32'd10149,32'd10200,32'd10251,32'd10302,32'd10353,32'd10404,32'd10455,32'd10506,32'd10557,32'd10608,32'd10659,32'd10710,32'd10761,32'd10812,32'd10863,32'd10914,32'd10965,32'd11016,32'd11067,32'd11118,32'd11169,32'd11220,32'd11271,32'd11322,32'd11373,32'd11424,32'd11475,32'd11526,32'd11577,32'd11628,32'd11679,32'd11730,32'd11781,32'd11832,32'd11883,32'd11934,32'd11985,32'd12036,32'd12087,32'd12138,32'd12189,32'd12240,32'd12291,32'd12342,32'd12393,32'd12444,32'd12495,32'd12546,32'd12597,32'd12648,32'd12699,32'd12750,32'd12801,32'd12852,32'd12903,32'd12954,32'd13005,32'd13056,32'd13107,32'd13158,32'd13209,32'd13260,32'd13311,32'd13362,32'd13413,32'd13464,32'd13515,32'd13566,32'd13617,32'd13668,32'd13719,32'd13770,32'd13821,32'd13872,32'd13923,32'd13974,32'd14025,32'd14076,32'd14127,32'd14178,32'd14229,32'd14280,32'd14331,32'd14382,32'd14433,32'd14484,32'd14535,32'd14586,32'd14637,32'd14688,32'd14739,32'd14790,32'd14841,32'd14892,32'd14943,32'd14994,32'd15045,32'd15096,32'd15147,32'd15198,32'd15249,32'd15300,32'd15351,32'd15402,32'd15453,32'd15504,32'd15555,32'd15606,32'd15657,32'd15708,32'd15759,32'd15810,32'd15861,32'd15912,32'd15963,32'd16014,32'd16065,32'd16116,32'd16167,32'd16218,32'd16269,32'd16320,32'd16371,32'd16422,32'd16473,32'd16524,32'd16575,32'd16626,32'd16677,32'd16728,32'd16779,32'd16830,32'd16881,32'd16932,32'd16983,32'd17034,32'd17085,32'd17136,32'd17187,32'd17238,32'd17289,32'd17340,32'd17391,32'd17442,32'd17493,32'd17544,32'd17595,32'd17646,32'd17697,32'd17748,32'd17799,32'd17850,32'd17901,32'd17952,32'd18003,32'd18054,32'd18105,32'd18156,32'd18207,32'd18258,32'd18309,32'd18360,32'd18411,32'd18462,32'd18513,32'd18564,32'd18615,32'd18666,32'd18717,32'd18768,32'd18819,32'd18870,32'd18921,32'd18972,32'd19023,32'd19074,32'd19125,32'd19176,32'd19227,32'd19278,32'd19329,32'd19380,32'd19431,32'd19482,32'd19533,32'd19584,32'd19635,32'd19686,32'd19737,32'd19788,32'd19839,32'd19890,32'd19941,32'd19992,32'd20043,32'd20094,32'd20145,32'd20196,32'd20247,32'd20298,32'd20349 };matrix[52]='{32'd0,32'd52,32'd104,32'd156,32'd208,32'd260,32'd312,32'd364,32'd416,32'd468,32'd520,32'd572,32'd624,32'd676,32'd728,32'd780,32'd832,32'd884,32'd936,32'd988,32'd1040,32'd1092,32'd1144,32'd1196,32'd1248,32'd1300,32'd1352,32'd1404,32'd1456,32'd1508,32'd1560,32'd1612,32'd1664,32'd1716,32'd1768,32'd1820,32'd1872,32'd1924,32'd1976,32'd2028,32'd2080,32'd2132,32'd2184,32'd2236,32'd2288,32'd2340,32'd2392,32'd2444,32'd2496,32'd2548,32'd2600,32'd2652,32'd2704,32'd2756,32'd2808,32'd2860,32'd2912,32'd2964,32'd3016,32'd3068,32'd3120,32'd3172,32'd3224,32'd3276,32'd3328,32'd3380,32'd3432,32'd3484,32'd3536,32'd3588,32'd3640,32'd3692,32'd3744,32'd3796,32'd3848,32'd3900,32'd3952,32'd4004,32'd4056,32'd4108,32'd4160,32'd4212,32'd4264,32'd4316,32'd4368,32'd4420,32'd4472,32'd4524,32'd4576,32'd4628,32'd4680,32'd4732,32'd4784,32'd4836,32'd4888,32'd4940,32'd4992,32'd5044,32'd5096,32'd5148,32'd5200,32'd5252,32'd5304,32'd5356,32'd5408,32'd5460,32'd5512,32'd5564,32'd5616,32'd5668,32'd5720,32'd5772,32'd5824,32'd5876,32'd5928,32'd5980,32'd6032,32'd6084,32'd6136,32'd6188,32'd6240,32'd6292,32'd6344,32'd6396,32'd6448,32'd6500,32'd6552,32'd6604,32'd6656,32'd6708,32'd6760,32'd6812,32'd6864,32'd6916,32'd6968,32'd7020,32'd7072,32'd7124,32'd7176,32'd7228,32'd7280,32'd7332,32'd7384,32'd7436,32'd7488,32'd7540,32'd7592,32'd7644,32'd7696,32'd7748,32'd7800,32'd7852,32'd7904,32'd7956,32'd8008,32'd8060,32'd8112,32'd8164,32'd8216,32'd8268,32'd8320,32'd8372,32'd8424,32'd8476,32'd8528,32'd8580,32'd8632,32'd8684,32'd8736,32'd8788,32'd8840,32'd8892,32'd8944,32'd8996,32'd9048,32'd9100,32'd9152,32'd9204,32'd9256,32'd9308,32'd9360,32'd9412,32'd9464,32'd9516,32'd9568,32'd9620,32'd9672,32'd9724,32'd9776,32'd9828,32'd9880,32'd9932,32'd9984,32'd10036,32'd10088,32'd10140,32'd10192,32'd10244,32'd10296,32'd10348,32'd10400,32'd10452,32'd10504,32'd10556,32'd10608,32'd10660,32'd10712,32'd10764,32'd10816,32'd10868,32'd10920,32'd10972,32'd11024,32'd11076,32'd11128,32'd11180,32'd11232,32'd11284,32'd11336,32'd11388,32'd11440,32'd11492,32'd11544,32'd11596,32'd11648,32'd11700,32'd11752,32'd11804,32'd11856,32'd11908,32'd11960,32'd12012,32'd12064,32'd12116,32'd12168,32'd12220,32'd12272,32'd12324,32'd12376,32'd12428,32'd12480,32'd12532,32'd12584,32'd12636,32'd12688,32'd12740,32'd12792,32'd12844,32'd12896,32'd12948,32'd13000,32'd13052,32'd13104,32'd13156,32'd13208,32'd13260,32'd13312,32'd13364,32'd13416,32'd13468,32'd13520,32'd13572,32'd13624,32'd13676,32'd13728,32'd13780,32'd13832,32'd13884,32'd13936,32'd13988,32'd14040,32'd14092,32'd14144,32'd14196,32'd14248,32'd14300,32'd14352,32'd14404,32'd14456,32'd14508,32'd14560,32'd14612,32'd14664,32'd14716,32'd14768,32'd14820,32'd14872,32'd14924,32'd14976,32'd15028,32'd15080,32'd15132,32'd15184,32'd15236,32'd15288,32'd15340,32'd15392,32'd15444,32'd15496,32'd15548,32'd15600,32'd15652,32'd15704,32'd15756,32'd15808,32'd15860,32'd15912,32'd15964,32'd16016,32'd16068,32'd16120,32'd16172,32'd16224,32'd16276,32'd16328,32'd16380,32'd16432,32'd16484,32'd16536,32'd16588,32'd16640,32'd16692,32'd16744,32'd16796,32'd16848,32'd16900,32'd16952,32'd17004,32'd17056,32'd17108,32'd17160,32'd17212,32'd17264,32'd17316,32'd17368,32'd17420,32'd17472,32'd17524,32'd17576,32'd17628,32'd17680,32'd17732,32'd17784,32'd17836,32'd17888,32'd17940,32'd17992,32'd18044,32'd18096,32'd18148,32'd18200,32'd18252,32'd18304,32'd18356,32'd18408,32'd18460,32'd18512,32'd18564,32'd18616,32'd18668,32'd18720,32'd18772,32'd18824,32'd18876,32'd18928,32'd18980,32'd19032,32'd19084,32'd19136,32'd19188,32'd19240,32'd19292,32'd19344,32'd19396,32'd19448,32'd19500,32'd19552,32'd19604,32'd19656,32'd19708,32'd19760,32'd19812,32'd19864,32'd19916,32'd19968,32'd20020,32'd20072,32'd20124,32'd20176,32'd20228,32'd20280,32'd20332,32'd20384,32'd20436,32'd20488,32'd20540,32'd20592,32'd20644,32'd20696,32'd20748 };matrix[53]='{32'd0,32'd53,32'd106,32'd159,32'd212,32'd265,32'd318,32'd371,32'd424,32'd477,32'd530,32'd583,32'd636,32'd689,32'd742,32'd795,32'd848,32'd901,32'd954,32'd1007,32'd1060,32'd1113,32'd1166,32'd1219,32'd1272,32'd1325,32'd1378,32'd1431,32'd1484,32'd1537,32'd1590,32'd1643,32'd1696,32'd1749,32'd1802,32'd1855,32'd1908,32'd1961,32'd2014,32'd2067,32'd2120,32'd2173,32'd2226,32'd2279,32'd2332,32'd2385,32'd2438,32'd2491,32'd2544,32'd2597,32'd2650,32'd2703,32'd2756,32'd2809,32'd2862,32'd2915,32'd2968,32'd3021,32'd3074,32'd3127,32'd3180,32'd3233,32'd3286,32'd3339,32'd3392,32'd3445,32'd3498,32'd3551,32'd3604,32'd3657,32'd3710,32'd3763,32'd3816,32'd3869,32'd3922,32'd3975,32'd4028,32'd4081,32'd4134,32'd4187,32'd4240,32'd4293,32'd4346,32'd4399,32'd4452,32'd4505,32'd4558,32'd4611,32'd4664,32'd4717,32'd4770,32'd4823,32'd4876,32'd4929,32'd4982,32'd5035,32'd5088,32'd5141,32'd5194,32'd5247,32'd5300,32'd5353,32'd5406,32'd5459,32'd5512,32'd5565,32'd5618,32'd5671,32'd5724,32'd5777,32'd5830,32'd5883,32'd5936,32'd5989,32'd6042,32'd6095,32'd6148,32'd6201,32'd6254,32'd6307,32'd6360,32'd6413,32'd6466,32'd6519,32'd6572,32'd6625,32'd6678,32'd6731,32'd6784,32'd6837,32'd6890,32'd6943,32'd6996,32'd7049,32'd7102,32'd7155,32'd7208,32'd7261,32'd7314,32'd7367,32'd7420,32'd7473,32'd7526,32'd7579,32'd7632,32'd7685,32'd7738,32'd7791,32'd7844,32'd7897,32'd7950,32'd8003,32'd8056,32'd8109,32'd8162,32'd8215,32'd8268,32'd8321,32'd8374,32'd8427,32'd8480,32'd8533,32'd8586,32'd8639,32'd8692,32'd8745,32'd8798,32'd8851,32'd8904,32'd8957,32'd9010,32'd9063,32'd9116,32'd9169,32'd9222,32'd9275,32'd9328,32'd9381,32'd9434,32'd9487,32'd9540,32'd9593,32'd9646,32'd9699,32'd9752,32'd9805,32'd9858,32'd9911,32'd9964,32'd10017,32'd10070,32'd10123,32'd10176,32'd10229,32'd10282,32'd10335,32'd10388,32'd10441,32'd10494,32'd10547,32'd10600,32'd10653,32'd10706,32'd10759,32'd10812,32'd10865,32'd10918,32'd10971,32'd11024,32'd11077,32'd11130,32'd11183,32'd11236,32'd11289,32'd11342,32'd11395,32'd11448,32'd11501,32'd11554,32'd11607,32'd11660,32'd11713,32'd11766,32'd11819,32'd11872,32'd11925,32'd11978,32'd12031,32'd12084,32'd12137,32'd12190,32'd12243,32'd12296,32'd12349,32'd12402,32'd12455,32'd12508,32'd12561,32'd12614,32'd12667,32'd12720,32'd12773,32'd12826,32'd12879,32'd12932,32'd12985,32'd13038,32'd13091,32'd13144,32'd13197,32'd13250,32'd13303,32'd13356,32'd13409,32'd13462,32'd13515,32'd13568,32'd13621,32'd13674,32'd13727,32'd13780,32'd13833,32'd13886,32'd13939,32'd13992,32'd14045,32'd14098,32'd14151,32'd14204,32'd14257,32'd14310,32'd14363,32'd14416,32'd14469,32'd14522,32'd14575,32'd14628,32'd14681,32'd14734,32'd14787,32'd14840,32'd14893,32'd14946,32'd14999,32'd15052,32'd15105,32'd15158,32'd15211,32'd15264,32'd15317,32'd15370,32'd15423,32'd15476,32'd15529,32'd15582,32'd15635,32'd15688,32'd15741,32'd15794,32'd15847,32'd15900,32'd15953,32'd16006,32'd16059,32'd16112,32'd16165,32'd16218,32'd16271,32'd16324,32'd16377,32'd16430,32'd16483,32'd16536,32'd16589,32'd16642,32'd16695,32'd16748,32'd16801,32'd16854,32'd16907,32'd16960,32'd17013,32'd17066,32'd17119,32'd17172,32'd17225,32'd17278,32'd17331,32'd17384,32'd17437,32'd17490,32'd17543,32'd17596,32'd17649,32'd17702,32'd17755,32'd17808,32'd17861,32'd17914,32'd17967,32'd18020,32'd18073,32'd18126,32'd18179,32'd18232,32'd18285,32'd18338,32'd18391,32'd18444,32'd18497,32'd18550,32'd18603,32'd18656,32'd18709,32'd18762,32'd18815,32'd18868,32'd18921,32'd18974,32'd19027,32'd19080,32'd19133,32'd19186,32'd19239,32'd19292,32'd19345,32'd19398,32'd19451,32'd19504,32'd19557,32'd19610,32'd19663,32'd19716,32'd19769,32'd19822,32'd19875,32'd19928,32'd19981,32'd20034,32'd20087,32'd20140,32'd20193,32'd20246,32'd20299,32'd20352,32'd20405,32'd20458,32'd20511,32'd20564,32'd20617,32'd20670,32'd20723,32'd20776,32'd20829,32'd20882,32'd20935,32'd20988,32'd21041,32'd21094,32'd21147 };matrix[54]='{32'd0,32'd54,32'd108,32'd162,32'd216,32'd270,32'd324,32'd378,32'd432,32'd486,32'd540,32'd594,32'd648,32'd702,32'd756,32'd810,32'd864,32'd918,32'd972,32'd1026,32'd1080,32'd1134,32'd1188,32'd1242,32'd1296,32'd1350,32'd1404,32'd1458,32'd1512,32'd1566,32'd1620,32'd1674,32'd1728,32'd1782,32'd1836,32'd1890,32'd1944,32'd1998,32'd2052,32'd2106,32'd2160,32'd2214,32'd2268,32'd2322,32'd2376,32'd2430,32'd2484,32'd2538,32'd2592,32'd2646,32'd2700,32'd2754,32'd2808,32'd2862,32'd2916,32'd2970,32'd3024,32'd3078,32'd3132,32'd3186,32'd3240,32'd3294,32'd3348,32'd3402,32'd3456,32'd3510,32'd3564,32'd3618,32'd3672,32'd3726,32'd3780,32'd3834,32'd3888,32'd3942,32'd3996,32'd4050,32'd4104,32'd4158,32'd4212,32'd4266,32'd4320,32'd4374,32'd4428,32'd4482,32'd4536,32'd4590,32'd4644,32'd4698,32'd4752,32'd4806,32'd4860,32'd4914,32'd4968,32'd5022,32'd5076,32'd5130,32'd5184,32'd5238,32'd5292,32'd5346,32'd5400,32'd5454,32'd5508,32'd5562,32'd5616,32'd5670,32'd5724,32'd5778,32'd5832,32'd5886,32'd5940,32'd5994,32'd6048,32'd6102,32'd6156,32'd6210,32'd6264,32'd6318,32'd6372,32'd6426,32'd6480,32'd6534,32'd6588,32'd6642,32'd6696,32'd6750,32'd6804,32'd6858,32'd6912,32'd6966,32'd7020,32'd7074,32'd7128,32'd7182,32'd7236,32'd7290,32'd7344,32'd7398,32'd7452,32'd7506,32'd7560,32'd7614,32'd7668,32'd7722,32'd7776,32'd7830,32'd7884,32'd7938,32'd7992,32'd8046,32'd8100,32'd8154,32'd8208,32'd8262,32'd8316,32'd8370,32'd8424,32'd8478,32'd8532,32'd8586,32'd8640,32'd8694,32'd8748,32'd8802,32'd8856,32'd8910,32'd8964,32'd9018,32'd9072,32'd9126,32'd9180,32'd9234,32'd9288,32'd9342,32'd9396,32'd9450,32'd9504,32'd9558,32'd9612,32'd9666,32'd9720,32'd9774,32'd9828,32'd9882,32'd9936,32'd9990,32'd10044,32'd10098,32'd10152,32'd10206,32'd10260,32'd10314,32'd10368,32'd10422,32'd10476,32'd10530,32'd10584,32'd10638,32'd10692,32'd10746,32'd10800,32'd10854,32'd10908,32'd10962,32'd11016,32'd11070,32'd11124,32'd11178,32'd11232,32'd11286,32'd11340,32'd11394,32'd11448,32'd11502,32'd11556,32'd11610,32'd11664,32'd11718,32'd11772,32'd11826,32'd11880,32'd11934,32'd11988,32'd12042,32'd12096,32'd12150,32'd12204,32'd12258,32'd12312,32'd12366,32'd12420,32'd12474,32'd12528,32'd12582,32'd12636,32'd12690,32'd12744,32'd12798,32'd12852,32'd12906,32'd12960,32'd13014,32'd13068,32'd13122,32'd13176,32'd13230,32'd13284,32'd13338,32'd13392,32'd13446,32'd13500,32'd13554,32'd13608,32'd13662,32'd13716,32'd13770,32'd13824,32'd13878,32'd13932,32'd13986,32'd14040,32'd14094,32'd14148,32'd14202,32'd14256,32'd14310,32'd14364,32'd14418,32'd14472,32'd14526,32'd14580,32'd14634,32'd14688,32'd14742,32'd14796,32'd14850,32'd14904,32'd14958,32'd15012,32'd15066,32'd15120,32'd15174,32'd15228,32'd15282,32'd15336,32'd15390,32'd15444,32'd15498,32'd15552,32'd15606,32'd15660,32'd15714,32'd15768,32'd15822,32'd15876,32'd15930,32'd15984,32'd16038,32'd16092,32'd16146,32'd16200,32'd16254,32'd16308,32'd16362,32'd16416,32'd16470,32'd16524,32'd16578,32'd16632,32'd16686,32'd16740,32'd16794,32'd16848,32'd16902,32'd16956,32'd17010,32'd17064,32'd17118,32'd17172,32'd17226,32'd17280,32'd17334,32'd17388,32'd17442,32'd17496,32'd17550,32'd17604,32'd17658,32'd17712,32'd17766,32'd17820,32'd17874,32'd17928,32'd17982,32'd18036,32'd18090,32'd18144,32'd18198,32'd18252,32'd18306,32'd18360,32'd18414,32'd18468,32'd18522,32'd18576,32'd18630,32'd18684,32'd18738,32'd18792,32'd18846,32'd18900,32'd18954,32'd19008,32'd19062,32'd19116,32'd19170,32'd19224,32'd19278,32'd19332,32'd19386,32'd19440,32'd19494,32'd19548,32'd19602,32'd19656,32'd19710,32'd19764,32'd19818,32'd19872,32'd19926,32'd19980,32'd20034,32'd20088,32'd20142,32'd20196,32'd20250,32'd20304,32'd20358,32'd20412,32'd20466,32'd20520,32'd20574,32'd20628,32'd20682,32'd20736,32'd20790,32'd20844,32'd20898,32'd20952,32'd21006,32'd21060,32'd21114,32'd21168,32'd21222,32'd21276,32'd21330,32'd21384,32'd21438,32'd21492,32'd21546 };matrix[55]='{32'd0,32'd55,32'd110,32'd165,32'd220,32'd275,32'd330,32'd385,32'd440,32'd495,32'd550,32'd605,32'd660,32'd715,32'd770,32'd825,32'd880,32'd935,32'd990,32'd1045,32'd1100,32'd1155,32'd1210,32'd1265,32'd1320,32'd1375,32'd1430,32'd1485,32'd1540,32'd1595,32'd1650,32'd1705,32'd1760,32'd1815,32'd1870,32'd1925,32'd1980,32'd2035,32'd2090,32'd2145,32'd2200,32'd2255,32'd2310,32'd2365,32'd2420,32'd2475,32'd2530,32'd2585,32'd2640,32'd2695,32'd2750,32'd2805,32'd2860,32'd2915,32'd2970,32'd3025,32'd3080,32'd3135,32'd3190,32'd3245,32'd3300,32'd3355,32'd3410,32'd3465,32'd3520,32'd3575,32'd3630,32'd3685,32'd3740,32'd3795,32'd3850,32'd3905,32'd3960,32'd4015,32'd4070,32'd4125,32'd4180,32'd4235,32'd4290,32'd4345,32'd4400,32'd4455,32'd4510,32'd4565,32'd4620,32'd4675,32'd4730,32'd4785,32'd4840,32'd4895,32'd4950,32'd5005,32'd5060,32'd5115,32'd5170,32'd5225,32'd5280,32'd5335,32'd5390,32'd5445,32'd5500,32'd5555,32'd5610,32'd5665,32'd5720,32'd5775,32'd5830,32'd5885,32'd5940,32'd5995,32'd6050,32'd6105,32'd6160,32'd6215,32'd6270,32'd6325,32'd6380,32'd6435,32'd6490,32'd6545,32'd6600,32'd6655,32'd6710,32'd6765,32'd6820,32'd6875,32'd6930,32'd6985,32'd7040,32'd7095,32'd7150,32'd7205,32'd7260,32'd7315,32'd7370,32'd7425,32'd7480,32'd7535,32'd7590,32'd7645,32'd7700,32'd7755,32'd7810,32'd7865,32'd7920,32'd7975,32'd8030,32'd8085,32'd8140,32'd8195,32'd8250,32'd8305,32'd8360,32'd8415,32'd8470,32'd8525,32'd8580,32'd8635,32'd8690,32'd8745,32'd8800,32'd8855,32'd8910,32'd8965,32'd9020,32'd9075,32'd9130,32'd9185,32'd9240,32'd9295,32'd9350,32'd9405,32'd9460,32'd9515,32'd9570,32'd9625,32'd9680,32'd9735,32'd9790,32'd9845,32'd9900,32'd9955,32'd10010,32'd10065,32'd10120,32'd10175,32'd10230,32'd10285,32'd10340,32'd10395,32'd10450,32'd10505,32'd10560,32'd10615,32'd10670,32'd10725,32'd10780,32'd10835,32'd10890,32'd10945,32'd11000,32'd11055,32'd11110,32'd11165,32'd11220,32'd11275,32'd11330,32'd11385,32'd11440,32'd11495,32'd11550,32'd11605,32'd11660,32'd11715,32'd11770,32'd11825,32'd11880,32'd11935,32'd11990,32'd12045,32'd12100,32'd12155,32'd12210,32'd12265,32'd12320,32'd12375,32'd12430,32'd12485,32'd12540,32'd12595,32'd12650,32'd12705,32'd12760,32'd12815,32'd12870,32'd12925,32'd12980,32'd13035,32'd13090,32'd13145,32'd13200,32'd13255,32'd13310,32'd13365,32'd13420,32'd13475,32'd13530,32'd13585,32'd13640,32'd13695,32'd13750,32'd13805,32'd13860,32'd13915,32'd13970,32'd14025,32'd14080,32'd14135,32'd14190,32'd14245,32'd14300,32'd14355,32'd14410,32'd14465,32'd14520,32'd14575,32'd14630,32'd14685,32'd14740,32'd14795,32'd14850,32'd14905,32'd14960,32'd15015,32'd15070,32'd15125,32'd15180,32'd15235,32'd15290,32'd15345,32'd15400,32'd15455,32'd15510,32'd15565,32'd15620,32'd15675,32'd15730,32'd15785,32'd15840,32'd15895,32'd15950,32'd16005,32'd16060,32'd16115,32'd16170,32'd16225,32'd16280,32'd16335,32'd16390,32'd16445,32'd16500,32'd16555,32'd16610,32'd16665,32'd16720,32'd16775,32'd16830,32'd16885,32'd16940,32'd16995,32'd17050,32'd17105,32'd17160,32'd17215,32'd17270,32'd17325,32'd17380,32'd17435,32'd17490,32'd17545,32'd17600,32'd17655,32'd17710,32'd17765,32'd17820,32'd17875,32'd17930,32'd17985,32'd18040,32'd18095,32'd18150,32'd18205,32'd18260,32'd18315,32'd18370,32'd18425,32'd18480,32'd18535,32'd18590,32'd18645,32'd18700,32'd18755,32'd18810,32'd18865,32'd18920,32'd18975,32'd19030,32'd19085,32'd19140,32'd19195,32'd19250,32'd19305,32'd19360,32'd19415,32'd19470,32'd19525,32'd19580,32'd19635,32'd19690,32'd19745,32'd19800,32'd19855,32'd19910,32'd19965,32'd20020,32'd20075,32'd20130,32'd20185,32'd20240,32'd20295,32'd20350,32'd20405,32'd20460,32'd20515,32'd20570,32'd20625,32'd20680,32'd20735,32'd20790,32'd20845,32'd20900,32'd20955,32'd21010,32'd21065,32'd21120,32'd21175,32'd21230,32'd21285,32'd21340,32'd21395,32'd21450,32'd21505,32'd21560,32'd21615,32'd21670,32'd21725,32'd21780,32'd21835,32'd21890,32'd21945 };matrix[56]='{32'd0,32'd56,32'd112,32'd168,32'd224,32'd280,32'd336,32'd392,32'd448,32'd504,32'd560,32'd616,32'd672,32'd728,32'd784,32'd840,32'd896,32'd952,32'd1008,32'd1064,32'd1120,32'd1176,32'd1232,32'd1288,32'd1344,32'd1400,32'd1456,32'd1512,32'd1568,32'd1624,32'd1680,32'd1736,32'd1792,32'd1848,32'd1904,32'd1960,32'd2016,32'd2072,32'd2128,32'd2184,32'd2240,32'd2296,32'd2352,32'd2408,32'd2464,32'd2520,32'd2576,32'd2632,32'd2688,32'd2744,32'd2800,32'd2856,32'd2912,32'd2968,32'd3024,32'd3080,32'd3136,32'd3192,32'd3248,32'd3304,32'd3360,32'd3416,32'd3472,32'd3528,32'd3584,32'd3640,32'd3696,32'd3752,32'd3808,32'd3864,32'd3920,32'd3976,32'd4032,32'd4088,32'd4144,32'd4200,32'd4256,32'd4312,32'd4368,32'd4424,32'd4480,32'd4536,32'd4592,32'd4648,32'd4704,32'd4760,32'd4816,32'd4872,32'd4928,32'd4984,32'd5040,32'd5096,32'd5152,32'd5208,32'd5264,32'd5320,32'd5376,32'd5432,32'd5488,32'd5544,32'd5600,32'd5656,32'd5712,32'd5768,32'd5824,32'd5880,32'd5936,32'd5992,32'd6048,32'd6104,32'd6160,32'd6216,32'd6272,32'd6328,32'd6384,32'd6440,32'd6496,32'd6552,32'd6608,32'd6664,32'd6720,32'd6776,32'd6832,32'd6888,32'd6944,32'd7000,32'd7056,32'd7112,32'd7168,32'd7224,32'd7280,32'd7336,32'd7392,32'd7448,32'd7504,32'd7560,32'd7616,32'd7672,32'd7728,32'd7784,32'd7840,32'd7896,32'd7952,32'd8008,32'd8064,32'd8120,32'd8176,32'd8232,32'd8288,32'd8344,32'd8400,32'd8456,32'd8512,32'd8568,32'd8624,32'd8680,32'd8736,32'd8792,32'd8848,32'd8904,32'd8960,32'd9016,32'd9072,32'd9128,32'd9184,32'd9240,32'd9296,32'd9352,32'd9408,32'd9464,32'd9520,32'd9576,32'd9632,32'd9688,32'd9744,32'd9800,32'd9856,32'd9912,32'd9968,32'd10024,32'd10080,32'd10136,32'd10192,32'd10248,32'd10304,32'd10360,32'd10416,32'd10472,32'd10528,32'd10584,32'd10640,32'd10696,32'd10752,32'd10808,32'd10864,32'd10920,32'd10976,32'd11032,32'd11088,32'd11144,32'd11200,32'd11256,32'd11312,32'd11368,32'd11424,32'd11480,32'd11536,32'd11592,32'd11648,32'd11704,32'd11760,32'd11816,32'd11872,32'd11928,32'd11984,32'd12040,32'd12096,32'd12152,32'd12208,32'd12264,32'd12320,32'd12376,32'd12432,32'd12488,32'd12544,32'd12600,32'd12656,32'd12712,32'd12768,32'd12824,32'd12880,32'd12936,32'd12992,32'd13048,32'd13104,32'd13160,32'd13216,32'd13272,32'd13328,32'd13384,32'd13440,32'd13496,32'd13552,32'd13608,32'd13664,32'd13720,32'd13776,32'd13832,32'd13888,32'd13944,32'd14000,32'd14056,32'd14112,32'd14168,32'd14224,32'd14280,32'd14336,32'd14392,32'd14448,32'd14504,32'd14560,32'd14616,32'd14672,32'd14728,32'd14784,32'd14840,32'd14896,32'd14952,32'd15008,32'd15064,32'd15120,32'd15176,32'd15232,32'd15288,32'd15344,32'd15400,32'd15456,32'd15512,32'd15568,32'd15624,32'd15680,32'd15736,32'd15792,32'd15848,32'd15904,32'd15960,32'd16016,32'd16072,32'd16128,32'd16184,32'd16240,32'd16296,32'd16352,32'd16408,32'd16464,32'd16520,32'd16576,32'd16632,32'd16688,32'd16744,32'd16800,32'd16856,32'd16912,32'd16968,32'd17024,32'd17080,32'd17136,32'd17192,32'd17248,32'd17304,32'd17360,32'd17416,32'd17472,32'd17528,32'd17584,32'd17640,32'd17696,32'd17752,32'd17808,32'd17864,32'd17920,32'd17976,32'd18032,32'd18088,32'd18144,32'd18200,32'd18256,32'd18312,32'd18368,32'd18424,32'd18480,32'd18536,32'd18592,32'd18648,32'd18704,32'd18760,32'd18816,32'd18872,32'd18928,32'd18984,32'd19040,32'd19096,32'd19152,32'd19208,32'd19264,32'd19320,32'd19376,32'd19432,32'd19488,32'd19544,32'd19600,32'd19656,32'd19712,32'd19768,32'd19824,32'd19880,32'd19936,32'd19992,32'd20048,32'd20104,32'd20160,32'd20216,32'd20272,32'd20328,32'd20384,32'd20440,32'd20496,32'd20552,32'd20608,32'd20664,32'd20720,32'd20776,32'd20832,32'd20888,32'd20944,32'd21000,32'd21056,32'd21112,32'd21168,32'd21224,32'd21280,32'd21336,32'd21392,32'd21448,32'd21504,32'd21560,32'd21616,32'd21672,32'd21728,32'd21784,32'd21840,32'd21896,32'd21952,32'd22008,32'd22064,32'd22120,32'd22176,32'd22232,32'd22288,32'd22344 };matrix[57]='{32'd0,32'd57,32'd114,32'd171,32'd228,32'd285,32'd342,32'd399,32'd456,32'd513,32'd570,32'd627,32'd684,32'd741,32'd798,32'd855,32'd912,32'd969,32'd1026,32'd1083,32'd1140,32'd1197,32'd1254,32'd1311,32'd1368,32'd1425,32'd1482,32'd1539,32'd1596,32'd1653,32'd1710,32'd1767,32'd1824,32'd1881,32'd1938,32'd1995,32'd2052,32'd2109,32'd2166,32'd2223,32'd2280,32'd2337,32'd2394,32'd2451,32'd2508,32'd2565,32'd2622,32'd2679,32'd2736,32'd2793,32'd2850,32'd2907,32'd2964,32'd3021,32'd3078,32'd3135,32'd3192,32'd3249,32'd3306,32'd3363,32'd3420,32'd3477,32'd3534,32'd3591,32'd3648,32'd3705,32'd3762,32'd3819,32'd3876,32'd3933,32'd3990,32'd4047,32'd4104,32'd4161,32'd4218,32'd4275,32'd4332,32'd4389,32'd4446,32'd4503,32'd4560,32'd4617,32'd4674,32'd4731,32'd4788,32'd4845,32'd4902,32'd4959,32'd5016,32'd5073,32'd5130,32'd5187,32'd5244,32'd5301,32'd5358,32'd5415,32'd5472,32'd5529,32'd5586,32'd5643,32'd5700,32'd5757,32'd5814,32'd5871,32'd5928,32'd5985,32'd6042,32'd6099,32'd6156,32'd6213,32'd6270,32'd6327,32'd6384,32'd6441,32'd6498,32'd6555,32'd6612,32'd6669,32'd6726,32'd6783,32'd6840,32'd6897,32'd6954,32'd7011,32'd7068,32'd7125,32'd7182,32'd7239,32'd7296,32'd7353,32'd7410,32'd7467,32'd7524,32'd7581,32'd7638,32'd7695,32'd7752,32'd7809,32'd7866,32'd7923,32'd7980,32'd8037,32'd8094,32'd8151,32'd8208,32'd8265,32'd8322,32'd8379,32'd8436,32'd8493,32'd8550,32'd8607,32'd8664,32'd8721,32'd8778,32'd8835,32'd8892,32'd8949,32'd9006,32'd9063,32'd9120,32'd9177,32'd9234,32'd9291,32'd9348,32'd9405,32'd9462,32'd9519,32'd9576,32'd9633,32'd9690,32'd9747,32'd9804,32'd9861,32'd9918,32'd9975,32'd10032,32'd10089,32'd10146,32'd10203,32'd10260,32'd10317,32'd10374,32'd10431,32'd10488,32'd10545,32'd10602,32'd10659,32'd10716,32'd10773,32'd10830,32'd10887,32'd10944,32'd11001,32'd11058,32'd11115,32'd11172,32'd11229,32'd11286,32'd11343,32'd11400,32'd11457,32'd11514,32'd11571,32'd11628,32'd11685,32'd11742,32'd11799,32'd11856,32'd11913,32'd11970,32'd12027,32'd12084,32'd12141,32'd12198,32'd12255,32'd12312,32'd12369,32'd12426,32'd12483,32'd12540,32'd12597,32'd12654,32'd12711,32'd12768,32'd12825,32'd12882,32'd12939,32'd12996,32'd13053,32'd13110,32'd13167,32'd13224,32'd13281,32'd13338,32'd13395,32'd13452,32'd13509,32'd13566,32'd13623,32'd13680,32'd13737,32'd13794,32'd13851,32'd13908,32'd13965,32'd14022,32'd14079,32'd14136,32'd14193,32'd14250,32'd14307,32'd14364,32'd14421,32'd14478,32'd14535,32'd14592,32'd14649,32'd14706,32'd14763,32'd14820,32'd14877,32'd14934,32'd14991,32'd15048,32'd15105,32'd15162,32'd15219,32'd15276,32'd15333,32'd15390,32'd15447,32'd15504,32'd15561,32'd15618,32'd15675,32'd15732,32'd15789,32'd15846,32'd15903,32'd15960,32'd16017,32'd16074,32'd16131,32'd16188,32'd16245,32'd16302,32'd16359,32'd16416,32'd16473,32'd16530,32'd16587,32'd16644,32'd16701,32'd16758,32'd16815,32'd16872,32'd16929,32'd16986,32'd17043,32'd17100,32'd17157,32'd17214,32'd17271,32'd17328,32'd17385,32'd17442,32'd17499,32'd17556,32'd17613,32'd17670,32'd17727,32'd17784,32'd17841,32'd17898,32'd17955,32'd18012,32'd18069,32'd18126,32'd18183,32'd18240,32'd18297,32'd18354,32'd18411,32'd18468,32'd18525,32'd18582,32'd18639,32'd18696,32'd18753,32'd18810,32'd18867,32'd18924,32'd18981,32'd19038,32'd19095,32'd19152,32'd19209,32'd19266,32'd19323,32'd19380,32'd19437,32'd19494,32'd19551,32'd19608,32'd19665,32'd19722,32'd19779,32'd19836,32'd19893,32'd19950,32'd20007,32'd20064,32'd20121,32'd20178,32'd20235,32'd20292,32'd20349,32'd20406,32'd20463,32'd20520,32'd20577,32'd20634,32'd20691,32'd20748,32'd20805,32'd20862,32'd20919,32'd20976,32'd21033,32'd21090,32'd21147,32'd21204,32'd21261,32'd21318,32'd21375,32'd21432,32'd21489,32'd21546,32'd21603,32'd21660,32'd21717,32'd21774,32'd21831,32'd21888,32'd21945,32'd22002,32'd22059,32'd22116,32'd22173,32'd22230,32'd22287,32'd22344,32'd22401,32'd22458,32'd22515,32'd22572,32'd22629,32'd22686,32'd22743 };matrix[58]='{32'd0,32'd58,32'd116,32'd174,32'd232,32'd290,32'd348,32'd406,32'd464,32'd522,32'd580,32'd638,32'd696,32'd754,32'd812,32'd870,32'd928,32'd986,32'd1044,32'd1102,32'd1160,32'd1218,32'd1276,32'd1334,32'd1392,32'd1450,32'd1508,32'd1566,32'd1624,32'd1682,32'd1740,32'd1798,32'd1856,32'd1914,32'd1972,32'd2030,32'd2088,32'd2146,32'd2204,32'd2262,32'd2320,32'd2378,32'd2436,32'd2494,32'd2552,32'd2610,32'd2668,32'd2726,32'd2784,32'd2842,32'd2900,32'd2958,32'd3016,32'd3074,32'd3132,32'd3190,32'd3248,32'd3306,32'd3364,32'd3422,32'd3480,32'd3538,32'd3596,32'd3654,32'd3712,32'd3770,32'd3828,32'd3886,32'd3944,32'd4002,32'd4060,32'd4118,32'd4176,32'd4234,32'd4292,32'd4350,32'd4408,32'd4466,32'd4524,32'd4582,32'd4640,32'd4698,32'd4756,32'd4814,32'd4872,32'd4930,32'd4988,32'd5046,32'd5104,32'd5162,32'd5220,32'd5278,32'd5336,32'd5394,32'd5452,32'd5510,32'd5568,32'd5626,32'd5684,32'd5742,32'd5800,32'd5858,32'd5916,32'd5974,32'd6032,32'd6090,32'd6148,32'd6206,32'd6264,32'd6322,32'd6380,32'd6438,32'd6496,32'd6554,32'd6612,32'd6670,32'd6728,32'd6786,32'd6844,32'd6902,32'd6960,32'd7018,32'd7076,32'd7134,32'd7192,32'd7250,32'd7308,32'd7366,32'd7424,32'd7482,32'd7540,32'd7598,32'd7656,32'd7714,32'd7772,32'd7830,32'd7888,32'd7946,32'd8004,32'd8062,32'd8120,32'd8178,32'd8236,32'd8294,32'd8352,32'd8410,32'd8468,32'd8526,32'd8584,32'd8642,32'd8700,32'd8758,32'd8816,32'd8874,32'd8932,32'd8990,32'd9048,32'd9106,32'd9164,32'd9222,32'd9280,32'd9338,32'd9396,32'd9454,32'd9512,32'd9570,32'd9628,32'd9686,32'd9744,32'd9802,32'd9860,32'd9918,32'd9976,32'd10034,32'd10092,32'd10150,32'd10208,32'd10266,32'd10324,32'd10382,32'd10440,32'd10498,32'd10556,32'd10614,32'd10672,32'd10730,32'd10788,32'd10846,32'd10904,32'd10962,32'd11020,32'd11078,32'd11136,32'd11194,32'd11252,32'd11310,32'd11368,32'd11426,32'd11484,32'd11542,32'd11600,32'd11658,32'd11716,32'd11774,32'd11832,32'd11890,32'd11948,32'd12006,32'd12064,32'd12122,32'd12180,32'd12238,32'd12296,32'd12354,32'd12412,32'd12470,32'd12528,32'd12586,32'd12644,32'd12702,32'd12760,32'd12818,32'd12876,32'd12934,32'd12992,32'd13050,32'd13108,32'd13166,32'd13224,32'd13282,32'd13340,32'd13398,32'd13456,32'd13514,32'd13572,32'd13630,32'd13688,32'd13746,32'd13804,32'd13862,32'd13920,32'd13978,32'd14036,32'd14094,32'd14152,32'd14210,32'd14268,32'd14326,32'd14384,32'd14442,32'd14500,32'd14558,32'd14616,32'd14674,32'd14732,32'd14790,32'd14848,32'd14906,32'd14964,32'd15022,32'd15080,32'd15138,32'd15196,32'd15254,32'd15312,32'd15370,32'd15428,32'd15486,32'd15544,32'd15602,32'd15660,32'd15718,32'd15776,32'd15834,32'd15892,32'd15950,32'd16008,32'd16066,32'd16124,32'd16182,32'd16240,32'd16298,32'd16356,32'd16414,32'd16472,32'd16530,32'd16588,32'd16646,32'd16704,32'd16762,32'd16820,32'd16878,32'd16936,32'd16994,32'd17052,32'd17110,32'd17168,32'd17226,32'd17284,32'd17342,32'd17400,32'd17458,32'd17516,32'd17574,32'd17632,32'd17690,32'd17748,32'd17806,32'd17864,32'd17922,32'd17980,32'd18038,32'd18096,32'd18154,32'd18212,32'd18270,32'd18328,32'd18386,32'd18444,32'd18502,32'd18560,32'd18618,32'd18676,32'd18734,32'd18792,32'd18850,32'd18908,32'd18966,32'd19024,32'd19082,32'd19140,32'd19198,32'd19256,32'd19314,32'd19372,32'd19430,32'd19488,32'd19546,32'd19604,32'd19662,32'd19720,32'd19778,32'd19836,32'd19894,32'd19952,32'd20010,32'd20068,32'd20126,32'd20184,32'd20242,32'd20300,32'd20358,32'd20416,32'd20474,32'd20532,32'd20590,32'd20648,32'd20706,32'd20764,32'd20822,32'd20880,32'd20938,32'd20996,32'd21054,32'd21112,32'd21170,32'd21228,32'd21286,32'd21344,32'd21402,32'd21460,32'd21518,32'd21576,32'd21634,32'd21692,32'd21750,32'd21808,32'd21866,32'd21924,32'd21982,32'd22040,32'd22098,32'd22156,32'd22214,32'd22272,32'd22330,32'd22388,32'd22446,32'd22504,32'd22562,32'd22620,32'd22678,32'd22736,32'd22794,32'd22852,32'd22910,32'd22968,32'd23026,32'd23084,32'd23142 };matrix[59]='{32'd0,32'd59,32'd118,32'd177,32'd236,32'd295,32'd354,32'd413,32'd472,32'd531,32'd590,32'd649,32'd708,32'd767,32'd826,32'd885,32'd944,32'd1003,32'd1062,32'd1121,32'd1180,32'd1239,32'd1298,32'd1357,32'd1416,32'd1475,32'd1534,32'd1593,32'd1652,32'd1711,32'd1770,32'd1829,32'd1888,32'd1947,32'd2006,32'd2065,32'd2124,32'd2183,32'd2242,32'd2301,32'd2360,32'd2419,32'd2478,32'd2537,32'd2596,32'd2655,32'd2714,32'd2773,32'd2832,32'd2891,32'd2950,32'd3009,32'd3068,32'd3127,32'd3186,32'd3245,32'd3304,32'd3363,32'd3422,32'd3481,32'd3540,32'd3599,32'd3658,32'd3717,32'd3776,32'd3835,32'd3894,32'd3953,32'd4012,32'd4071,32'd4130,32'd4189,32'd4248,32'd4307,32'd4366,32'd4425,32'd4484,32'd4543,32'd4602,32'd4661,32'd4720,32'd4779,32'd4838,32'd4897,32'd4956,32'd5015,32'd5074,32'd5133,32'd5192,32'd5251,32'd5310,32'd5369,32'd5428,32'd5487,32'd5546,32'd5605,32'd5664,32'd5723,32'd5782,32'd5841,32'd5900,32'd5959,32'd6018,32'd6077,32'd6136,32'd6195,32'd6254,32'd6313,32'd6372,32'd6431,32'd6490,32'd6549,32'd6608,32'd6667,32'd6726,32'd6785,32'd6844,32'd6903,32'd6962,32'd7021,32'd7080,32'd7139,32'd7198,32'd7257,32'd7316,32'd7375,32'd7434,32'd7493,32'd7552,32'd7611,32'd7670,32'd7729,32'd7788,32'd7847,32'd7906,32'd7965,32'd8024,32'd8083,32'd8142,32'd8201,32'd8260,32'd8319,32'd8378,32'd8437,32'd8496,32'd8555,32'd8614,32'd8673,32'd8732,32'd8791,32'd8850,32'd8909,32'd8968,32'd9027,32'd9086,32'd9145,32'd9204,32'd9263,32'd9322,32'd9381,32'd9440,32'd9499,32'd9558,32'd9617,32'd9676,32'd9735,32'd9794,32'd9853,32'd9912,32'd9971,32'd10030,32'd10089,32'd10148,32'd10207,32'd10266,32'd10325,32'd10384,32'd10443,32'd10502,32'd10561,32'd10620,32'd10679,32'd10738,32'd10797,32'd10856,32'd10915,32'd10974,32'd11033,32'd11092,32'd11151,32'd11210,32'd11269,32'd11328,32'd11387,32'd11446,32'd11505,32'd11564,32'd11623,32'd11682,32'd11741,32'd11800,32'd11859,32'd11918,32'd11977,32'd12036,32'd12095,32'd12154,32'd12213,32'd12272,32'd12331,32'd12390,32'd12449,32'd12508,32'd12567,32'd12626,32'd12685,32'd12744,32'd12803,32'd12862,32'd12921,32'd12980,32'd13039,32'd13098,32'd13157,32'd13216,32'd13275,32'd13334,32'd13393,32'd13452,32'd13511,32'd13570,32'd13629,32'd13688,32'd13747,32'd13806,32'd13865,32'd13924,32'd13983,32'd14042,32'd14101,32'd14160,32'd14219,32'd14278,32'd14337,32'd14396,32'd14455,32'd14514,32'd14573,32'd14632,32'd14691,32'd14750,32'd14809,32'd14868,32'd14927,32'd14986,32'd15045,32'd15104,32'd15163,32'd15222,32'd15281,32'd15340,32'd15399,32'd15458,32'd15517,32'd15576,32'd15635,32'd15694,32'd15753,32'd15812,32'd15871,32'd15930,32'd15989,32'd16048,32'd16107,32'd16166,32'd16225,32'd16284,32'd16343,32'd16402,32'd16461,32'd16520,32'd16579,32'd16638,32'd16697,32'd16756,32'd16815,32'd16874,32'd16933,32'd16992,32'd17051,32'd17110,32'd17169,32'd17228,32'd17287,32'd17346,32'd17405,32'd17464,32'd17523,32'd17582,32'd17641,32'd17700,32'd17759,32'd17818,32'd17877,32'd17936,32'd17995,32'd18054,32'd18113,32'd18172,32'd18231,32'd18290,32'd18349,32'd18408,32'd18467,32'd18526,32'd18585,32'd18644,32'd18703,32'd18762,32'd18821,32'd18880,32'd18939,32'd18998,32'd19057,32'd19116,32'd19175,32'd19234,32'd19293,32'd19352,32'd19411,32'd19470,32'd19529,32'd19588,32'd19647,32'd19706,32'd19765,32'd19824,32'd19883,32'd19942,32'd20001,32'd20060,32'd20119,32'd20178,32'd20237,32'd20296,32'd20355,32'd20414,32'd20473,32'd20532,32'd20591,32'd20650,32'd20709,32'd20768,32'd20827,32'd20886,32'd20945,32'd21004,32'd21063,32'd21122,32'd21181,32'd21240,32'd21299,32'd21358,32'd21417,32'd21476,32'd21535,32'd21594,32'd21653,32'd21712,32'd21771,32'd21830,32'd21889,32'd21948,32'd22007,32'd22066,32'd22125,32'd22184,32'd22243,32'd22302,32'd22361,32'd22420,32'd22479,32'd22538,32'd22597,32'd22656,32'd22715,32'd22774,32'd22833,32'd22892,32'd22951,32'd23010,32'd23069,32'd23128,32'd23187,32'd23246,32'd23305,32'd23364,32'd23423,32'd23482,32'd23541 };matrix[60]='{32'd0,32'd60,32'd120,32'd180,32'd240,32'd300,32'd360,32'd420,32'd480,32'd540,32'd600,32'd660,32'd720,32'd780,32'd840,32'd900,32'd960,32'd1020,32'd1080,32'd1140,32'd1200,32'd1260,32'd1320,32'd1380,32'd1440,32'd1500,32'd1560,32'd1620,32'd1680,32'd1740,32'd1800,32'd1860,32'd1920,32'd1980,32'd2040,32'd2100,32'd2160,32'd2220,32'd2280,32'd2340,32'd2400,32'd2460,32'd2520,32'd2580,32'd2640,32'd2700,32'd2760,32'd2820,32'd2880,32'd2940,32'd3000,32'd3060,32'd3120,32'd3180,32'd3240,32'd3300,32'd3360,32'd3420,32'd3480,32'd3540,32'd3600,32'd3660,32'd3720,32'd3780,32'd3840,32'd3900,32'd3960,32'd4020,32'd4080,32'd4140,32'd4200,32'd4260,32'd4320,32'd4380,32'd4440,32'd4500,32'd4560,32'd4620,32'd4680,32'd4740,32'd4800,32'd4860,32'd4920,32'd4980,32'd5040,32'd5100,32'd5160,32'd5220,32'd5280,32'd5340,32'd5400,32'd5460,32'd5520,32'd5580,32'd5640,32'd5700,32'd5760,32'd5820,32'd5880,32'd5940,32'd6000,32'd6060,32'd6120,32'd6180,32'd6240,32'd6300,32'd6360,32'd6420,32'd6480,32'd6540,32'd6600,32'd6660,32'd6720,32'd6780,32'd6840,32'd6900,32'd6960,32'd7020,32'd7080,32'd7140,32'd7200,32'd7260,32'd7320,32'd7380,32'd7440,32'd7500,32'd7560,32'd7620,32'd7680,32'd7740,32'd7800,32'd7860,32'd7920,32'd7980,32'd8040,32'd8100,32'd8160,32'd8220,32'd8280,32'd8340,32'd8400,32'd8460,32'd8520,32'd8580,32'd8640,32'd8700,32'd8760,32'd8820,32'd8880,32'd8940,32'd9000,32'd9060,32'd9120,32'd9180,32'd9240,32'd9300,32'd9360,32'd9420,32'd9480,32'd9540,32'd9600,32'd9660,32'd9720,32'd9780,32'd9840,32'd9900,32'd9960,32'd10020,32'd10080,32'd10140,32'd10200,32'd10260,32'd10320,32'd10380,32'd10440,32'd10500,32'd10560,32'd10620,32'd10680,32'd10740,32'd10800,32'd10860,32'd10920,32'd10980,32'd11040,32'd11100,32'd11160,32'd11220,32'd11280,32'd11340,32'd11400,32'd11460,32'd11520,32'd11580,32'd11640,32'd11700,32'd11760,32'd11820,32'd11880,32'd11940,32'd12000,32'd12060,32'd12120,32'd12180,32'd12240,32'd12300,32'd12360,32'd12420,32'd12480,32'd12540,32'd12600,32'd12660,32'd12720,32'd12780,32'd12840,32'd12900,32'd12960,32'd13020,32'd13080,32'd13140,32'd13200,32'd13260,32'd13320,32'd13380,32'd13440,32'd13500,32'd13560,32'd13620,32'd13680,32'd13740,32'd13800,32'd13860,32'd13920,32'd13980,32'd14040,32'd14100,32'd14160,32'd14220,32'd14280,32'd14340,32'd14400,32'd14460,32'd14520,32'd14580,32'd14640,32'd14700,32'd14760,32'd14820,32'd14880,32'd14940,32'd15000,32'd15060,32'd15120,32'd15180,32'd15240,32'd15300,32'd15360,32'd15420,32'd15480,32'd15540,32'd15600,32'd15660,32'd15720,32'd15780,32'd15840,32'd15900,32'd15960,32'd16020,32'd16080,32'd16140,32'd16200,32'd16260,32'd16320,32'd16380,32'd16440,32'd16500,32'd16560,32'd16620,32'd16680,32'd16740,32'd16800,32'd16860,32'd16920,32'd16980,32'd17040,32'd17100,32'd17160,32'd17220,32'd17280,32'd17340,32'd17400,32'd17460,32'd17520,32'd17580,32'd17640,32'd17700,32'd17760,32'd17820,32'd17880,32'd17940,32'd18000,32'd18060,32'd18120,32'd18180,32'd18240,32'd18300,32'd18360,32'd18420,32'd18480,32'd18540,32'd18600,32'd18660,32'd18720,32'd18780,32'd18840,32'd18900,32'd18960,32'd19020,32'd19080,32'd19140,32'd19200,32'd19260,32'd19320,32'd19380,32'd19440,32'd19500,32'd19560,32'd19620,32'd19680,32'd19740,32'd19800,32'd19860,32'd19920,32'd19980,32'd20040,32'd20100,32'd20160,32'd20220,32'd20280,32'd20340,32'd20400,32'd20460,32'd20520,32'd20580,32'd20640,32'd20700,32'd20760,32'd20820,32'd20880,32'd20940,32'd21000,32'd21060,32'd21120,32'd21180,32'd21240,32'd21300,32'd21360,32'd21420,32'd21480,32'd21540,32'd21600,32'd21660,32'd21720,32'd21780,32'd21840,32'd21900,32'd21960,32'd22020,32'd22080,32'd22140,32'd22200,32'd22260,32'd22320,32'd22380,32'd22440,32'd22500,32'd22560,32'd22620,32'd22680,32'd22740,32'd22800,32'd22860,32'd22920,32'd22980,32'd23040,32'd23100,32'd23160,32'd23220,32'd23280,32'd23340,32'd23400,32'd23460,32'd23520,32'd23580,32'd23640,32'd23700,32'd23760,32'd23820,32'd23880,32'd23940 };matrix[61]='{32'd0,32'd61,32'd122,32'd183,32'd244,32'd305,32'd366,32'd427,32'd488,32'd549,32'd610,32'd671,32'd732,32'd793,32'd854,32'd915,32'd976,32'd1037,32'd1098,32'd1159,32'd1220,32'd1281,32'd1342,32'd1403,32'd1464,32'd1525,32'd1586,32'd1647,32'd1708,32'd1769,32'd1830,32'd1891,32'd1952,32'd2013,32'd2074,32'd2135,32'd2196,32'd2257,32'd2318,32'd2379,32'd2440,32'd2501,32'd2562,32'd2623,32'd2684,32'd2745,32'd2806,32'd2867,32'd2928,32'd2989,32'd3050,32'd3111,32'd3172,32'd3233,32'd3294,32'd3355,32'd3416,32'd3477,32'd3538,32'd3599,32'd3660,32'd3721,32'd3782,32'd3843,32'd3904,32'd3965,32'd4026,32'd4087,32'd4148,32'd4209,32'd4270,32'd4331,32'd4392,32'd4453,32'd4514,32'd4575,32'd4636,32'd4697,32'd4758,32'd4819,32'd4880,32'd4941,32'd5002,32'd5063,32'd5124,32'd5185,32'd5246,32'd5307,32'd5368,32'd5429,32'd5490,32'd5551,32'd5612,32'd5673,32'd5734,32'd5795,32'd5856,32'd5917,32'd5978,32'd6039,32'd6100,32'd6161,32'd6222,32'd6283,32'd6344,32'd6405,32'd6466,32'd6527,32'd6588,32'd6649,32'd6710,32'd6771,32'd6832,32'd6893,32'd6954,32'd7015,32'd7076,32'd7137,32'd7198,32'd7259,32'd7320,32'd7381,32'd7442,32'd7503,32'd7564,32'd7625,32'd7686,32'd7747,32'd7808,32'd7869,32'd7930,32'd7991,32'd8052,32'd8113,32'd8174,32'd8235,32'd8296,32'd8357,32'd8418,32'd8479,32'd8540,32'd8601,32'd8662,32'd8723,32'd8784,32'd8845,32'd8906,32'd8967,32'd9028,32'd9089,32'd9150,32'd9211,32'd9272,32'd9333,32'd9394,32'd9455,32'd9516,32'd9577,32'd9638,32'd9699,32'd9760,32'd9821,32'd9882,32'd9943,32'd10004,32'd10065,32'd10126,32'd10187,32'd10248,32'd10309,32'd10370,32'd10431,32'd10492,32'd10553,32'd10614,32'd10675,32'd10736,32'd10797,32'd10858,32'd10919,32'd10980,32'd11041,32'd11102,32'd11163,32'd11224,32'd11285,32'd11346,32'd11407,32'd11468,32'd11529,32'd11590,32'd11651,32'd11712,32'd11773,32'd11834,32'd11895,32'd11956,32'd12017,32'd12078,32'd12139,32'd12200,32'd12261,32'd12322,32'd12383,32'd12444,32'd12505,32'd12566,32'd12627,32'd12688,32'd12749,32'd12810,32'd12871,32'd12932,32'd12993,32'd13054,32'd13115,32'd13176,32'd13237,32'd13298,32'd13359,32'd13420,32'd13481,32'd13542,32'd13603,32'd13664,32'd13725,32'd13786,32'd13847,32'd13908,32'd13969,32'd14030,32'd14091,32'd14152,32'd14213,32'd14274,32'd14335,32'd14396,32'd14457,32'd14518,32'd14579,32'd14640,32'd14701,32'd14762,32'd14823,32'd14884,32'd14945,32'd15006,32'd15067,32'd15128,32'd15189,32'd15250,32'd15311,32'd15372,32'd15433,32'd15494,32'd15555,32'd15616,32'd15677,32'd15738,32'd15799,32'd15860,32'd15921,32'd15982,32'd16043,32'd16104,32'd16165,32'd16226,32'd16287,32'd16348,32'd16409,32'd16470,32'd16531,32'd16592,32'd16653,32'd16714,32'd16775,32'd16836,32'd16897,32'd16958,32'd17019,32'd17080,32'd17141,32'd17202,32'd17263,32'd17324,32'd17385,32'd17446,32'd17507,32'd17568,32'd17629,32'd17690,32'd17751,32'd17812,32'd17873,32'd17934,32'd17995,32'd18056,32'd18117,32'd18178,32'd18239,32'd18300,32'd18361,32'd18422,32'd18483,32'd18544,32'd18605,32'd18666,32'd18727,32'd18788,32'd18849,32'd18910,32'd18971,32'd19032,32'd19093,32'd19154,32'd19215,32'd19276,32'd19337,32'd19398,32'd19459,32'd19520,32'd19581,32'd19642,32'd19703,32'd19764,32'd19825,32'd19886,32'd19947,32'd20008,32'd20069,32'd20130,32'd20191,32'd20252,32'd20313,32'd20374,32'd20435,32'd20496,32'd20557,32'd20618,32'd20679,32'd20740,32'd20801,32'd20862,32'd20923,32'd20984,32'd21045,32'd21106,32'd21167,32'd21228,32'd21289,32'd21350,32'd21411,32'd21472,32'd21533,32'd21594,32'd21655,32'd21716,32'd21777,32'd21838,32'd21899,32'd21960,32'd22021,32'd22082,32'd22143,32'd22204,32'd22265,32'd22326,32'd22387,32'd22448,32'd22509,32'd22570,32'd22631,32'd22692,32'd22753,32'd22814,32'd22875,32'd22936,32'd22997,32'd23058,32'd23119,32'd23180,32'd23241,32'd23302,32'd23363,32'd23424,32'd23485,32'd23546,32'd23607,32'd23668,32'd23729,32'd23790,32'd23851,32'd23912,32'd23973,32'd24034,32'd24095,32'd24156,32'd24217,32'd24278,32'd24339 };matrix[62]='{32'd0,32'd62,32'd124,32'd186,32'd248,32'd310,32'd372,32'd434,32'd496,32'd558,32'd620,32'd682,32'd744,32'd806,32'd868,32'd930,32'd992,32'd1054,32'd1116,32'd1178,32'd1240,32'd1302,32'd1364,32'd1426,32'd1488,32'd1550,32'd1612,32'd1674,32'd1736,32'd1798,32'd1860,32'd1922,32'd1984,32'd2046,32'd2108,32'd2170,32'd2232,32'd2294,32'd2356,32'd2418,32'd2480,32'd2542,32'd2604,32'd2666,32'd2728,32'd2790,32'd2852,32'd2914,32'd2976,32'd3038,32'd3100,32'd3162,32'd3224,32'd3286,32'd3348,32'd3410,32'd3472,32'd3534,32'd3596,32'd3658,32'd3720,32'd3782,32'd3844,32'd3906,32'd3968,32'd4030,32'd4092,32'd4154,32'd4216,32'd4278,32'd4340,32'd4402,32'd4464,32'd4526,32'd4588,32'd4650,32'd4712,32'd4774,32'd4836,32'd4898,32'd4960,32'd5022,32'd5084,32'd5146,32'd5208,32'd5270,32'd5332,32'd5394,32'd5456,32'd5518,32'd5580,32'd5642,32'd5704,32'd5766,32'd5828,32'd5890,32'd5952,32'd6014,32'd6076,32'd6138,32'd6200,32'd6262,32'd6324,32'd6386,32'd6448,32'd6510,32'd6572,32'd6634,32'd6696,32'd6758,32'd6820,32'd6882,32'd6944,32'd7006,32'd7068,32'd7130,32'd7192,32'd7254,32'd7316,32'd7378,32'd7440,32'd7502,32'd7564,32'd7626,32'd7688,32'd7750,32'd7812,32'd7874,32'd7936,32'd7998,32'd8060,32'd8122,32'd8184,32'd8246,32'd8308,32'd8370,32'd8432,32'd8494,32'd8556,32'd8618,32'd8680,32'd8742,32'd8804,32'd8866,32'd8928,32'd8990,32'd9052,32'd9114,32'd9176,32'd9238,32'd9300,32'd9362,32'd9424,32'd9486,32'd9548,32'd9610,32'd9672,32'd9734,32'd9796,32'd9858,32'd9920,32'd9982,32'd10044,32'd10106,32'd10168,32'd10230,32'd10292,32'd10354,32'd10416,32'd10478,32'd10540,32'd10602,32'd10664,32'd10726,32'd10788,32'd10850,32'd10912,32'd10974,32'd11036,32'd11098,32'd11160,32'd11222,32'd11284,32'd11346,32'd11408,32'd11470,32'd11532,32'd11594,32'd11656,32'd11718,32'd11780,32'd11842,32'd11904,32'd11966,32'd12028,32'd12090,32'd12152,32'd12214,32'd12276,32'd12338,32'd12400,32'd12462,32'd12524,32'd12586,32'd12648,32'd12710,32'd12772,32'd12834,32'd12896,32'd12958,32'd13020,32'd13082,32'd13144,32'd13206,32'd13268,32'd13330,32'd13392,32'd13454,32'd13516,32'd13578,32'd13640,32'd13702,32'd13764,32'd13826,32'd13888,32'd13950,32'd14012,32'd14074,32'd14136,32'd14198,32'd14260,32'd14322,32'd14384,32'd14446,32'd14508,32'd14570,32'd14632,32'd14694,32'd14756,32'd14818,32'd14880,32'd14942,32'd15004,32'd15066,32'd15128,32'd15190,32'd15252,32'd15314,32'd15376,32'd15438,32'd15500,32'd15562,32'd15624,32'd15686,32'd15748,32'd15810,32'd15872,32'd15934,32'd15996,32'd16058,32'd16120,32'd16182,32'd16244,32'd16306,32'd16368,32'd16430,32'd16492,32'd16554,32'd16616,32'd16678,32'd16740,32'd16802,32'd16864,32'd16926,32'd16988,32'd17050,32'd17112,32'd17174,32'd17236,32'd17298,32'd17360,32'd17422,32'd17484,32'd17546,32'd17608,32'd17670,32'd17732,32'd17794,32'd17856,32'd17918,32'd17980,32'd18042,32'd18104,32'd18166,32'd18228,32'd18290,32'd18352,32'd18414,32'd18476,32'd18538,32'd18600,32'd18662,32'd18724,32'd18786,32'd18848,32'd18910,32'd18972,32'd19034,32'd19096,32'd19158,32'd19220,32'd19282,32'd19344,32'd19406,32'd19468,32'd19530,32'd19592,32'd19654,32'd19716,32'd19778,32'd19840,32'd19902,32'd19964,32'd20026,32'd20088,32'd20150,32'd20212,32'd20274,32'd20336,32'd20398,32'd20460,32'd20522,32'd20584,32'd20646,32'd20708,32'd20770,32'd20832,32'd20894,32'd20956,32'd21018,32'd21080,32'd21142,32'd21204,32'd21266,32'd21328,32'd21390,32'd21452,32'd21514,32'd21576,32'd21638,32'd21700,32'd21762,32'd21824,32'd21886,32'd21948,32'd22010,32'd22072,32'd22134,32'd22196,32'd22258,32'd22320,32'd22382,32'd22444,32'd22506,32'd22568,32'd22630,32'd22692,32'd22754,32'd22816,32'd22878,32'd22940,32'd23002,32'd23064,32'd23126,32'd23188,32'd23250,32'd23312,32'd23374,32'd23436,32'd23498,32'd23560,32'd23622,32'd23684,32'd23746,32'd23808,32'd23870,32'd23932,32'd23994,32'd24056,32'd24118,32'd24180,32'd24242,32'd24304,32'd24366,32'd24428,32'd24490,32'd24552,32'd24614,32'd24676,32'd24738 };matrix[63]='{32'd0,32'd63,32'd126,32'd189,32'd252,32'd315,32'd378,32'd441,32'd504,32'd567,32'd630,32'd693,32'd756,32'd819,32'd882,32'd945,32'd1008,32'd1071,32'd1134,32'd1197,32'd1260,32'd1323,32'd1386,32'd1449,32'd1512,32'd1575,32'd1638,32'd1701,32'd1764,32'd1827,32'd1890,32'd1953,32'd2016,32'd2079,32'd2142,32'd2205,32'd2268,32'd2331,32'd2394,32'd2457,32'd2520,32'd2583,32'd2646,32'd2709,32'd2772,32'd2835,32'd2898,32'd2961,32'd3024,32'd3087,32'd3150,32'd3213,32'd3276,32'd3339,32'd3402,32'd3465,32'd3528,32'd3591,32'd3654,32'd3717,32'd3780,32'd3843,32'd3906,32'd3969,32'd4032,32'd4095,32'd4158,32'd4221,32'd4284,32'd4347,32'd4410,32'd4473,32'd4536,32'd4599,32'd4662,32'd4725,32'd4788,32'd4851,32'd4914,32'd4977,32'd5040,32'd5103,32'd5166,32'd5229,32'd5292,32'd5355,32'd5418,32'd5481,32'd5544,32'd5607,32'd5670,32'd5733,32'd5796,32'd5859,32'd5922,32'd5985,32'd6048,32'd6111,32'd6174,32'd6237,32'd6300,32'd6363,32'd6426,32'd6489,32'd6552,32'd6615,32'd6678,32'd6741,32'd6804,32'd6867,32'd6930,32'd6993,32'd7056,32'd7119,32'd7182,32'd7245,32'd7308,32'd7371,32'd7434,32'd7497,32'd7560,32'd7623,32'd7686,32'd7749,32'd7812,32'd7875,32'd7938,32'd8001,32'd8064,32'd8127,32'd8190,32'd8253,32'd8316,32'd8379,32'd8442,32'd8505,32'd8568,32'd8631,32'd8694,32'd8757,32'd8820,32'd8883,32'd8946,32'd9009,32'd9072,32'd9135,32'd9198,32'd9261,32'd9324,32'd9387,32'd9450,32'd9513,32'd9576,32'd9639,32'd9702,32'd9765,32'd9828,32'd9891,32'd9954,32'd10017,32'd10080,32'd10143,32'd10206,32'd10269,32'd10332,32'd10395,32'd10458,32'd10521,32'd10584,32'd10647,32'd10710,32'd10773,32'd10836,32'd10899,32'd10962,32'd11025,32'd11088,32'd11151,32'd11214,32'd11277,32'd11340,32'd11403,32'd11466,32'd11529,32'd11592,32'd11655,32'd11718,32'd11781,32'd11844,32'd11907,32'd11970,32'd12033,32'd12096,32'd12159,32'd12222,32'd12285,32'd12348,32'd12411,32'd12474,32'd12537,32'd12600,32'd12663,32'd12726,32'd12789,32'd12852,32'd12915,32'd12978,32'd13041,32'd13104,32'd13167,32'd13230,32'd13293,32'd13356,32'd13419,32'd13482,32'd13545,32'd13608,32'd13671,32'd13734,32'd13797,32'd13860,32'd13923,32'd13986,32'd14049,32'd14112,32'd14175,32'd14238,32'd14301,32'd14364,32'd14427,32'd14490,32'd14553,32'd14616,32'd14679,32'd14742,32'd14805,32'd14868,32'd14931,32'd14994,32'd15057,32'd15120,32'd15183,32'd15246,32'd15309,32'd15372,32'd15435,32'd15498,32'd15561,32'd15624,32'd15687,32'd15750,32'd15813,32'd15876,32'd15939,32'd16002,32'd16065,32'd16128,32'd16191,32'd16254,32'd16317,32'd16380,32'd16443,32'd16506,32'd16569,32'd16632,32'd16695,32'd16758,32'd16821,32'd16884,32'd16947,32'd17010,32'd17073,32'd17136,32'd17199,32'd17262,32'd17325,32'd17388,32'd17451,32'd17514,32'd17577,32'd17640,32'd17703,32'd17766,32'd17829,32'd17892,32'd17955,32'd18018,32'd18081,32'd18144,32'd18207,32'd18270,32'd18333,32'd18396,32'd18459,32'd18522,32'd18585,32'd18648,32'd18711,32'd18774,32'd18837,32'd18900,32'd18963,32'd19026,32'd19089,32'd19152,32'd19215,32'd19278,32'd19341,32'd19404,32'd19467,32'd19530,32'd19593,32'd19656,32'd19719,32'd19782,32'd19845,32'd19908,32'd19971,32'd20034,32'd20097,32'd20160,32'd20223,32'd20286,32'd20349,32'd20412,32'd20475,32'd20538,32'd20601,32'd20664,32'd20727,32'd20790,32'd20853,32'd20916,32'd20979,32'd21042,32'd21105,32'd21168,32'd21231,32'd21294,32'd21357,32'd21420,32'd21483,32'd21546,32'd21609,32'd21672,32'd21735,32'd21798,32'd21861,32'd21924,32'd21987,32'd22050,32'd22113,32'd22176,32'd22239,32'd22302,32'd22365,32'd22428,32'd22491,32'd22554,32'd22617,32'd22680,32'd22743,32'd22806,32'd22869,32'd22932,32'd22995,32'd23058,32'd23121,32'd23184,32'd23247,32'd23310,32'd23373,32'd23436,32'd23499,32'd23562,32'd23625,32'd23688,32'd23751,32'd23814,32'd23877,32'd23940,32'd24003,32'd24066,32'd24129,32'd24192,32'd24255,32'd24318,32'd24381,32'd24444,32'd24507,32'd24570,32'd24633,32'd24696,32'd24759,32'd24822,32'd24885,32'd24948,32'd25011,32'd25074,32'd25137 };matrix[64]='{32'd0,32'd64,32'd128,32'd192,32'd256,32'd320,32'd384,32'd448,32'd512,32'd576,32'd640,32'd704,32'd768,32'd832,32'd896,32'd960,32'd1024,32'd1088,32'd1152,32'd1216,32'd1280,32'd1344,32'd1408,32'd1472,32'd1536,32'd1600,32'd1664,32'd1728,32'd1792,32'd1856,32'd1920,32'd1984,32'd2048,32'd2112,32'd2176,32'd2240,32'd2304,32'd2368,32'd2432,32'd2496,32'd2560,32'd2624,32'd2688,32'd2752,32'd2816,32'd2880,32'd2944,32'd3008,32'd3072,32'd3136,32'd3200,32'd3264,32'd3328,32'd3392,32'd3456,32'd3520,32'd3584,32'd3648,32'd3712,32'd3776,32'd3840,32'd3904,32'd3968,32'd4032,32'd4096,32'd4160,32'd4224,32'd4288,32'd4352,32'd4416,32'd4480,32'd4544,32'd4608,32'd4672,32'd4736,32'd4800,32'd4864,32'd4928,32'd4992,32'd5056,32'd5120,32'd5184,32'd5248,32'd5312,32'd5376,32'd5440,32'd5504,32'd5568,32'd5632,32'd5696,32'd5760,32'd5824,32'd5888,32'd5952,32'd6016,32'd6080,32'd6144,32'd6208,32'd6272,32'd6336,32'd6400,32'd6464,32'd6528,32'd6592,32'd6656,32'd6720,32'd6784,32'd6848,32'd6912,32'd6976,32'd7040,32'd7104,32'd7168,32'd7232,32'd7296,32'd7360,32'd7424,32'd7488,32'd7552,32'd7616,32'd7680,32'd7744,32'd7808,32'd7872,32'd7936,32'd8000,32'd8064,32'd8128,32'd8192,32'd8256,32'd8320,32'd8384,32'd8448,32'd8512,32'd8576,32'd8640,32'd8704,32'd8768,32'd8832,32'd8896,32'd8960,32'd9024,32'd9088,32'd9152,32'd9216,32'd9280,32'd9344,32'd9408,32'd9472,32'd9536,32'd9600,32'd9664,32'd9728,32'd9792,32'd9856,32'd9920,32'd9984,32'd10048,32'd10112,32'd10176,32'd10240,32'd10304,32'd10368,32'd10432,32'd10496,32'd10560,32'd10624,32'd10688,32'd10752,32'd10816,32'd10880,32'd10944,32'd11008,32'd11072,32'd11136,32'd11200,32'd11264,32'd11328,32'd11392,32'd11456,32'd11520,32'd11584,32'd11648,32'd11712,32'd11776,32'd11840,32'd11904,32'd11968,32'd12032,32'd12096,32'd12160,32'd12224,32'd12288,32'd12352,32'd12416,32'd12480,32'd12544,32'd12608,32'd12672,32'd12736,32'd12800,32'd12864,32'd12928,32'd12992,32'd13056,32'd13120,32'd13184,32'd13248,32'd13312,32'd13376,32'd13440,32'd13504,32'd13568,32'd13632,32'd13696,32'd13760,32'd13824,32'd13888,32'd13952,32'd14016,32'd14080,32'd14144,32'd14208,32'd14272,32'd14336,32'd14400,32'd14464,32'd14528,32'd14592,32'd14656,32'd14720,32'd14784,32'd14848,32'd14912,32'd14976,32'd15040,32'd15104,32'd15168,32'd15232,32'd15296,32'd15360,32'd15424,32'd15488,32'd15552,32'd15616,32'd15680,32'd15744,32'd15808,32'd15872,32'd15936,32'd16000,32'd16064,32'd16128,32'd16192,32'd16256,32'd16320,32'd16384,32'd16448,32'd16512,32'd16576,32'd16640,32'd16704,32'd16768,32'd16832,32'd16896,32'd16960,32'd17024,32'd17088,32'd17152,32'd17216,32'd17280,32'd17344,32'd17408,32'd17472,32'd17536,32'd17600,32'd17664,32'd17728,32'd17792,32'd17856,32'd17920,32'd17984,32'd18048,32'd18112,32'd18176,32'd18240,32'd18304,32'd18368,32'd18432,32'd18496,32'd18560,32'd18624,32'd18688,32'd18752,32'd18816,32'd18880,32'd18944,32'd19008,32'd19072,32'd19136,32'd19200,32'd19264,32'd19328,32'd19392,32'd19456,32'd19520,32'd19584,32'd19648,32'd19712,32'd19776,32'd19840,32'd19904,32'd19968,32'd20032,32'd20096,32'd20160,32'd20224,32'd20288,32'd20352,32'd20416,32'd20480,32'd20544,32'd20608,32'd20672,32'd20736,32'd20800,32'd20864,32'd20928,32'd20992,32'd21056,32'd21120,32'd21184,32'd21248,32'd21312,32'd21376,32'd21440,32'd21504,32'd21568,32'd21632,32'd21696,32'd21760,32'd21824,32'd21888,32'd21952,32'd22016,32'd22080,32'd22144,32'd22208,32'd22272,32'd22336,32'd22400,32'd22464,32'd22528,32'd22592,32'd22656,32'd22720,32'd22784,32'd22848,32'd22912,32'd22976,32'd23040,32'd23104,32'd23168,32'd23232,32'd23296,32'd23360,32'd23424,32'd23488,32'd23552,32'd23616,32'd23680,32'd23744,32'd23808,32'd23872,32'd23936,32'd24000,32'd24064,32'd24128,32'd24192,32'd24256,32'd24320,32'd24384,32'd24448,32'd24512,32'd24576,32'd24640,32'd24704,32'd24768,32'd24832,32'd24896,32'd24960,32'd25024,32'd25088,32'd25152,32'd25216,32'd25280,32'd25344,32'd25408,32'd25472,32'd25536 };matrix[65]='{32'd0,32'd65,32'd130,32'd195,32'd260,32'd325,32'd390,32'd455,32'd520,32'd585,32'd650,32'd715,32'd780,32'd845,32'd910,32'd975,32'd1040,32'd1105,32'd1170,32'd1235,32'd1300,32'd1365,32'd1430,32'd1495,32'd1560,32'd1625,32'd1690,32'd1755,32'd1820,32'd1885,32'd1950,32'd2015,32'd2080,32'd2145,32'd2210,32'd2275,32'd2340,32'd2405,32'd2470,32'd2535,32'd2600,32'd2665,32'd2730,32'd2795,32'd2860,32'd2925,32'd2990,32'd3055,32'd3120,32'd3185,32'd3250,32'd3315,32'd3380,32'd3445,32'd3510,32'd3575,32'd3640,32'd3705,32'd3770,32'd3835,32'd3900,32'd3965,32'd4030,32'd4095,32'd4160,32'd4225,32'd4290,32'd4355,32'd4420,32'd4485,32'd4550,32'd4615,32'd4680,32'd4745,32'd4810,32'd4875,32'd4940,32'd5005,32'd5070,32'd5135,32'd5200,32'd5265,32'd5330,32'd5395,32'd5460,32'd5525,32'd5590,32'd5655,32'd5720,32'd5785,32'd5850,32'd5915,32'd5980,32'd6045,32'd6110,32'd6175,32'd6240,32'd6305,32'd6370,32'd6435,32'd6500,32'd6565,32'd6630,32'd6695,32'd6760,32'd6825,32'd6890,32'd6955,32'd7020,32'd7085,32'd7150,32'd7215,32'd7280,32'd7345,32'd7410,32'd7475,32'd7540,32'd7605,32'd7670,32'd7735,32'd7800,32'd7865,32'd7930,32'd7995,32'd8060,32'd8125,32'd8190,32'd8255,32'd8320,32'd8385,32'd8450,32'd8515,32'd8580,32'd8645,32'd8710,32'd8775,32'd8840,32'd8905,32'd8970,32'd9035,32'd9100,32'd9165,32'd9230,32'd9295,32'd9360,32'd9425,32'd9490,32'd9555,32'd9620,32'd9685,32'd9750,32'd9815,32'd9880,32'd9945,32'd10010,32'd10075,32'd10140,32'd10205,32'd10270,32'd10335,32'd10400,32'd10465,32'd10530,32'd10595,32'd10660,32'd10725,32'd10790,32'd10855,32'd10920,32'd10985,32'd11050,32'd11115,32'd11180,32'd11245,32'd11310,32'd11375,32'd11440,32'd11505,32'd11570,32'd11635,32'd11700,32'd11765,32'd11830,32'd11895,32'd11960,32'd12025,32'd12090,32'd12155,32'd12220,32'd12285,32'd12350,32'd12415,32'd12480,32'd12545,32'd12610,32'd12675,32'd12740,32'd12805,32'd12870,32'd12935,32'd13000,32'd13065,32'd13130,32'd13195,32'd13260,32'd13325,32'd13390,32'd13455,32'd13520,32'd13585,32'd13650,32'd13715,32'd13780,32'd13845,32'd13910,32'd13975,32'd14040,32'd14105,32'd14170,32'd14235,32'd14300,32'd14365,32'd14430,32'd14495,32'd14560,32'd14625,32'd14690,32'd14755,32'd14820,32'd14885,32'd14950,32'd15015,32'd15080,32'd15145,32'd15210,32'd15275,32'd15340,32'd15405,32'd15470,32'd15535,32'd15600,32'd15665,32'd15730,32'd15795,32'd15860,32'd15925,32'd15990,32'd16055,32'd16120,32'd16185,32'd16250,32'd16315,32'd16380,32'd16445,32'd16510,32'd16575,32'd16640,32'd16705,32'd16770,32'd16835,32'd16900,32'd16965,32'd17030,32'd17095,32'd17160,32'd17225,32'd17290,32'd17355,32'd17420,32'd17485,32'd17550,32'd17615,32'd17680,32'd17745,32'd17810,32'd17875,32'd17940,32'd18005,32'd18070,32'd18135,32'd18200,32'd18265,32'd18330,32'd18395,32'd18460,32'd18525,32'd18590,32'd18655,32'd18720,32'd18785,32'd18850,32'd18915,32'd18980,32'd19045,32'd19110,32'd19175,32'd19240,32'd19305,32'd19370,32'd19435,32'd19500,32'd19565,32'd19630,32'd19695,32'd19760,32'd19825,32'd19890,32'd19955,32'd20020,32'd20085,32'd20150,32'd20215,32'd20280,32'd20345,32'd20410,32'd20475,32'd20540,32'd20605,32'd20670,32'd20735,32'd20800,32'd20865,32'd20930,32'd20995,32'd21060,32'd21125,32'd21190,32'd21255,32'd21320,32'd21385,32'd21450,32'd21515,32'd21580,32'd21645,32'd21710,32'd21775,32'd21840,32'd21905,32'd21970,32'd22035,32'd22100,32'd22165,32'd22230,32'd22295,32'd22360,32'd22425,32'd22490,32'd22555,32'd22620,32'd22685,32'd22750,32'd22815,32'd22880,32'd22945,32'd23010,32'd23075,32'd23140,32'd23205,32'd23270,32'd23335,32'd23400,32'd23465,32'd23530,32'd23595,32'd23660,32'd23725,32'd23790,32'd23855,32'd23920,32'd23985,32'd24050,32'd24115,32'd24180,32'd24245,32'd24310,32'd24375,32'd24440,32'd24505,32'd24570,32'd24635,32'd24700,32'd24765,32'd24830,32'd24895,32'd24960,32'd25025,32'd25090,32'd25155,32'd25220,32'd25285,32'd25350,32'd25415,32'd25480,32'd25545,32'd25610,32'd25675,32'd25740,32'd25805,32'd25870,32'd25935 };matrix[66]='{32'd0,32'd66,32'd132,32'd198,32'd264,32'd330,32'd396,32'd462,32'd528,32'd594,32'd660,32'd726,32'd792,32'd858,32'd924,32'd990,32'd1056,32'd1122,32'd1188,32'd1254,32'd1320,32'd1386,32'd1452,32'd1518,32'd1584,32'd1650,32'd1716,32'd1782,32'd1848,32'd1914,32'd1980,32'd2046,32'd2112,32'd2178,32'd2244,32'd2310,32'd2376,32'd2442,32'd2508,32'd2574,32'd2640,32'd2706,32'd2772,32'd2838,32'd2904,32'd2970,32'd3036,32'd3102,32'd3168,32'd3234,32'd3300,32'd3366,32'd3432,32'd3498,32'd3564,32'd3630,32'd3696,32'd3762,32'd3828,32'd3894,32'd3960,32'd4026,32'd4092,32'd4158,32'd4224,32'd4290,32'd4356,32'd4422,32'd4488,32'd4554,32'd4620,32'd4686,32'd4752,32'd4818,32'd4884,32'd4950,32'd5016,32'd5082,32'd5148,32'd5214,32'd5280,32'd5346,32'd5412,32'd5478,32'd5544,32'd5610,32'd5676,32'd5742,32'd5808,32'd5874,32'd5940,32'd6006,32'd6072,32'd6138,32'd6204,32'd6270,32'd6336,32'd6402,32'd6468,32'd6534,32'd6600,32'd6666,32'd6732,32'd6798,32'd6864,32'd6930,32'd6996,32'd7062,32'd7128,32'd7194,32'd7260,32'd7326,32'd7392,32'd7458,32'd7524,32'd7590,32'd7656,32'd7722,32'd7788,32'd7854,32'd7920,32'd7986,32'd8052,32'd8118,32'd8184,32'd8250,32'd8316,32'd8382,32'd8448,32'd8514,32'd8580,32'd8646,32'd8712,32'd8778,32'd8844,32'd8910,32'd8976,32'd9042,32'd9108,32'd9174,32'd9240,32'd9306,32'd9372,32'd9438,32'd9504,32'd9570,32'd9636,32'd9702,32'd9768,32'd9834,32'd9900,32'd9966,32'd10032,32'd10098,32'd10164,32'd10230,32'd10296,32'd10362,32'd10428,32'd10494,32'd10560,32'd10626,32'd10692,32'd10758,32'd10824,32'd10890,32'd10956,32'd11022,32'd11088,32'd11154,32'd11220,32'd11286,32'd11352,32'd11418,32'd11484,32'd11550,32'd11616,32'd11682,32'd11748,32'd11814,32'd11880,32'd11946,32'd12012,32'd12078,32'd12144,32'd12210,32'd12276,32'd12342,32'd12408,32'd12474,32'd12540,32'd12606,32'd12672,32'd12738,32'd12804,32'd12870,32'd12936,32'd13002,32'd13068,32'd13134,32'd13200,32'd13266,32'd13332,32'd13398,32'd13464,32'd13530,32'd13596,32'd13662,32'd13728,32'd13794,32'd13860,32'd13926,32'd13992,32'd14058,32'd14124,32'd14190,32'd14256,32'd14322,32'd14388,32'd14454,32'd14520,32'd14586,32'd14652,32'd14718,32'd14784,32'd14850,32'd14916,32'd14982,32'd15048,32'd15114,32'd15180,32'd15246,32'd15312,32'd15378,32'd15444,32'd15510,32'd15576,32'd15642,32'd15708,32'd15774,32'd15840,32'd15906,32'd15972,32'd16038,32'd16104,32'd16170,32'd16236,32'd16302,32'd16368,32'd16434,32'd16500,32'd16566,32'd16632,32'd16698,32'd16764,32'd16830,32'd16896,32'd16962,32'd17028,32'd17094,32'd17160,32'd17226,32'd17292,32'd17358,32'd17424,32'd17490,32'd17556,32'd17622,32'd17688,32'd17754,32'd17820,32'd17886,32'd17952,32'd18018,32'd18084,32'd18150,32'd18216,32'd18282,32'd18348,32'd18414,32'd18480,32'd18546,32'd18612,32'd18678,32'd18744,32'd18810,32'd18876,32'd18942,32'd19008,32'd19074,32'd19140,32'd19206,32'd19272,32'd19338,32'd19404,32'd19470,32'd19536,32'd19602,32'd19668,32'd19734,32'd19800,32'd19866,32'd19932,32'd19998,32'd20064,32'd20130,32'd20196,32'd20262,32'd20328,32'd20394,32'd20460,32'd20526,32'd20592,32'd20658,32'd20724,32'd20790,32'd20856,32'd20922,32'd20988,32'd21054,32'd21120,32'd21186,32'd21252,32'd21318,32'd21384,32'd21450,32'd21516,32'd21582,32'd21648,32'd21714,32'd21780,32'd21846,32'd21912,32'd21978,32'd22044,32'd22110,32'd22176,32'd22242,32'd22308,32'd22374,32'd22440,32'd22506,32'd22572,32'd22638,32'd22704,32'd22770,32'd22836,32'd22902,32'd22968,32'd23034,32'd23100,32'd23166,32'd23232,32'd23298,32'd23364,32'd23430,32'd23496,32'd23562,32'd23628,32'd23694,32'd23760,32'd23826,32'd23892,32'd23958,32'd24024,32'd24090,32'd24156,32'd24222,32'd24288,32'd24354,32'd24420,32'd24486,32'd24552,32'd24618,32'd24684,32'd24750,32'd24816,32'd24882,32'd24948,32'd25014,32'd25080,32'd25146,32'd25212,32'd25278,32'd25344,32'd25410,32'd25476,32'd25542,32'd25608,32'd25674,32'd25740,32'd25806,32'd25872,32'd25938,32'd26004,32'd26070,32'd26136,32'd26202,32'd26268,32'd26334 };matrix[67]='{32'd0,32'd67,32'd134,32'd201,32'd268,32'd335,32'd402,32'd469,32'd536,32'd603,32'd670,32'd737,32'd804,32'd871,32'd938,32'd1005,32'd1072,32'd1139,32'd1206,32'd1273,32'd1340,32'd1407,32'd1474,32'd1541,32'd1608,32'd1675,32'd1742,32'd1809,32'd1876,32'd1943,32'd2010,32'd2077,32'd2144,32'd2211,32'd2278,32'd2345,32'd2412,32'd2479,32'd2546,32'd2613,32'd2680,32'd2747,32'd2814,32'd2881,32'd2948,32'd3015,32'd3082,32'd3149,32'd3216,32'd3283,32'd3350,32'd3417,32'd3484,32'd3551,32'd3618,32'd3685,32'd3752,32'd3819,32'd3886,32'd3953,32'd4020,32'd4087,32'd4154,32'd4221,32'd4288,32'd4355,32'd4422,32'd4489,32'd4556,32'd4623,32'd4690,32'd4757,32'd4824,32'd4891,32'd4958,32'd5025,32'd5092,32'd5159,32'd5226,32'd5293,32'd5360,32'd5427,32'd5494,32'd5561,32'd5628,32'd5695,32'd5762,32'd5829,32'd5896,32'd5963,32'd6030,32'd6097,32'd6164,32'd6231,32'd6298,32'd6365,32'd6432,32'd6499,32'd6566,32'd6633,32'd6700,32'd6767,32'd6834,32'd6901,32'd6968,32'd7035,32'd7102,32'd7169,32'd7236,32'd7303,32'd7370,32'd7437,32'd7504,32'd7571,32'd7638,32'd7705,32'd7772,32'd7839,32'd7906,32'd7973,32'd8040,32'd8107,32'd8174,32'd8241,32'd8308,32'd8375,32'd8442,32'd8509,32'd8576,32'd8643,32'd8710,32'd8777,32'd8844,32'd8911,32'd8978,32'd9045,32'd9112,32'd9179,32'd9246,32'd9313,32'd9380,32'd9447,32'd9514,32'd9581,32'd9648,32'd9715,32'd9782,32'd9849,32'd9916,32'd9983,32'd10050,32'd10117,32'd10184,32'd10251,32'd10318,32'd10385,32'd10452,32'd10519,32'd10586,32'd10653,32'd10720,32'd10787,32'd10854,32'd10921,32'd10988,32'd11055,32'd11122,32'd11189,32'd11256,32'd11323,32'd11390,32'd11457,32'd11524,32'd11591,32'd11658,32'd11725,32'd11792,32'd11859,32'd11926,32'd11993,32'd12060,32'd12127,32'd12194,32'd12261,32'd12328,32'd12395,32'd12462,32'd12529,32'd12596,32'd12663,32'd12730,32'd12797,32'd12864,32'd12931,32'd12998,32'd13065,32'd13132,32'd13199,32'd13266,32'd13333,32'd13400,32'd13467,32'd13534,32'd13601,32'd13668,32'd13735,32'd13802,32'd13869,32'd13936,32'd14003,32'd14070,32'd14137,32'd14204,32'd14271,32'd14338,32'd14405,32'd14472,32'd14539,32'd14606,32'd14673,32'd14740,32'd14807,32'd14874,32'd14941,32'd15008,32'd15075,32'd15142,32'd15209,32'd15276,32'd15343,32'd15410,32'd15477,32'd15544,32'd15611,32'd15678,32'd15745,32'd15812,32'd15879,32'd15946,32'd16013,32'd16080,32'd16147,32'd16214,32'd16281,32'd16348,32'd16415,32'd16482,32'd16549,32'd16616,32'd16683,32'd16750,32'd16817,32'd16884,32'd16951,32'd17018,32'd17085,32'd17152,32'd17219,32'd17286,32'd17353,32'd17420,32'd17487,32'd17554,32'd17621,32'd17688,32'd17755,32'd17822,32'd17889,32'd17956,32'd18023,32'd18090,32'd18157,32'd18224,32'd18291,32'd18358,32'd18425,32'd18492,32'd18559,32'd18626,32'd18693,32'd18760,32'd18827,32'd18894,32'd18961,32'd19028,32'd19095,32'd19162,32'd19229,32'd19296,32'd19363,32'd19430,32'd19497,32'd19564,32'd19631,32'd19698,32'd19765,32'd19832,32'd19899,32'd19966,32'd20033,32'd20100,32'd20167,32'd20234,32'd20301,32'd20368,32'd20435,32'd20502,32'd20569,32'd20636,32'd20703,32'd20770,32'd20837,32'd20904,32'd20971,32'd21038,32'd21105,32'd21172,32'd21239,32'd21306,32'd21373,32'd21440,32'd21507,32'd21574,32'd21641,32'd21708,32'd21775,32'd21842,32'd21909,32'd21976,32'd22043,32'd22110,32'd22177,32'd22244,32'd22311,32'd22378,32'd22445,32'd22512,32'd22579,32'd22646,32'd22713,32'd22780,32'd22847,32'd22914,32'd22981,32'd23048,32'd23115,32'd23182,32'd23249,32'd23316,32'd23383,32'd23450,32'd23517,32'd23584,32'd23651,32'd23718,32'd23785,32'd23852,32'd23919,32'd23986,32'd24053,32'd24120,32'd24187,32'd24254,32'd24321,32'd24388,32'd24455,32'd24522,32'd24589,32'd24656,32'd24723,32'd24790,32'd24857,32'd24924,32'd24991,32'd25058,32'd25125,32'd25192,32'd25259,32'd25326,32'd25393,32'd25460,32'd25527,32'd25594,32'd25661,32'd25728,32'd25795,32'd25862,32'd25929,32'd25996,32'd26063,32'd26130,32'd26197,32'd26264,32'd26331,32'd26398,32'd26465,32'd26532,32'd26599,32'd26666,32'd26733 };matrix[68]='{32'd0,32'd68,32'd136,32'd204,32'd272,32'd340,32'd408,32'd476,32'd544,32'd612,32'd680,32'd748,32'd816,32'd884,32'd952,32'd1020,32'd1088,32'd1156,32'd1224,32'd1292,32'd1360,32'd1428,32'd1496,32'd1564,32'd1632,32'd1700,32'd1768,32'd1836,32'd1904,32'd1972,32'd2040,32'd2108,32'd2176,32'd2244,32'd2312,32'd2380,32'd2448,32'd2516,32'd2584,32'd2652,32'd2720,32'd2788,32'd2856,32'd2924,32'd2992,32'd3060,32'd3128,32'd3196,32'd3264,32'd3332,32'd3400,32'd3468,32'd3536,32'd3604,32'd3672,32'd3740,32'd3808,32'd3876,32'd3944,32'd4012,32'd4080,32'd4148,32'd4216,32'd4284,32'd4352,32'd4420,32'd4488,32'd4556,32'd4624,32'd4692,32'd4760,32'd4828,32'd4896,32'd4964,32'd5032,32'd5100,32'd5168,32'd5236,32'd5304,32'd5372,32'd5440,32'd5508,32'd5576,32'd5644,32'd5712,32'd5780,32'd5848,32'd5916,32'd5984,32'd6052,32'd6120,32'd6188,32'd6256,32'd6324,32'd6392,32'd6460,32'd6528,32'd6596,32'd6664,32'd6732,32'd6800,32'd6868,32'd6936,32'd7004,32'd7072,32'd7140,32'd7208,32'd7276,32'd7344,32'd7412,32'd7480,32'd7548,32'd7616,32'd7684,32'd7752,32'd7820,32'd7888,32'd7956,32'd8024,32'd8092,32'd8160,32'd8228,32'd8296,32'd8364,32'd8432,32'd8500,32'd8568,32'd8636,32'd8704,32'd8772,32'd8840,32'd8908,32'd8976,32'd9044,32'd9112,32'd9180,32'd9248,32'd9316,32'd9384,32'd9452,32'd9520,32'd9588,32'd9656,32'd9724,32'd9792,32'd9860,32'd9928,32'd9996,32'd10064,32'd10132,32'd10200,32'd10268,32'd10336,32'd10404,32'd10472,32'd10540,32'd10608,32'd10676,32'd10744,32'd10812,32'd10880,32'd10948,32'd11016,32'd11084,32'd11152,32'd11220,32'd11288,32'd11356,32'd11424,32'd11492,32'd11560,32'd11628,32'd11696,32'd11764,32'd11832,32'd11900,32'd11968,32'd12036,32'd12104,32'd12172,32'd12240,32'd12308,32'd12376,32'd12444,32'd12512,32'd12580,32'd12648,32'd12716,32'd12784,32'd12852,32'd12920,32'd12988,32'd13056,32'd13124,32'd13192,32'd13260,32'd13328,32'd13396,32'd13464,32'd13532,32'd13600,32'd13668,32'd13736,32'd13804,32'd13872,32'd13940,32'd14008,32'd14076,32'd14144,32'd14212,32'd14280,32'd14348,32'd14416,32'd14484,32'd14552,32'd14620,32'd14688,32'd14756,32'd14824,32'd14892,32'd14960,32'd15028,32'd15096,32'd15164,32'd15232,32'd15300,32'd15368,32'd15436,32'd15504,32'd15572,32'd15640,32'd15708,32'd15776,32'd15844,32'd15912,32'd15980,32'd16048,32'd16116,32'd16184,32'd16252,32'd16320,32'd16388,32'd16456,32'd16524,32'd16592,32'd16660,32'd16728,32'd16796,32'd16864,32'd16932,32'd17000,32'd17068,32'd17136,32'd17204,32'd17272,32'd17340,32'd17408,32'd17476,32'd17544,32'd17612,32'd17680,32'd17748,32'd17816,32'd17884,32'd17952,32'd18020,32'd18088,32'd18156,32'd18224,32'd18292,32'd18360,32'd18428,32'd18496,32'd18564,32'd18632,32'd18700,32'd18768,32'd18836,32'd18904,32'd18972,32'd19040,32'd19108,32'd19176,32'd19244,32'd19312,32'd19380,32'd19448,32'd19516,32'd19584,32'd19652,32'd19720,32'd19788,32'd19856,32'd19924,32'd19992,32'd20060,32'd20128,32'd20196,32'd20264,32'd20332,32'd20400,32'd20468,32'd20536,32'd20604,32'd20672,32'd20740,32'd20808,32'd20876,32'd20944,32'd21012,32'd21080,32'd21148,32'd21216,32'd21284,32'd21352,32'd21420,32'd21488,32'd21556,32'd21624,32'd21692,32'd21760,32'd21828,32'd21896,32'd21964,32'd22032,32'd22100,32'd22168,32'd22236,32'd22304,32'd22372,32'd22440,32'd22508,32'd22576,32'd22644,32'd22712,32'd22780,32'd22848,32'd22916,32'd22984,32'd23052,32'd23120,32'd23188,32'd23256,32'd23324,32'd23392,32'd23460,32'd23528,32'd23596,32'd23664,32'd23732,32'd23800,32'd23868,32'd23936,32'd24004,32'd24072,32'd24140,32'd24208,32'd24276,32'd24344,32'd24412,32'd24480,32'd24548,32'd24616,32'd24684,32'd24752,32'd24820,32'd24888,32'd24956,32'd25024,32'd25092,32'd25160,32'd25228,32'd25296,32'd25364,32'd25432,32'd25500,32'd25568,32'd25636,32'd25704,32'd25772,32'd25840,32'd25908,32'd25976,32'd26044,32'd26112,32'd26180,32'd26248,32'd26316,32'd26384,32'd26452,32'd26520,32'd26588,32'd26656,32'd26724,32'd26792,32'd26860,32'd26928,32'd26996,32'd27064,32'd27132 };matrix[69]='{32'd0,32'd69,32'd138,32'd207,32'd276,32'd345,32'd414,32'd483,32'd552,32'd621,32'd690,32'd759,32'd828,32'd897,32'd966,32'd1035,32'd1104,32'd1173,32'd1242,32'd1311,32'd1380,32'd1449,32'd1518,32'd1587,32'd1656,32'd1725,32'd1794,32'd1863,32'd1932,32'd2001,32'd2070,32'd2139,32'd2208,32'd2277,32'd2346,32'd2415,32'd2484,32'd2553,32'd2622,32'd2691,32'd2760,32'd2829,32'd2898,32'd2967,32'd3036,32'd3105,32'd3174,32'd3243,32'd3312,32'd3381,32'd3450,32'd3519,32'd3588,32'd3657,32'd3726,32'd3795,32'd3864,32'd3933,32'd4002,32'd4071,32'd4140,32'd4209,32'd4278,32'd4347,32'd4416,32'd4485,32'd4554,32'd4623,32'd4692,32'd4761,32'd4830,32'd4899,32'd4968,32'd5037,32'd5106,32'd5175,32'd5244,32'd5313,32'd5382,32'd5451,32'd5520,32'd5589,32'd5658,32'd5727,32'd5796,32'd5865,32'd5934,32'd6003,32'd6072,32'd6141,32'd6210,32'd6279,32'd6348,32'd6417,32'd6486,32'd6555,32'd6624,32'd6693,32'd6762,32'd6831,32'd6900,32'd6969,32'd7038,32'd7107,32'd7176,32'd7245,32'd7314,32'd7383,32'd7452,32'd7521,32'd7590,32'd7659,32'd7728,32'd7797,32'd7866,32'd7935,32'd8004,32'd8073,32'd8142,32'd8211,32'd8280,32'd8349,32'd8418,32'd8487,32'd8556,32'd8625,32'd8694,32'd8763,32'd8832,32'd8901,32'd8970,32'd9039,32'd9108,32'd9177,32'd9246,32'd9315,32'd9384,32'd9453,32'd9522,32'd9591,32'd9660,32'd9729,32'd9798,32'd9867,32'd9936,32'd10005,32'd10074,32'd10143,32'd10212,32'd10281,32'd10350,32'd10419,32'd10488,32'd10557,32'd10626,32'd10695,32'd10764,32'd10833,32'd10902,32'd10971,32'd11040,32'd11109,32'd11178,32'd11247,32'd11316,32'd11385,32'd11454,32'd11523,32'd11592,32'd11661,32'd11730,32'd11799,32'd11868,32'd11937,32'd12006,32'd12075,32'd12144,32'd12213,32'd12282,32'd12351,32'd12420,32'd12489,32'd12558,32'd12627,32'd12696,32'd12765,32'd12834,32'd12903,32'd12972,32'd13041,32'd13110,32'd13179,32'd13248,32'd13317,32'd13386,32'd13455,32'd13524,32'd13593,32'd13662,32'd13731,32'd13800,32'd13869,32'd13938,32'd14007,32'd14076,32'd14145,32'd14214,32'd14283,32'd14352,32'd14421,32'd14490,32'd14559,32'd14628,32'd14697,32'd14766,32'd14835,32'd14904,32'd14973,32'd15042,32'd15111,32'd15180,32'd15249,32'd15318,32'd15387,32'd15456,32'd15525,32'd15594,32'd15663,32'd15732,32'd15801,32'd15870,32'd15939,32'd16008,32'd16077,32'd16146,32'd16215,32'd16284,32'd16353,32'd16422,32'd16491,32'd16560,32'd16629,32'd16698,32'd16767,32'd16836,32'd16905,32'd16974,32'd17043,32'd17112,32'd17181,32'd17250,32'd17319,32'd17388,32'd17457,32'd17526,32'd17595,32'd17664,32'd17733,32'd17802,32'd17871,32'd17940,32'd18009,32'd18078,32'd18147,32'd18216,32'd18285,32'd18354,32'd18423,32'd18492,32'd18561,32'd18630,32'd18699,32'd18768,32'd18837,32'd18906,32'd18975,32'd19044,32'd19113,32'd19182,32'd19251,32'd19320,32'd19389,32'd19458,32'd19527,32'd19596,32'd19665,32'd19734,32'd19803,32'd19872,32'd19941,32'd20010,32'd20079,32'd20148,32'd20217,32'd20286,32'd20355,32'd20424,32'd20493,32'd20562,32'd20631,32'd20700,32'd20769,32'd20838,32'd20907,32'd20976,32'd21045,32'd21114,32'd21183,32'd21252,32'd21321,32'd21390,32'd21459,32'd21528,32'd21597,32'd21666,32'd21735,32'd21804,32'd21873,32'd21942,32'd22011,32'd22080,32'd22149,32'd22218,32'd22287,32'd22356,32'd22425,32'd22494,32'd22563,32'd22632,32'd22701,32'd22770,32'd22839,32'd22908,32'd22977,32'd23046,32'd23115,32'd23184,32'd23253,32'd23322,32'd23391,32'd23460,32'd23529,32'd23598,32'd23667,32'd23736,32'd23805,32'd23874,32'd23943,32'd24012,32'd24081,32'd24150,32'd24219,32'd24288,32'd24357,32'd24426,32'd24495,32'd24564,32'd24633,32'd24702,32'd24771,32'd24840,32'd24909,32'd24978,32'd25047,32'd25116,32'd25185,32'd25254,32'd25323,32'd25392,32'd25461,32'd25530,32'd25599,32'd25668,32'd25737,32'd25806,32'd25875,32'd25944,32'd26013,32'd26082,32'd26151,32'd26220,32'd26289,32'd26358,32'd26427,32'd26496,32'd26565,32'd26634,32'd26703,32'd26772,32'd26841,32'd26910,32'd26979,32'd27048,32'd27117,32'd27186,32'd27255,32'd27324,32'd27393,32'd27462,32'd27531 };matrix[70]='{32'd0,32'd70,32'd140,32'd210,32'd280,32'd350,32'd420,32'd490,32'd560,32'd630,32'd700,32'd770,32'd840,32'd910,32'd980,32'd1050,32'd1120,32'd1190,32'd1260,32'd1330,32'd1400,32'd1470,32'd1540,32'd1610,32'd1680,32'd1750,32'd1820,32'd1890,32'd1960,32'd2030,32'd2100,32'd2170,32'd2240,32'd2310,32'd2380,32'd2450,32'd2520,32'd2590,32'd2660,32'd2730,32'd2800,32'd2870,32'd2940,32'd3010,32'd3080,32'd3150,32'd3220,32'd3290,32'd3360,32'd3430,32'd3500,32'd3570,32'd3640,32'd3710,32'd3780,32'd3850,32'd3920,32'd3990,32'd4060,32'd4130,32'd4200,32'd4270,32'd4340,32'd4410,32'd4480,32'd4550,32'd4620,32'd4690,32'd4760,32'd4830,32'd4900,32'd4970,32'd5040,32'd5110,32'd5180,32'd5250,32'd5320,32'd5390,32'd5460,32'd5530,32'd5600,32'd5670,32'd5740,32'd5810,32'd5880,32'd5950,32'd6020,32'd6090,32'd6160,32'd6230,32'd6300,32'd6370,32'd6440,32'd6510,32'd6580,32'd6650,32'd6720,32'd6790,32'd6860,32'd6930,32'd7000,32'd7070,32'd7140,32'd7210,32'd7280,32'd7350,32'd7420,32'd7490,32'd7560,32'd7630,32'd7700,32'd7770,32'd7840,32'd7910,32'd7980,32'd8050,32'd8120,32'd8190,32'd8260,32'd8330,32'd8400,32'd8470,32'd8540,32'd8610,32'd8680,32'd8750,32'd8820,32'd8890,32'd8960,32'd9030,32'd9100,32'd9170,32'd9240,32'd9310,32'd9380,32'd9450,32'd9520,32'd9590,32'd9660,32'd9730,32'd9800,32'd9870,32'd9940,32'd10010,32'd10080,32'd10150,32'd10220,32'd10290,32'd10360,32'd10430,32'd10500,32'd10570,32'd10640,32'd10710,32'd10780,32'd10850,32'd10920,32'd10990,32'd11060,32'd11130,32'd11200,32'd11270,32'd11340,32'd11410,32'd11480,32'd11550,32'd11620,32'd11690,32'd11760,32'd11830,32'd11900,32'd11970,32'd12040,32'd12110,32'd12180,32'd12250,32'd12320,32'd12390,32'd12460,32'd12530,32'd12600,32'd12670,32'd12740,32'd12810,32'd12880,32'd12950,32'd13020,32'd13090,32'd13160,32'd13230,32'd13300,32'd13370,32'd13440,32'd13510,32'd13580,32'd13650,32'd13720,32'd13790,32'd13860,32'd13930,32'd14000,32'd14070,32'd14140,32'd14210,32'd14280,32'd14350,32'd14420,32'd14490,32'd14560,32'd14630,32'd14700,32'd14770,32'd14840,32'd14910,32'd14980,32'd15050,32'd15120,32'd15190,32'd15260,32'd15330,32'd15400,32'd15470,32'd15540,32'd15610,32'd15680,32'd15750,32'd15820,32'd15890,32'd15960,32'd16030,32'd16100,32'd16170,32'd16240,32'd16310,32'd16380,32'd16450,32'd16520,32'd16590,32'd16660,32'd16730,32'd16800,32'd16870,32'd16940,32'd17010,32'd17080,32'd17150,32'd17220,32'd17290,32'd17360,32'd17430,32'd17500,32'd17570,32'd17640,32'd17710,32'd17780,32'd17850,32'd17920,32'd17990,32'd18060,32'd18130,32'd18200,32'd18270,32'd18340,32'd18410,32'd18480,32'd18550,32'd18620,32'd18690,32'd18760,32'd18830,32'd18900,32'd18970,32'd19040,32'd19110,32'd19180,32'd19250,32'd19320,32'd19390,32'd19460,32'd19530,32'd19600,32'd19670,32'd19740,32'd19810,32'd19880,32'd19950,32'd20020,32'd20090,32'd20160,32'd20230,32'd20300,32'd20370,32'd20440,32'd20510,32'd20580,32'd20650,32'd20720,32'd20790,32'd20860,32'd20930,32'd21000,32'd21070,32'd21140,32'd21210,32'd21280,32'd21350,32'd21420,32'd21490,32'd21560,32'd21630,32'd21700,32'd21770,32'd21840,32'd21910,32'd21980,32'd22050,32'd22120,32'd22190,32'd22260,32'd22330,32'd22400,32'd22470,32'd22540,32'd22610,32'd22680,32'd22750,32'd22820,32'd22890,32'd22960,32'd23030,32'd23100,32'd23170,32'd23240,32'd23310,32'd23380,32'd23450,32'd23520,32'd23590,32'd23660,32'd23730,32'd23800,32'd23870,32'd23940,32'd24010,32'd24080,32'd24150,32'd24220,32'd24290,32'd24360,32'd24430,32'd24500,32'd24570,32'd24640,32'd24710,32'd24780,32'd24850,32'd24920,32'd24990,32'd25060,32'd25130,32'd25200,32'd25270,32'd25340,32'd25410,32'd25480,32'd25550,32'd25620,32'd25690,32'd25760,32'd25830,32'd25900,32'd25970,32'd26040,32'd26110,32'd26180,32'd26250,32'd26320,32'd26390,32'd26460,32'd26530,32'd26600,32'd26670,32'd26740,32'd26810,32'd26880,32'd26950,32'd27020,32'd27090,32'd27160,32'd27230,32'd27300,32'd27370,32'd27440,32'd27510,32'd27580,32'd27650,32'd27720,32'd27790,32'd27860,32'd27930 };matrix[71]='{32'd0,32'd71,32'd142,32'd213,32'd284,32'd355,32'd426,32'd497,32'd568,32'd639,32'd710,32'd781,32'd852,32'd923,32'd994,32'd1065,32'd1136,32'd1207,32'd1278,32'd1349,32'd1420,32'd1491,32'd1562,32'd1633,32'd1704,32'd1775,32'd1846,32'd1917,32'd1988,32'd2059,32'd2130,32'd2201,32'd2272,32'd2343,32'd2414,32'd2485,32'd2556,32'd2627,32'd2698,32'd2769,32'd2840,32'd2911,32'd2982,32'd3053,32'd3124,32'd3195,32'd3266,32'd3337,32'd3408,32'd3479,32'd3550,32'd3621,32'd3692,32'd3763,32'd3834,32'd3905,32'd3976,32'd4047,32'd4118,32'd4189,32'd4260,32'd4331,32'd4402,32'd4473,32'd4544,32'd4615,32'd4686,32'd4757,32'd4828,32'd4899,32'd4970,32'd5041,32'd5112,32'd5183,32'd5254,32'd5325,32'd5396,32'd5467,32'd5538,32'd5609,32'd5680,32'd5751,32'd5822,32'd5893,32'd5964,32'd6035,32'd6106,32'd6177,32'd6248,32'd6319,32'd6390,32'd6461,32'd6532,32'd6603,32'd6674,32'd6745,32'd6816,32'd6887,32'd6958,32'd7029,32'd7100,32'd7171,32'd7242,32'd7313,32'd7384,32'd7455,32'd7526,32'd7597,32'd7668,32'd7739,32'd7810,32'd7881,32'd7952,32'd8023,32'd8094,32'd8165,32'd8236,32'd8307,32'd8378,32'd8449,32'd8520,32'd8591,32'd8662,32'd8733,32'd8804,32'd8875,32'd8946,32'd9017,32'd9088,32'd9159,32'd9230,32'd9301,32'd9372,32'd9443,32'd9514,32'd9585,32'd9656,32'd9727,32'd9798,32'd9869,32'd9940,32'd10011,32'd10082,32'd10153,32'd10224,32'd10295,32'd10366,32'd10437,32'd10508,32'd10579,32'd10650,32'd10721,32'd10792,32'd10863,32'd10934,32'd11005,32'd11076,32'd11147,32'd11218,32'd11289,32'd11360,32'd11431,32'd11502,32'd11573,32'd11644,32'd11715,32'd11786,32'd11857,32'd11928,32'd11999,32'd12070,32'd12141,32'd12212,32'd12283,32'd12354,32'd12425,32'd12496,32'd12567,32'd12638,32'd12709,32'd12780,32'd12851,32'd12922,32'd12993,32'd13064,32'd13135,32'd13206,32'd13277,32'd13348,32'd13419,32'd13490,32'd13561,32'd13632,32'd13703,32'd13774,32'd13845,32'd13916,32'd13987,32'd14058,32'd14129,32'd14200,32'd14271,32'd14342,32'd14413,32'd14484,32'd14555,32'd14626,32'd14697,32'd14768,32'd14839,32'd14910,32'd14981,32'd15052,32'd15123,32'd15194,32'd15265,32'd15336,32'd15407,32'd15478,32'd15549,32'd15620,32'd15691,32'd15762,32'd15833,32'd15904,32'd15975,32'd16046,32'd16117,32'd16188,32'd16259,32'd16330,32'd16401,32'd16472,32'd16543,32'd16614,32'd16685,32'd16756,32'd16827,32'd16898,32'd16969,32'd17040,32'd17111,32'd17182,32'd17253,32'd17324,32'd17395,32'd17466,32'd17537,32'd17608,32'd17679,32'd17750,32'd17821,32'd17892,32'd17963,32'd18034,32'd18105,32'd18176,32'd18247,32'd18318,32'd18389,32'd18460,32'd18531,32'd18602,32'd18673,32'd18744,32'd18815,32'd18886,32'd18957,32'd19028,32'd19099,32'd19170,32'd19241,32'd19312,32'd19383,32'd19454,32'd19525,32'd19596,32'd19667,32'd19738,32'd19809,32'd19880,32'd19951,32'd20022,32'd20093,32'd20164,32'd20235,32'd20306,32'd20377,32'd20448,32'd20519,32'd20590,32'd20661,32'd20732,32'd20803,32'd20874,32'd20945,32'd21016,32'd21087,32'd21158,32'd21229,32'd21300,32'd21371,32'd21442,32'd21513,32'd21584,32'd21655,32'd21726,32'd21797,32'd21868,32'd21939,32'd22010,32'd22081,32'd22152,32'd22223,32'd22294,32'd22365,32'd22436,32'd22507,32'd22578,32'd22649,32'd22720,32'd22791,32'd22862,32'd22933,32'd23004,32'd23075,32'd23146,32'd23217,32'd23288,32'd23359,32'd23430,32'd23501,32'd23572,32'd23643,32'd23714,32'd23785,32'd23856,32'd23927,32'd23998,32'd24069,32'd24140,32'd24211,32'd24282,32'd24353,32'd24424,32'd24495,32'd24566,32'd24637,32'd24708,32'd24779,32'd24850,32'd24921,32'd24992,32'd25063,32'd25134,32'd25205,32'd25276,32'd25347,32'd25418,32'd25489,32'd25560,32'd25631,32'd25702,32'd25773,32'd25844,32'd25915,32'd25986,32'd26057,32'd26128,32'd26199,32'd26270,32'd26341,32'd26412,32'd26483,32'd26554,32'd26625,32'd26696,32'd26767,32'd26838,32'd26909,32'd26980,32'd27051,32'd27122,32'd27193,32'd27264,32'd27335,32'd27406,32'd27477,32'd27548,32'd27619,32'd27690,32'd27761,32'd27832,32'd27903,32'd27974,32'd28045,32'd28116,32'd28187,32'd28258,32'd28329 };matrix[72]='{32'd0,32'd72,32'd144,32'd216,32'd288,32'd360,32'd432,32'd504,32'd576,32'd648,32'd720,32'd792,32'd864,32'd936,32'd1008,32'd1080,32'd1152,32'd1224,32'd1296,32'd1368,32'd1440,32'd1512,32'd1584,32'd1656,32'd1728,32'd1800,32'd1872,32'd1944,32'd2016,32'd2088,32'd2160,32'd2232,32'd2304,32'd2376,32'd2448,32'd2520,32'd2592,32'd2664,32'd2736,32'd2808,32'd2880,32'd2952,32'd3024,32'd3096,32'd3168,32'd3240,32'd3312,32'd3384,32'd3456,32'd3528,32'd3600,32'd3672,32'd3744,32'd3816,32'd3888,32'd3960,32'd4032,32'd4104,32'd4176,32'd4248,32'd4320,32'd4392,32'd4464,32'd4536,32'd4608,32'd4680,32'd4752,32'd4824,32'd4896,32'd4968,32'd5040,32'd5112,32'd5184,32'd5256,32'd5328,32'd5400,32'd5472,32'd5544,32'd5616,32'd5688,32'd5760,32'd5832,32'd5904,32'd5976,32'd6048,32'd6120,32'd6192,32'd6264,32'd6336,32'd6408,32'd6480,32'd6552,32'd6624,32'd6696,32'd6768,32'd6840,32'd6912,32'd6984,32'd7056,32'd7128,32'd7200,32'd7272,32'd7344,32'd7416,32'd7488,32'd7560,32'd7632,32'd7704,32'd7776,32'd7848,32'd7920,32'd7992,32'd8064,32'd8136,32'd8208,32'd8280,32'd8352,32'd8424,32'd8496,32'd8568,32'd8640,32'd8712,32'd8784,32'd8856,32'd8928,32'd9000,32'd9072,32'd9144,32'd9216,32'd9288,32'd9360,32'd9432,32'd9504,32'd9576,32'd9648,32'd9720,32'd9792,32'd9864,32'd9936,32'd10008,32'd10080,32'd10152,32'd10224,32'd10296,32'd10368,32'd10440,32'd10512,32'd10584,32'd10656,32'd10728,32'd10800,32'd10872,32'd10944,32'd11016,32'd11088,32'd11160,32'd11232,32'd11304,32'd11376,32'd11448,32'd11520,32'd11592,32'd11664,32'd11736,32'd11808,32'd11880,32'd11952,32'd12024,32'd12096,32'd12168,32'd12240,32'd12312,32'd12384,32'd12456,32'd12528,32'd12600,32'd12672,32'd12744,32'd12816,32'd12888,32'd12960,32'd13032,32'd13104,32'd13176,32'd13248,32'd13320,32'd13392,32'd13464,32'd13536,32'd13608,32'd13680,32'd13752,32'd13824,32'd13896,32'd13968,32'd14040,32'd14112,32'd14184,32'd14256,32'd14328,32'd14400,32'd14472,32'd14544,32'd14616,32'd14688,32'd14760,32'd14832,32'd14904,32'd14976,32'd15048,32'd15120,32'd15192,32'd15264,32'd15336,32'd15408,32'd15480,32'd15552,32'd15624,32'd15696,32'd15768,32'd15840,32'd15912,32'd15984,32'd16056,32'd16128,32'd16200,32'd16272,32'd16344,32'd16416,32'd16488,32'd16560,32'd16632,32'd16704,32'd16776,32'd16848,32'd16920,32'd16992,32'd17064,32'd17136,32'd17208,32'd17280,32'd17352,32'd17424,32'd17496,32'd17568,32'd17640,32'd17712,32'd17784,32'd17856,32'd17928,32'd18000,32'd18072,32'd18144,32'd18216,32'd18288,32'd18360,32'd18432,32'd18504,32'd18576,32'd18648,32'd18720,32'd18792,32'd18864,32'd18936,32'd19008,32'd19080,32'd19152,32'd19224,32'd19296,32'd19368,32'd19440,32'd19512,32'd19584,32'd19656,32'd19728,32'd19800,32'd19872,32'd19944,32'd20016,32'd20088,32'd20160,32'd20232,32'd20304,32'd20376,32'd20448,32'd20520,32'd20592,32'd20664,32'd20736,32'd20808,32'd20880,32'd20952,32'd21024,32'd21096,32'd21168,32'd21240,32'd21312,32'd21384,32'd21456,32'd21528,32'd21600,32'd21672,32'd21744,32'd21816,32'd21888,32'd21960,32'd22032,32'd22104,32'd22176,32'd22248,32'd22320,32'd22392,32'd22464,32'd22536,32'd22608,32'd22680,32'd22752,32'd22824,32'd22896,32'd22968,32'd23040,32'd23112,32'd23184,32'd23256,32'd23328,32'd23400,32'd23472,32'd23544,32'd23616,32'd23688,32'd23760,32'd23832,32'd23904,32'd23976,32'd24048,32'd24120,32'd24192,32'd24264,32'd24336,32'd24408,32'd24480,32'd24552,32'd24624,32'd24696,32'd24768,32'd24840,32'd24912,32'd24984,32'd25056,32'd25128,32'd25200,32'd25272,32'd25344,32'd25416,32'd25488,32'd25560,32'd25632,32'd25704,32'd25776,32'd25848,32'd25920,32'd25992,32'd26064,32'd26136,32'd26208,32'd26280,32'd26352,32'd26424,32'd26496,32'd26568,32'd26640,32'd26712,32'd26784,32'd26856,32'd26928,32'd27000,32'd27072,32'd27144,32'd27216,32'd27288,32'd27360,32'd27432,32'd27504,32'd27576,32'd27648,32'd27720,32'd27792,32'd27864,32'd27936,32'd28008,32'd28080,32'd28152,32'd28224,32'd28296,32'd28368,32'd28440,32'd28512,32'd28584,32'd28656,32'd28728 };matrix[73]='{32'd0,32'd73,32'd146,32'd219,32'd292,32'd365,32'd438,32'd511,32'd584,32'd657,32'd730,32'd803,32'd876,32'd949,32'd1022,32'd1095,32'd1168,32'd1241,32'd1314,32'd1387,32'd1460,32'd1533,32'd1606,32'd1679,32'd1752,32'd1825,32'd1898,32'd1971,32'd2044,32'd2117,32'd2190,32'd2263,32'd2336,32'd2409,32'd2482,32'd2555,32'd2628,32'd2701,32'd2774,32'd2847,32'd2920,32'd2993,32'd3066,32'd3139,32'd3212,32'd3285,32'd3358,32'd3431,32'd3504,32'd3577,32'd3650,32'd3723,32'd3796,32'd3869,32'd3942,32'd4015,32'd4088,32'd4161,32'd4234,32'd4307,32'd4380,32'd4453,32'd4526,32'd4599,32'd4672,32'd4745,32'd4818,32'd4891,32'd4964,32'd5037,32'd5110,32'd5183,32'd5256,32'd5329,32'd5402,32'd5475,32'd5548,32'd5621,32'd5694,32'd5767,32'd5840,32'd5913,32'd5986,32'd6059,32'd6132,32'd6205,32'd6278,32'd6351,32'd6424,32'd6497,32'd6570,32'd6643,32'd6716,32'd6789,32'd6862,32'd6935,32'd7008,32'd7081,32'd7154,32'd7227,32'd7300,32'd7373,32'd7446,32'd7519,32'd7592,32'd7665,32'd7738,32'd7811,32'd7884,32'd7957,32'd8030,32'd8103,32'd8176,32'd8249,32'd8322,32'd8395,32'd8468,32'd8541,32'd8614,32'd8687,32'd8760,32'd8833,32'd8906,32'd8979,32'd9052,32'd9125,32'd9198,32'd9271,32'd9344,32'd9417,32'd9490,32'd9563,32'd9636,32'd9709,32'd9782,32'd9855,32'd9928,32'd10001,32'd10074,32'd10147,32'd10220,32'd10293,32'd10366,32'd10439,32'd10512,32'd10585,32'd10658,32'd10731,32'd10804,32'd10877,32'd10950,32'd11023,32'd11096,32'd11169,32'd11242,32'd11315,32'd11388,32'd11461,32'd11534,32'd11607,32'd11680,32'd11753,32'd11826,32'd11899,32'd11972,32'd12045,32'd12118,32'd12191,32'd12264,32'd12337,32'd12410,32'd12483,32'd12556,32'd12629,32'd12702,32'd12775,32'd12848,32'd12921,32'd12994,32'd13067,32'd13140,32'd13213,32'd13286,32'd13359,32'd13432,32'd13505,32'd13578,32'd13651,32'd13724,32'd13797,32'd13870,32'd13943,32'd14016,32'd14089,32'd14162,32'd14235,32'd14308,32'd14381,32'd14454,32'd14527,32'd14600,32'd14673,32'd14746,32'd14819,32'd14892,32'd14965,32'd15038,32'd15111,32'd15184,32'd15257,32'd15330,32'd15403,32'd15476,32'd15549,32'd15622,32'd15695,32'd15768,32'd15841,32'd15914,32'd15987,32'd16060,32'd16133,32'd16206,32'd16279,32'd16352,32'd16425,32'd16498,32'd16571,32'd16644,32'd16717,32'd16790,32'd16863,32'd16936,32'd17009,32'd17082,32'd17155,32'd17228,32'd17301,32'd17374,32'd17447,32'd17520,32'd17593,32'd17666,32'd17739,32'd17812,32'd17885,32'd17958,32'd18031,32'd18104,32'd18177,32'd18250,32'd18323,32'd18396,32'd18469,32'd18542,32'd18615,32'd18688,32'd18761,32'd18834,32'd18907,32'd18980,32'd19053,32'd19126,32'd19199,32'd19272,32'd19345,32'd19418,32'd19491,32'd19564,32'd19637,32'd19710,32'd19783,32'd19856,32'd19929,32'd20002,32'd20075,32'd20148,32'd20221,32'd20294,32'd20367,32'd20440,32'd20513,32'd20586,32'd20659,32'd20732,32'd20805,32'd20878,32'd20951,32'd21024,32'd21097,32'd21170,32'd21243,32'd21316,32'd21389,32'd21462,32'd21535,32'd21608,32'd21681,32'd21754,32'd21827,32'd21900,32'd21973,32'd22046,32'd22119,32'd22192,32'd22265,32'd22338,32'd22411,32'd22484,32'd22557,32'd22630,32'd22703,32'd22776,32'd22849,32'd22922,32'd22995,32'd23068,32'd23141,32'd23214,32'd23287,32'd23360,32'd23433,32'd23506,32'd23579,32'd23652,32'd23725,32'd23798,32'd23871,32'd23944,32'd24017,32'd24090,32'd24163,32'd24236,32'd24309,32'd24382,32'd24455,32'd24528,32'd24601,32'd24674,32'd24747,32'd24820,32'd24893,32'd24966,32'd25039,32'd25112,32'd25185,32'd25258,32'd25331,32'd25404,32'd25477,32'd25550,32'd25623,32'd25696,32'd25769,32'd25842,32'd25915,32'd25988,32'd26061,32'd26134,32'd26207,32'd26280,32'd26353,32'd26426,32'd26499,32'd26572,32'd26645,32'd26718,32'd26791,32'd26864,32'd26937,32'd27010,32'd27083,32'd27156,32'd27229,32'd27302,32'd27375,32'd27448,32'd27521,32'd27594,32'd27667,32'd27740,32'd27813,32'd27886,32'd27959,32'd28032,32'd28105,32'd28178,32'd28251,32'd28324,32'd28397,32'd28470,32'd28543,32'd28616,32'd28689,32'd28762,32'd28835,32'd28908,32'd28981,32'd29054,32'd29127 };matrix[74]='{32'd0,32'd74,32'd148,32'd222,32'd296,32'd370,32'd444,32'd518,32'd592,32'd666,32'd740,32'd814,32'd888,32'd962,32'd1036,32'd1110,32'd1184,32'd1258,32'd1332,32'd1406,32'd1480,32'd1554,32'd1628,32'd1702,32'd1776,32'd1850,32'd1924,32'd1998,32'd2072,32'd2146,32'd2220,32'd2294,32'd2368,32'd2442,32'd2516,32'd2590,32'd2664,32'd2738,32'd2812,32'd2886,32'd2960,32'd3034,32'd3108,32'd3182,32'd3256,32'd3330,32'd3404,32'd3478,32'd3552,32'd3626,32'd3700,32'd3774,32'd3848,32'd3922,32'd3996,32'd4070,32'd4144,32'd4218,32'd4292,32'd4366,32'd4440,32'd4514,32'd4588,32'd4662,32'd4736,32'd4810,32'd4884,32'd4958,32'd5032,32'd5106,32'd5180,32'd5254,32'd5328,32'd5402,32'd5476,32'd5550,32'd5624,32'd5698,32'd5772,32'd5846,32'd5920,32'd5994,32'd6068,32'd6142,32'd6216,32'd6290,32'd6364,32'd6438,32'd6512,32'd6586,32'd6660,32'd6734,32'd6808,32'd6882,32'd6956,32'd7030,32'd7104,32'd7178,32'd7252,32'd7326,32'd7400,32'd7474,32'd7548,32'd7622,32'd7696,32'd7770,32'd7844,32'd7918,32'd7992,32'd8066,32'd8140,32'd8214,32'd8288,32'd8362,32'd8436,32'd8510,32'd8584,32'd8658,32'd8732,32'd8806,32'd8880,32'd8954,32'd9028,32'd9102,32'd9176,32'd9250,32'd9324,32'd9398,32'd9472,32'd9546,32'd9620,32'd9694,32'd9768,32'd9842,32'd9916,32'd9990,32'd10064,32'd10138,32'd10212,32'd10286,32'd10360,32'd10434,32'd10508,32'd10582,32'd10656,32'd10730,32'd10804,32'd10878,32'd10952,32'd11026,32'd11100,32'd11174,32'd11248,32'd11322,32'd11396,32'd11470,32'd11544,32'd11618,32'd11692,32'd11766,32'd11840,32'd11914,32'd11988,32'd12062,32'd12136,32'd12210,32'd12284,32'd12358,32'd12432,32'd12506,32'd12580,32'd12654,32'd12728,32'd12802,32'd12876,32'd12950,32'd13024,32'd13098,32'd13172,32'd13246,32'd13320,32'd13394,32'd13468,32'd13542,32'd13616,32'd13690,32'd13764,32'd13838,32'd13912,32'd13986,32'd14060,32'd14134,32'd14208,32'd14282,32'd14356,32'd14430,32'd14504,32'd14578,32'd14652,32'd14726,32'd14800,32'd14874,32'd14948,32'd15022,32'd15096,32'd15170,32'd15244,32'd15318,32'd15392,32'd15466,32'd15540,32'd15614,32'd15688,32'd15762,32'd15836,32'd15910,32'd15984,32'd16058,32'd16132,32'd16206,32'd16280,32'd16354,32'd16428,32'd16502,32'd16576,32'd16650,32'd16724,32'd16798,32'd16872,32'd16946,32'd17020,32'd17094,32'd17168,32'd17242,32'd17316,32'd17390,32'd17464,32'd17538,32'd17612,32'd17686,32'd17760,32'd17834,32'd17908,32'd17982,32'd18056,32'd18130,32'd18204,32'd18278,32'd18352,32'd18426,32'd18500,32'd18574,32'd18648,32'd18722,32'd18796,32'd18870,32'd18944,32'd19018,32'd19092,32'd19166,32'd19240,32'd19314,32'd19388,32'd19462,32'd19536,32'd19610,32'd19684,32'd19758,32'd19832,32'd19906,32'd19980,32'd20054,32'd20128,32'd20202,32'd20276,32'd20350,32'd20424,32'd20498,32'd20572,32'd20646,32'd20720,32'd20794,32'd20868,32'd20942,32'd21016,32'd21090,32'd21164,32'd21238,32'd21312,32'd21386,32'd21460,32'd21534,32'd21608,32'd21682,32'd21756,32'd21830,32'd21904,32'd21978,32'd22052,32'd22126,32'd22200,32'd22274,32'd22348,32'd22422,32'd22496,32'd22570,32'd22644,32'd22718,32'd22792,32'd22866,32'd22940,32'd23014,32'd23088,32'd23162,32'd23236,32'd23310,32'd23384,32'd23458,32'd23532,32'd23606,32'd23680,32'd23754,32'd23828,32'd23902,32'd23976,32'd24050,32'd24124,32'd24198,32'd24272,32'd24346,32'd24420,32'd24494,32'd24568,32'd24642,32'd24716,32'd24790,32'd24864,32'd24938,32'd25012,32'd25086,32'd25160,32'd25234,32'd25308,32'd25382,32'd25456,32'd25530,32'd25604,32'd25678,32'd25752,32'd25826,32'd25900,32'd25974,32'd26048,32'd26122,32'd26196,32'd26270,32'd26344,32'd26418,32'd26492,32'd26566,32'd26640,32'd26714,32'd26788,32'd26862,32'd26936,32'd27010,32'd27084,32'd27158,32'd27232,32'd27306,32'd27380,32'd27454,32'd27528,32'd27602,32'd27676,32'd27750,32'd27824,32'd27898,32'd27972,32'd28046,32'd28120,32'd28194,32'd28268,32'd28342,32'd28416,32'd28490,32'd28564,32'd28638,32'd28712,32'd28786,32'd28860,32'd28934,32'd29008,32'd29082,32'd29156,32'd29230,32'd29304,32'd29378,32'd29452,32'd29526 };matrix[75]='{32'd0,32'd75,32'd150,32'd225,32'd300,32'd375,32'd450,32'd525,32'd600,32'd675,32'd750,32'd825,32'd900,32'd975,32'd1050,32'd1125,32'd1200,32'd1275,32'd1350,32'd1425,32'd1500,32'd1575,32'd1650,32'd1725,32'd1800,32'd1875,32'd1950,32'd2025,32'd2100,32'd2175,32'd2250,32'd2325,32'd2400,32'd2475,32'd2550,32'd2625,32'd2700,32'd2775,32'd2850,32'd2925,32'd3000,32'd3075,32'd3150,32'd3225,32'd3300,32'd3375,32'd3450,32'd3525,32'd3600,32'd3675,32'd3750,32'd3825,32'd3900,32'd3975,32'd4050,32'd4125,32'd4200,32'd4275,32'd4350,32'd4425,32'd4500,32'd4575,32'd4650,32'd4725,32'd4800,32'd4875,32'd4950,32'd5025,32'd5100,32'd5175,32'd5250,32'd5325,32'd5400,32'd5475,32'd5550,32'd5625,32'd5700,32'd5775,32'd5850,32'd5925,32'd6000,32'd6075,32'd6150,32'd6225,32'd6300,32'd6375,32'd6450,32'd6525,32'd6600,32'd6675,32'd6750,32'd6825,32'd6900,32'd6975,32'd7050,32'd7125,32'd7200,32'd7275,32'd7350,32'd7425,32'd7500,32'd7575,32'd7650,32'd7725,32'd7800,32'd7875,32'd7950,32'd8025,32'd8100,32'd8175,32'd8250,32'd8325,32'd8400,32'd8475,32'd8550,32'd8625,32'd8700,32'd8775,32'd8850,32'd8925,32'd9000,32'd9075,32'd9150,32'd9225,32'd9300,32'd9375,32'd9450,32'd9525,32'd9600,32'd9675,32'd9750,32'd9825,32'd9900,32'd9975,32'd10050,32'd10125,32'd10200,32'd10275,32'd10350,32'd10425,32'd10500,32'd10575,32'd10650,32'd10725,32'd10800,32'd10875,32'd10950,32'd11025,32'd11100,32'd11175,32'd11250,32'd11325,32'd11400,32'd11475,32'd11550,32'd11625,32'd11700,32'd11775,32'd11850,32'd11925,32'd12000,32'd12075,32'd12150,32'd12225,32'd12300,32'd12375,32'd12450,32'd12525,32'd12600,32'd12675,32'd12750,32'd12825,32'd12900,32'd12975,32'd13050,32'd13125,32'd13200,32'd13275,32'd13350,32'd13425,32'd13500,32'd13575,32'd13650,32'd13725,32'd13800,32'd13875,32'd13950,32'd14025,32'd14100,32'd14175,32'd14250,32'd14325,32'd14400,32'd14475,32'd14550,32'd14625,32'd14700,32'd14775,32'd14850,32'd14925,32'd15000,32'd15075,32'd15150,32'd15225,32'd15300,32'd15375,32'd15450,32'd15525,32'd15600,32'd15675,32'd15750,32'd15825,32'd15900,32'd15975,32'd16050,32'd16125,32'd16200,32'd16275,32'd16350,32'd16425,32'd16500,32'd16575,32'd16650,32'd16725,32'd16800,32'd16875,32'd16950,32'd17025,32'd17100,32'd17175,32'd17250,32'd17325,32'd17400,32'd17475,32'd17550,32'd17625,32'd17700,32'd17775,32'd17850,32'd17925,32'd18000,32'd18075,32'd18150,32'd18225,32'd18300,32'd18375,32'd18450,32'd18525,32'd18600,32'd18675,32'd18750,32'd18825,32'd18900,32'd18975,32'd19050,32'd19125,32'd19200,32'd19275,32'd19350,32'd19425,32'd19500,32'd19575,32'd19650,32'd19725,32'd19800,32'd19875,32'd19950,32'd20025,32'd20100,32'd20175,32'd20250,32'd20325,32'd20400,32'd20475,32'd20550,32'd20625,32'd20700,32'd20775,32'd20850,32'd20925,32'd21000,32'd21075,32'd21150,32'd21225,32'd21300,32'd21375,32'd21450,32'd21525,32'd21600,32'd21675,32'd21750,32'd21825,32'd21900,32'd21975,32'd22050,32'd22125,32'd22200,32'd22275,32'd22350,32'd22425,32'd22500,32'd22575,32'd22650,32'd22725,32'd22800,32'd22875,32'd22950,32'd23025,32'd23100,32'd23175,32'd23250,32'd23325,32'd23400,32'd23475,32'd23550,32'd23625,32'd23700,32'd23775,32'd23850,32'd23925,32'd24000,32'd24075,32'd24150,32'd24225,32'd24300,32'd24375,32'd24450,32'd24525,32'd24600,32'd24675,32'd24750,32'd24825,32'd24900,32'd24975,32'd25050,32'd25125,32'd25200,32'd25275,32'd25350,32'd25425,32'd25500,32'd25575,32'd25650,32'd25725,32'd25800,32'd25875,32'd25950,32'd26025,32'd26100,32'd26175,32'd26250,32'd26325,32'd26400,32'd26475,32'd26550,32'd26625,32'd26700,32'd26775,32'd26850,32'd26925,32'd27000,32'd27075,32'd27150,32'd27225,32'd27300,32'd27375,32'd27450,32'd27525,32'd27600,32'd27675,32'd27750,32'd27825,32'd27900,32'd27975,32'd28050,32'd28125,32'd28200,32'd28275,32'd28350,32'd28425,32'd28500,32'd28575,32'd28650,32'd28725,32'd28800,32'd28875,32'd28950,32'd29025,32'd29100,32'd29175,32'd29250,32'd29325,32'd29400,32'd29475,32'd29550,32'd29625,32'd29700,32'd29775,32'd29850,32'd29925 };matrix[76]='{32'd0,32'd76,32'd152,32'd228,32'd304,32'd380,32'd456,32'd532,32'd608,32'd684,32'd760,32'd836,32'd912,32'd988,32'd1064,32'd1140,32'd1216,32'd1292,32'd1368,32'd1444,32'd1520,32'd1596,32'd1672,32'd1748,32'd1824,32'd1900,32'd1976,32'd2052,32'd2128,32'd2204,32'd2280,32'd2356,32'd2432,32'd2508,32'd2584,32'd2660,32'd2736,32'd2812,32'd2888,32'd2964,32'd3040,32'd3116,32'd3192,32'd3268,32'd3344,32'd3420,32'd3496,32'd3572,32'd3648,32'd3724,32'd3800,32'd3876,32'd3952,32'd4028,32'd4104,32'd4180,32'd4256,32'd4332,32'd4408,32'd4484,32'd4560,32'd4636,32'd4712,32'd4788,32'd4864,32'd4940,32'd5016,32'd5092,32'd5168,32'd5244,32'd5320,32'd5396,32'd5472,32'd5548,32'd5624,32'd5700,32'd5776,32'd5852,32'd5928,32'd6004,32'd6080,32'd6156,32'd6232,32'd6308,32'd6384,32'd6460,32'd6536,32'd6612,32'd6688,32'd6764,32'd6840,32'd6916,32'd6992,32'd7068,32'd7144,32'd7220,32'd7296,32'd7372,32'd7448,32'd7524,32'd7600,32'd7676,32'd7752,32'd7828,32'd7904,32'd7980,32'd8056,32'd8132,32'd8208,32'd8284,32'd8360,32'd8436,32'd8512,32'd8588,32'd8664,32'd8740,32'd8816,32'd8892,32'd8968,32'd9044,32'd9120,32'd9196,32'd9272,32'd9348,32'd9424,32'd9500,32'd9576,32'd9652,32'd9728,32'd9804,32'd9880,32'd9956,32'd10032,32'd10108,32'd10184,32'd10260,32'd10336,32'd10412,32'd10488,32'd10564,32'd10640,32'd10716,32'd10792,32'd10868,32'd10944,32'd11020,32'd11096,32'd11172,32'd11248,32'd11324,32'd11400,32'd11476,32'd11552,32'd11628,32'd11704,32'd11780,32'd11856,32'd11932,32'd12008,32'd12084,32'd12160,32'd12236,32'd12312,32'd12388,32'd12464,32'd12540,32'd12616,32'd12692,32'd12768,32'd12844,32'd12920,32'd12996,32'd13072,32'd13148,32'd13224,32'd13300,32'd13376,32'd13452,32'd13528,32'd13604,32'd13680,32'd13756,32'd13832,32'd13908,32'd13984,32'd14060,32'd14136,32'd14212,32'd14288,32'd14364,32'd14440,32'd14516,32'd14592,32'd14668,32'd14744,32'd14820,32'd14896,32'd14972,32'd15048,32'd15124,32'd15200,32'd15276,32'd15352,32'd15428,32'd15504,32'd15580,32'd15656,32'd15732,32'd15808,32'd15884,32'd15960,32'd16036,32'd16112,32'd16188,32'd16264,32'd16340,32'd16416,32'd16492,32'd16568,32'd16644,32'd16720,32'd16796,32'd16872,32'd16948,32'd17024,32'd17100,32'd17176,32'd17252,32'd17328,32'd17404,32'd17480,32'd17556,32'd17632,32'd17708,32'd17784,32'd17860,32'd17936,32'd18012,32'd18088,32'd18164,32'd18240,32'd18316,32'd18392,32'd18468,32'd18544,32'd18620,32'd18696,32'd18772,32'd18848,32'd18924,32'd19000,32'd19076,32'd19152,32'd19228,32'd19304,32'd19380,32'd19456,32'd19532,32'd19608,32'd19684,32'd19760,32'd19836,32'd19912,32'd19988,32'd20064,32'd20140,32'd20216,32'd20292,32'd20368,32'd20444,32'd20520,32'd20596,32'd20672,32'd20748,32'd20824,32'd20900,32'd20976,32'd21052,32'd21128,32'd21204,32'd21280,32'd21356,32'd21432,32'd21508,32'd21584,32'd21660,32'd21736,32'd21812,32'd21888,32'd21964,32'd22040,32'd22116,32'd22192,32'd22268,32'd22344,32'd22420,32'd22496,32'd22572,32'd22648,32'd22724,32'd22800,32'd22876,32'd22952,32'd23028,32'd23104,32'd23180,32'd23256,32'd23332,32'd23408,32'd23484,32'd23560,32'd23636,32'd23712,32'd23788,32'd23864,32'd23940,32'd24016,32'd24092,32'd24168,32'd24244,32'd24320,32'd24396,32'd24472,32'd24548,32'd24624,32'd24700,32'd24776,32'd24852,32'd24928,32'd25004,32'd25080,32'd25156,32'd25232,32'd25308,32'd25384,32'd25460,32'd25536,32'd25612,32'd25688,32'd25764,32'd25840,32'd25916,32'd25992,32'd26068,32'd26144,32'd26220,32'd26296,32'd26372,32'd26448,32'd26524,32'd26600,32'd26676,32'd26752,32'd26828,32'd26904,32'd26980,32'd27056,32'd27132,32'd27208,32'd27284,32'd27360,32'd27436,32'd27512,32'd27588,32'd27664,32'd27740,32'd27816,32'd27892,32'd27968,32'd28044,32'd28120,32'd28196,32'd28272,32'd28348,32'd28424,32'd28500,32'd28576,32'd28652,32'd28728,32'd28804,32'd28880,32'd28956,32'd29032,32'd29108,32'd29184,32'd29260,32'd29336,32'd29412,32'd29488,32'd29564,32'd29640,32'd29716,32'd29792,32'd29868,32'd29944,32'd30020,32'd30096,32'd30172,32'd30248,32'd30324 };matrix[77]='{32'd0,32'd77,32'd154,32'd231,32'd308,32'd385,32'd462,32'd539,32'd616,32'd693,32'd770,32'd847,32'd924,32'd1001,32'd1078,32'd1155,32'd1232,32'd1309,32'd1386,32'd1463,32'd1540,32'd1617,32'd1694,32'd1771,32'd1848,32'd1925,32'd2002,32'd2079,32'd2156,32'd2233,32'd2310,32'd2387,32'd2464,32'd2541,32'd2618,32'd2695,32'd2772,32'd2849,32'd2926,32'd3003,32'd3080,32'd3157,32'd3234,32'd3311,32'd3388,32'd3465,32'd3542,32'd3619,32'd3696,32'd3773,32'd3850,32'd3927,32'd4004,32'd4081,32'd4158,32'd4235,32'd4312,32'd4389,32'd4466,32'd4543,32'd4620,32'd4697,32'd4774,32'd4851,32'd4928,32'd5005,32'd5082,32'd5159,32'd5236,32'd5313,32'd5390,32'd5467,32'd5544,32'd5621,32'd5698,32'd5775,32'd5852,32'd5929,32'd6006,32'd6083,32'd6160,32'd6237,32'd6314,32'd6391,32'd6468,32'd6545,32'd6622,32'd6699,32'd6776,32'd6853,32'd6930,32'd7007,32'd7084,32'd7161,32'd7238,32'd7315,32'd7392,32'd7469,32'd7546,32'd7623,32'd7700,32'd7777,32'd7854,32'd7931,32'd8008,32'd8085,32'd8162,32'd8239,32'd8316,32'd8393,32'd8470,32'd8547,32'd8624,32'd8701,32'd8778,32'd8855,32'd8932,32'd9009,32'd9086,32'd9163,32'd9240,32'd9317,32'd9394,32'd9471,32'd9548,32'd9625,32'd9702,32'd9779,32'd9856,32'd9933,32'd10010,32'd10087,32'd10164,32'd10241,32'd10318,32'd10395,32'd10472,32'd10549,32'd10626,32'd10703,32'd10780,32'd10857,32'd10934,32'd11011,32'd11088,32'd11165,32'd11242,32'd11319,32'd11396,32'd11473,32'd11550,32'd11627,32'd11704,32'd11781,32'd11858,32'd11935,32'd12012,32'd12089,32'd12166,32'd12243,32'd12320,32'd12397,32'd12474,32'd12551,32'd12628,32'd12705,32'd12782,32'd12859,32'd12936,32'd13013,32'd13090,32'd13167,32'd13244,32'd13321,32'd13398,32'd13475,32'd13552,32'd13629,32'd13706,32'd13783,32'd13860,32'd13937,32'd14014,32'd14091,32'd14168,32'd14245,32'd14322,32'd14399,32'd14476,32'd14553,32'd14630,32'd14707,32'd14784,32'd14861,32'd14938,32'd15015,32'd15092,32'd15169,32'd15246,32'd15323,32'd15400,32'd15477,32'd15554,32'd15631,32'd15708,32'd15785,32'd15862,32'd15939,32'd16016,32'd16093,32'd16170,32'd16247,32'd16324,32'd16401,32'd16478,32'd16555,32'd16632,32'd16709,32'd16786,32'd16863,32'd16940,32'd17017,32'd17094,32'd17171,32'd17248,32'd17325,32'd17402,32'd17479,32'd17556,32'd17633,32'd17710,32'd17787,32'd17864,32'd17941,32'd18018,32'd18095,32'd18172,32'd18249,32'd18326,32'd18403,32'd18480,32'd18557,32'd18634,32'd18711,32'd18788,32'd18865,32'd18942,32'd19019,32'd19096,32'd19173,32'd19250,32'd19327,32'd19404,32'd19481,32'd19558,32'd19635,32'd19712,32'd19789,32'd19866,32'd19943,32'd20020,32'd20097,32'd20174,32'd20251,32'd20328,32'd20405,32'd20482,32'd20559,32'd20636,32'd20713,32'd20790,32'd20867,32'd20944,32'd21021,32'd21098,32'd21175,32'd21252,32'd21329,32'd21406,32'd21483,32'd21560,32'd21637,32'd21714,32'd21791,32'd21868,32'd21945,32'd22022,32'd22099,32'd22176,32'd22253,32'd22330,32'd22407,32'd22484,32'd22561,32'd22638,32'd22715,32'd22792,32'd22869,32'd22946,32'd23023,32'd23100,32'd23177,32'd23254,32'd23331,32'd23408,32'd23485,32'd23562,32'd23639,32'd23716,32'd23793,32'd23870,32'd23947,32'd24024,32'd24101,32'd24178,32'd24255,32'd24332,32'd24409,32'd24486,32'd24563,32'd24640,32'd24717,32'd24794,32'd24871,32'd24948,32'd25025,32'd25102,32'd25179,32'd25256,32'd25333,32'd25410,32'd25487,32'd25564,32'd25641,32'd25718,32'd25795,32'd25872,32'd25949,32'd26026,32'd26103,32'd26180,32'd26257,32'd26334,32'd26411,32'd26488,32'd26565,32'd26642,32'd26719,32'd26796,32'd26873,32'd26950,32'd27027,32'd27104,32'd27181,32'd27258,32'd27335,32'd27412,32'd27489,32'd27566,32'd27643,32'd27720,32'd27797,32'd27874,32'd27951,32'd28028,32'd28105,32'd28182,32'd28259,32'd28336,32'd28413,32'd28490,32'd28567,32'd28644,32'd28721,32'd28798,32'd28875,32'd28952,32'd29029,32'd29106,32'd29183,32'd29260,32'd29337,32'd29414,32'd29491,32'd29568,32'd29645,32'd29722,32'd29799,32'd29876,32'd29953,32'd30030,32'd30107,32'd30184,32'd30261,32'd30338,32'd30415,32'd30492,32'd30569,32'd30646,32'd30723 };matrix[78]='{32'd0,32'd78,32'd156,32'd234,32'd312,32'd390,32'd468,32'd546,32'd624,32'd702,32'd780,32'd858,32'd936,32'd1014,32'd1092,32'd1170,32'd1248,32'd1326,32'd1404,32'd1482,32'd1560,32'd1638,32'd1716,32'd1794,32'd1872,32'd1950,32'd2028,32'd2106,32'd2184,32'd2262,32'd2340,32'd2418,32'd2496,32'd2574,32'd2652,32'd2730,32'd2808,32'd2886,32'd2964,32'd3042,32'd3120,32'd3198,32'd3276,32'd3354,32'd3432,32'd3510,32'd3588,32'd3666,32'd3744,32'd3822,32'd3900,32'd3978,32'd4056,32'd4134,32'd4212,32'd4290,32'd4368,32'd4446,32'd4524,32'd4602,32'd4680,32'd4758,32'd4836,32'd4914,32'd4992,32'd5070,32'd5148,32'd5226,32'd5304,32'd5382,32'd5460,32'd5538,32'd5616,32'd5694,32'd5772,32'd5850,32'd5928,32'd6006,32'd6084,32'd6162,32'd6240,32'd6318,32'd6396,32'd6474,32'd6552,32'd6630,32'd6708,32'd6786,32'd6864,32'd6942,32'd7020,32'd7098,32'd7176,32'd7254,32'd7332,32'd7410,32'd7488,32'd7566,32'd7644,32'd7722,32'd7800,32'd7878,32'd7956,32'd8034,32'd8112,32'd8190,32'd8268,32'd8346,32'd8424,32'd8502,32'd8580,32'd8658,32'd8736,32'd8814,32'd8892,32'd8970,32'd9048,32'd9126,32'd9204,32'd9282,32'd9360,32'd9438,32'd9516,32'd9594,32'd9672,32'd9750,32'd9828,32'd9906,32'd9984,32'd10062,32'd10140,32'd10218,32'd10296,32'd10374,32'd10452,32'd10530,32'd10608,32'd10686,32'd10764,32'd10842,32'd10920,32'd10998,32'd11076,32'd11154,32'd11232,32'd11310,32'd11388,32'd11466,32'd11544,32'd11622,32'd11700,32'd11778,32'd11856,32'd11934,32'd12012,32'd12090,32'd12168,32'd12246,32'd12324,32'd12402,32'd12480,32'd12558,32'd12636,32'd12714,32'd12792,32'd12870,32'd12948,32'd13026,32'd13104,32'd13182,32'd13260,32'd13338,32'd13416,32'd13494,32'd13572,32'd13650,32'd13728,32'd13806,32'd13884,32'd13962,32'd14040,32'd14118,32'd14196,32'd14274,32'd14352,32'd14430,32'd14508,32'd14586,32'd14664,32'd14742,32'd14820,32'd14898,32'd14976,32'd15054,32'd15132,32'd15210,32'd15288,32'd15366,32'd15444,32'd15522,32'd15600,32'd15678,32'd15756,32'd15834,32'd15912,32'd15990,32'd16068,32'd16146,32'd16224,32'd16302,32'd16380,32'd16458,32'd16536,32'd16614,32'd16692,32'd16770,32'd16848,32'd16926,32'd17004,32'd17082,32'd17160,32'd17238,32'd17316,32'd17394,32'd17472,32'd17550,32'd17628,32'd17706,32'd17784,32'd17862,32'd17940,32'd18018,32'd18096,32'd18174,32'd18252,32'd18330,32'd18408,32'd18486,32'd18564,32'd18642,32'd18720,32'd18798,32'd18876,32'd18954,32'd19032,32'd19110,32'd19188,32'd19266,32'd19344,32'd19422,32'd19500,32'd19578,32'd19656,32'd19734,32'd19812,32'd19890,32'd19968,32'd20046,32'd20124,32'd20202,32'd20280,32'd20358,32'd20436,32'd20514,32'd20592,32'd20670,32'd20748,32'd20826,32'd20904,32'd20982,32'd21060,32'd21138,32'd21216,32'd21294,32'd21372,32'd21450,32'd21528,32'd21606,32'd21684,32'd21762,32'd21840,32'd21918,32'd21996,32'd22074,32'd22152,32'd22230,32'd22308,32'd22386,32'd22464,32'd22542,32'd22620,32'd22698,32'd22776,32'd22854,32'd22932,32'd23010,32'd23088,32'd23166,32'd23244,32'd23322,32'd23400,32'd23478,32'd23556,32'd23634,32'd23712,32'd23790,32'd23868,32'd23946,32'd24024,32'd24102,32'd24180,32'd24258,32'd24336,32'd24414,32'd24492,32'd24570,32'd24648,32'd24726,32'd24804,32'd24882,32'd24960,32'd25038,32'd25116,32'd25194,32'd25272,32'd25350,32'd25428,32'd25506,32'd25584,32'd25662,32'd25740,32'd25818,32'd25896,32'd25974,32'd26052,32'd26130,32'd26208,32'd26286,32'd26364,32'd26442,32'd26520,32'd26598,32'd26676,32'd26754,32'd26832,32'd26910,32'd26988,32'd27066,32'd27144,32'd27222,32'd27300,32'd27378,32'd27456,32'd27534,32'd27612,32'd27690,32'd27768,32'd27846,32'd27924,32'd28002,32'd28080,32'd28158,32'd28236,32'd28314,32'd28392,32'd28470,32'd28548,32'd28626,32'd28704,32'd28782,32'd28860,32'd28938,32'd29016,32'd29094,32'd29172,32'd29250,32'd29328,32'd29406,32'd29484,32'd29562,32'd29640,32'd29718,32'd29796,32'd29874,32'd29952,32'd30030,32'd30108,32'd30186,32'd30264,32'd30342,32'd30420,32'd30498,32'd30576,32'd30654,32'd30732,32'd30810,32'd30888,32'd30966,32'd31044,32'd31122 };matrix[79]='{32'd0,32'd79,32'd158,32'd237,32'd316,32'd395,32'd474,32'd553,32'd632,32'd711,32'd790,32'd869,32'd948,32'd1027,32'd1106,32'd1185,32'd1264,32'd1343,32'd1422,32'd1501,32'd1580,32'd1659,32'd1738,32'd1817,32'd1896,32'd1975,32'd2054,32'd2133,32'd2212,32'd2291,32'd2370,32'd2449,32'd2528,32'd2607,32'd2686,32'd2765,32'd2844,32'd2923,32'd3002,32'd3081,32'd3160,32'd3239,32'd3318,32'd3397,32'd3476,32'd3555,32'd3634,32'd3713,32'd3792,32'd3871,32'd3950,32'd4029,32'd4108,32'd4187,32'd4266,32'd4345,32'd4424,32'd4503,32'd4582,32'd4661,32'd4740,32'd4819,32'd4898,32'd4977,32'd5056,32'd5135,32'd5214,32'd5293,32'd5372,32'd5451,32'd5530,32'd5609,32'd5688,32'd5767,32'd5846,32'd5925,32'd6004,32'd6083,32'd6162,32'd6241,32'd6320,32'd6399,32'd6478,32'd6557,32'd6636,32'd6715,32'd6794,32'd6873,32'd6952,32'd7031,32'd7110,32'd7189,32'd7268,32'd7347,32'd7426,32'd7505,32'd7584,32'd7663,32'd7742,32'd7821,32'd7900,32'd7979,32'd8058,32'd8137,32'd8216,32'd8295,32'd8374,32'd8453,32'd8532,32'd8611,32'd8690,32'd8769,32'd8848,32'd8927,32'd9006,32'd9085,32'd9164,32'd9243,32'd9322,32'd9401,32'd9480,32'd9559,32'd9638,32'd9717,32'd9796,32'd9875,32'd9954,32'd10033,32'd10112,32'd10191,32'd10270,32'd10349,32'd10428,32'd10507,32'd10586,32'd10665,32'd10744,32'd10823,32'd10902,32'd10981,32'd11060,32'd11139,32'd11218,32'd11297,32'd11376,32'd11455,32'd11534,32'd11613,32'd11692,32'd11771,32'd11850,32'd11929,32'd12008,32'd12087,32'd12166,32'd12245,32'd12324,32'd12403,32'd12482,32'd12561,32'd12640,32'd12719,32'd12798,32'd12877,32'd12956,32'd13035,32'd13114,32'd13193,32'd13272,32'd13351,32'd13430,32'd13509,32'd13588,32'd13667,32'd13746,32'd13825,32'd13904,32'd13983,32'd14062,32'd14141,32'd14220,32'd14299,32'd14378,32'd14457,32'd14536,32'd14615,32'd14694,32'd14773,32'd14852,32'd14931,32'd15010,32'd15089,32'd15168,32'd15247,32'd15326,32'd15405,32'd15484,32'd15563,32'd15642,32'd15721,32'd15800,32'd15879,32'd15958,32'd16037,32'd16116,32'd16195,32'd16274,32'd16353,32'd16432,32'd16511,32'd16590,32'd16669,32'd16748,32'd16827,32'd16906,32'd16985,32'd17064,32'd17143,32'd17222,32'd17301,32'd17380,32'd17459,32'd17538,32'd17617,32'd17696,32'd17775,32'd17854,32'd17933,32'd18012,32'd18091,32'd18170,32'd18249,32'd18328,32'd18407,32'd18486,32'd18565,32'd18644,32'd18723,32'd18802,32'd18881,32'd18960,32'd19039,32'd19118,32'd19197,32'd19276,32'd19355,32'd19434,32'd19513,32'd19592,32'd19671,32'd19750,32'd19829,32'd19908,32'd19987,32'd20066,32'd20145,32'd20224,32'd20303,32'd20382,32'd20461,32'd20540,32'd20619,32'd20698,32'd20777,32'd20856,32'd20935,32'd21014,32'd21093,32'd21172,32'd21251,32'd21330,32'd21409,32'd21488,32'd21567,32'd21646,32'd21725,32'd21804,32'd21883,32'd21962,32'd22041,32'd22120,32'd22199,32'd22278,32'd22357,32'd22436,32'd22515,32'd22594,32'd22673,32'd22752,32'd22831,32'd22910,32'd22989,32'd23068,32'd23147,32'd23226,32'd23305,32'd23384,32'd23463,32'd23542,32'd23621,32'd23700,32'd23779,32'd23858,32'd23937,32'd24016,32'd24095,32'd24174,32'd24253,32'd24332,32'd24411,32'd24490,32'd24569,32'd24648,32'd24727,32'd24806,32'd24885,32'd24964,32'd25043,32'd25122,32'd25201,32'd25280,32'd25359,32'd25438,32'd25517,32'd25596,32'd25675,32'd25754,32'd25833,32'd25912,32'd25991,32'd26070,32'd26149,32'd26228,32'd26307,32'd26386,32'd26465,32'd26544,32'd26623,32'd26702,32'd26781,32'd26860,32'd26939,32'd27018,32'd27097,32'd27176,32'd27255,32'd27334,32'd27413,32'd27492,32'd27571,32'd27650,32'd27729,32'd27808,32'd27887,32'd27966,32'd28045,32'd28124,32'd28203,32'd28282,32'd28361,32'd28440,32'd28519,32'd28598,32'd28677,32'd28756,32'd28835,32'd28914,32'd28993,32'd29072,32'd29151,32'd29230,32'd29309,32'd29388,32'd29467,32'd29546,32'd29625,32'd29704,32'd29783,32'd29862,32'd29941,32'd30020,32'd30099,32'd30178,32'd30257,32'd30336,32'd30415,32'd30494,32'd30573,32'd30652,32'd30731,32'd30810,32'd30889,32'd30968,32'd31047,32'd31126,32'd31205,32'd31284,32'd31363,32'd31442,32'd31521 };matrix[80]='{32'd0,32'd80,32'd160,32'd240,32'd320,32'd400,32'd480,32'd560,32'd640,32'd720,32'd800,32'd880,32'd960,32'd1040,32'd1120,32'd1200,32'd1280,32'd1360,32'd1440,32'd1520,32'd1600,32'd1680,32'd1760,32'd1840,32'd1920,32'd2000,32'd2080,32'd2160,32'd2240,32'd2320,32'd2400,32'd2480,32'd2560,32'd2640,32'd2720,32'd2800,32'd2880,32'd2960,32'd3040,32'd3120,32'd3200,32'd3280,32'd3360,32'd3440,32'd3520,32'd3600,32'd3680,32'd3760,32'd3840,32'd3920,32'd4000,32'd4080,32'd4160,32'd4240,32'd4320,32'd4400,32'd4480,32'd4560,32'd4640,32'd4720,32'd4800,32'd4880,32'd4960,32'd5040,32'd5120,32'd5200,32'd5280,32'd5360,32'd5440,32'd5520,32'd5600,32'd5680,32'd5760,32'd5840,32'd5920,32'd6000,32'd6080,32'd6160,32'd6240,32'd6320,32'd6400,32'd6480,32'd6560,32'd6640,32'd6720,32'd6800,32'd6880,32'd6960,32'd7040,32'd7120,32'd7200,32'd7280,32'd7360,32'd7440,32'd7520,32'd7600,32'd7680,32'd7760,32'd7840,32'd7920,32'd8000,32'd8080,32'd8160,32'd8240,32'd8320,32'd8400,32'd8480,32'd8560,32'd8640,32'd8720,32'd8800,32'd8880,32'd8960,32'd9040,32'd9120,32'd9200,32'd9280,32'd9360,32'd9440,32'd9520,32'd9600,32'd9680,32'd9760,32'd9840,32'd9920,32'd10000,32'd10080,32'd10160,32'd10240,32'd10320,32'd10400,32'd10480,32'd10560,32'd10640,32'd10720,32'd10800,32'd10880,32'd10960,32'd11040,32'd11120,32'd11200,32'd11280,32'd11360,32'd11440,32'd11520,32'd11600,32'd11680,32'd11760,32'd11840,32'd11920,32'd12000,32'd12080,32'd12160,32'd12240,32'd12320,32'd12400,32'd12480,32'd12560,32'd12640,32'd12720,32'd12800,32'd12880,32'd12960,32'd13040,32'd13120,32'd13200,32'd13280,32'd13360,32'd13440,32'd13520,32'd13600,32'd13680,32'd13760,32'd13840,32'd13920,32'd14000,32'd14080,32'd14160,32'd14240,32'd14320,32'd14400,32'd14480,32'd14560,32'd14640,32'd14720,32'd14800,32'd14880,32'd14960,32'd15040,32'd15120,32'd15200,32'd15280,32'd15360,32'd15440,32'd15520,32'd15600,32'd15680,32'd15760,32'd15840,32'd15920,32'd16000,32'd16080,32'd16160,32'd16240,32'd16320,32'd16400,32'd16480,32'd16560,32'd16640,32'd16720,32'd16800,32'd16880,32'd16960,32'd17040,32'd17120,32'd17200,32'd17280,32'd17360,32'd17440,32'd17520,32'd17600,32'd17680,32'd17760,32'd17840,32'd17920,32'd18000,32'd18080,32'd18160,32'd18240,32'd18320,32'd18400,32'd18480,32'd18560,32'd18640,32'd18720,32'd18800,32'd18880,32'd18960,32'd19040,32'd19120,32'd19200,32'd19280,32'd19360,32'd19440,32'd19520,32'd19600,32'd19680,32'd19760,32'd19840,32'd19920,32'd20000,32'd20080,32'd20160,32'd20240,32'd20320,32'd20400,32'd20480,32'd20560,32'd20640,32'd20720,32'd20800,32'd20880,32'd20960,32'd21040,32'd21120,32'd21200,32'd21280,32'd21360,32'd21440,32'd21520,32'd21600,32'd21680,32'd21760,32'd21840,32'd21920,32'd22000,32'd22080,32'd22160,32'd22240,32'd22320,32'd22400,32'd22480,32'd22560,32'd22640,32'd22720,32'd22800,32'd22880,32'd22960,32'd23040,32'd23120,32'd23200,32'd23280,32'd23360,32'd23440,32'd23520,32'd23600,32'd23680,32'd23760,32'd23840,32'd23920,32'd24000,32'd24080,32'd24160,32'd24240,32'd24320,32'd24400,32'd24480,32'd24560,32'd24640,32'd24720,32'd24800,32'd24880,32'd24960,32'd25040,32'd25120,32'd25200,32'd25280,32'd25360,32'd25440,32'd25520,32'd25600,32'd25680,32'd25760,32'd25840,32'd25920,32'd26000,32'd26080,32'd26160,32'd26240,32'd26320,32'd26400,32'd26480,32'd26560,32'd26640,32'd26720,32'd26800,32'd26880,32'd26960,32'd27040,32'd27120,32'd27200,32'd27280,32'd27360,32'd27440,32'd27520,32'd27600,32'd27680,32'd27760,32'd27840,32'd27920,32'd28000,32'd28080,32'd28160,32'd28240,32'd28320,32'd28400,32'd28480,32'd28560,32'd28640,32'd28720,32'd28800,32'd28880,32'd28960,32'd29040,32'd29120,32'd29200,32'd29280,32'd29360,32'd29440,32'd29520,32'd29600,32'd29680,32'd29760,32'd29840,32'd29920,32'd30000,32'd30080,32'd30160,32'd30240,32'd30320,32'd30400,32'd30480,32'd30560,32'd30640,32'd30720,32'd30800,32'd30880,32'd30960,32'd31040,32'd31120,32'd31200,32'd31280,32'd31360,32'd31440,32'd31520,32'd31600,32'd31680,32'd31760,32'd31840,32'd31920 };matrix[81]='{32'd0,32'd81,32'd162,32'd243,32'd324,32'd405,32'd486,32'd567,32'd648,32'd729,32'd810,32'd891,32'd972,32'd1053,32'd1134,32'd1215,32'd1296,32'd1377,32'd1458,32'd1539,32'd1620,32'd1701,32'd1782,32'd1863,32'd1944,32'd2025,32'd2106,32'd2187,32'd2268,32'd2349,32'd2430,32'd2511,32'd2592,32'd2673,32'd2754,32'd2835,32'd2916,32'd2997,32'd3078,32'd3159,32'd3240,32'd3321,32'd3402,32'd3483,32'd3564,32'd3645,32'd3726,32'd3807,32'd3888,32'd3969,32'd4050,32'd4131,32'd4212,32'd4293,32'd4374,32'd4455,32'd4536,32'd4617,32'd4698,32'd4779,32'd4860,32'd4941,32'd5022,32'd5103,32'd5184,32'd5265,32'd5346,32'd5427,32'd5508,32'd5589,32'd5670,32'd5751,32'd5832,32'd5913,32'd5994,32'd6075,32'd6156,32'd6237,32'd6318,32'd6399,32'd6480,32'd6561,32'd6642,32'd6723,32'd6804,32'd6885,32'd6966,32'd7047,32'd7128,32'd7209,32'd7290,32'd7371,32'd7452,32'd7533,32'd7614,32'd7695,32'd7776,32'd7857,32'd7938,32'd8019,32'd8100,32'd8181,32'd8262,32'd8343,32'd8424,32'd8505,32'd8586,32'd8667,32'd8748,32'd8829,32'd8910,32'd8991,32'd9072,32'd9153,32'd9234,32'd9315,32'd9396,32'd9477,32'd9558,32'd9639,32'd9720,32'd9801,32'd9882,32'd9963,32'd10044,32'd10125,32'd10206,32'd10287,32'd10368,32'd10449,32'd10530,32'd10611,32'd10692,32'd10773,32'd10854,32'd10935,32'd11016,32'd11097,32'd11178,32'd11259,32'd11340,32'd11421,32'd11502,32'd11583,32'd11664,32'd11745,32'd11826,32'd11907,32'd11988,32'd12069,32'd12150,32'd12231,32'd12312,32'd12393,32'd12474,32'd12555,32'd12636,32'd12717,32'd12798,32'd12879,32'd12960,32'd13041,32'd13122,32'd13203,32'd13284,32'd13365,32'd13446,32'd13527,32'd13608,32'd13689,32'd13770,32'd13851,32'd13932,32'd14013,32'd14094,32'd14175,32'd14256,32'd14337,32'd14418,32'd14499,32'd14580,32'd14661,32'd14742,32'd14823,32'd14904,32'd14985,32'd15066,32'd15147,32'd15228,32'd15309,32'd15390,32'd15471,32'd15552,32'd15633,32'd15714,32'd15795,32'd15876,32'd15957,32'd16038,32'd16119,32'd16200,32'd16281,32'd16362,32'd16443,32'd16524,32'd16605,32'd16686,32'd16767,32'd16848,32'd16929,32'd17010,32'd17091,32'd17172,32'd17253,32'd17334,32'd17415,32'd17496,32'd17577,32'd17658,32'd17739,32'd17820,32'd17901,32'd17982,32'd18063,32'd18144,32'd18225,32'd18306,32'd18387,32'd18468,32'd18549,32'd18630,32'd18711,32'd18792,32'd18873,32'd18954,32'd19035,32'd19116,32'd19197,32'd19278,32'd19359,32'd19440,32'd19521,32'd19602,32'd19683,32'd19764,32'd19845,32'd19926,32'd20007,32'd20088,32'd20169,32'd20250,32'd20331,32'd20412,32'd20493,32'd20574,32'd20655,32'd20736,32'd20817,32'd20898,32'd20979,32'd21060,32'd21141,32'd21222,32'd21303,32'd21384,32'd21465,32'd21546,32'd21627,32'd21708,32'd21789,32'd21870,32'd21951,32'd22032,32'd22113,32'd22194,32'd22275,32'd22356,32'd22437,32'd22518,32'd22599,32'd22680,32'd22761,32'd22842,32'd22923,32'd23004,32'd23085,32'd23166,32'd23247,32'd23328,32'd23409,32'd23490,32'd23571,32'd23652,32'd23733,32'd23814,32'd23895,32'd23976,32'd24057,32'd24138,32'd24219,32'd24300,32'd24381,32'd24462,32'd24543,32'd24624,32'd24705,32'd24786,32'd24867,32'd24948,32'd25029,32'd25110,32'd25191,32'd25272,32'd25353,32'd25434,32'd25515,32'd25596,32'd25677,32'd25758,32'd25839,32'd25920,32'd26001,32'd26082,32'd26163,32'd26244,32'd26325,32'd26406,32'd26487,32'd26568,32'd26649,32'd26730,32'd26811,32'd26892,32'd26973,32'd27054,32'd27135,32'd27216,32'd27297,32'd27378,32'd27459,32'd27540,32'd27621,32'd27702,32'd27783,32'd27864,32'd27945,32'd28026,32'd28107,32'd28188,32'd28269,32'd28350,32'd28431,32'd28512,32'd28593,32'd28674,32'd28755,32'd28836,32'd28917,32'd28998,32'd29079,32'd29160,32'd29241,32'd29322,32'd29403,32'd29484,32'd29565,32'd29646,32'd29727,32'd29808,32'd29889,32'd29970,32'd30051,32'd30132,32'd30213,32'd30294,32'd30375,32'd30456,32'd30537,32'd30618,32'd30699,32'd30780,32'd30861,32'd30942,32'd31023,32'd31104,32'd31185,32'd31266,32'd31347,32'd31428,32'd31509,32'd31590,32'd31671,32'd31752,32'd31833,32'd31914,32'd31995,32'd32076,32'd32157,32'd32238,32'd32319 };matrix[82]='{32'd0,32'd82,32'd164,32'd246,32'd328,32'd410,32'd492,32'd574,32'd656,32'd738,32'd820,32'd902,32'd984,32'd1066,32'd1148,32'd1230,32'd1312,32'd1394,32'd1476,32'd1558,32'd1640,32'd1722,32'd1804,32'd1886,32'd1968,32'd2050,32'd2132,32'd2214,32'd2296,32'd2378,32'd2460,32'd2542,32'd2624,32'd2706,32'd2788,32'd2870,32'd2952,32'd3034,32'd3116,32'd3198,32'd3280,32'd3362,32'd3444,32'd3526,32'd3608,32'd3690,32'd3772,32'd3854,32'd3936,32'd4018,32'd4100,32'd4182,32'd4264,32'd4346,32'd4428,32'd4510,32'd4592,32'd4674,32'd4756,32'd4838,32'd4920,32'd5002,32'd5084,32'd5166,32'd5248,32'd5330,32'd5412,32'd5494,32'd5576,32'd5658,32'd5740,32'd5822,32'd5904,32'd5986,32'd6068,32'd6150,32'd6232,32'd6314,32'd6396,32'd6478,32'd6560,32'd6642,32'd6724,32'd6806,32'd6888,32'd6970,32'd7052,32'd7134,32'd7216,32'd7298,32'd7380,32'd7462,32'd7544,32'd7626,32'd7708,32'd7790,32'd7872,32'd7954,32'd8036,32'd8118,32'd8200,32'd8282,32'd8364,32'd8446,32'd8528,32'd8610,32'd8692,32'd8774,32'd8856,32'd8938,32'd9020,32'd9102,32'd9184,32'd9266,32'd9348,32'd9430,32'd9512,32'd9594,32'd9676,32'd9758,32'd9840,32'd9922,32'd10004,32'd10086,32'd10168,32'd10250,32'd10332,32'd10414,32'd10496,32'd10578,32'd10660,32'd10742,32'd10824,32'd10906,32'd10988,32'd11070,32'd11152,32'd11234,32'd11316,32'd11398,32'd11480,32'd11562,32'd11644,32'd11726,32'd11808,32'd11890,32'd11972,32'd12054,32'd12136,32'd12218,32'd12300,32'd12382,32'd12464,32'd12546,32'd12628,32'd12710,32'd12792,32'd12874,32'd12956,32'd13038,32'd13120,32'd13202,32'd13284,32'd13366,32'd13448,32'd13530,32'd13612,32'd13694,32'd13776,32'd13858,32'd13940,32'd14022,32'd14104,32'd14186,32'd14268,32'd14350,32'd14432,32'd14514,32'd14596,32'd14678,32'd14760,32'd14842,32'd14924,32'd15006,32'd15088,32'd15170,32'd15252,32'd15334,32'd15416,32'd15498,32'd15580,32'd15662,32'd15744,32'd15826,32'd15908,32'd15990,32'd16072,32'd16154,32'd16236,32'd16318,32'd16400,32'd16482,32'd16564,32'd16646,32'd16728,32'd16810,32'd16892,32'd16974,32'd17056,32'd17138,32'd17220,32'd17302,32'd17384,32'd17466,32'd17548,32'd17630,32'd17712,32'd17794,32'd17876,32'd17958,32'd18040,32'd18122,32'd18204,32'd18286,32'd18368,32'd18450,32'd18532,32'd18614,32'd18696,32'd18778,32'd18860,32'd18942,32'd19024,32'd19106,32'd19188,32'd19270,32'd19352,32'd19434,32'd19516,32'd19598,32'd19680,32'd19762,32'd19844,32'd19926,32'd20008,32'd20090,32'd20172,32'd20254,32'd20336,32'd20418,32'd20500,32'd20582,32'd20664,32'd20746,32'd20828,32'd20910,32'd20992,32'd21074,32'd21156,32'd21238,32'd21320,32'd21402,32'd21484,32'd21566,32'd21648,32'd21730,32'd21812,32'd21894,32'd21976,32'd22058,32'd22140,32'd22222,32'd22304,32'd22386,32'd22468,32'd22550,32'd22632,32'd22714,32'd22796,32'd22878,32'd22960,32'd23042,32'd23124,32'd23206,32'd23288,32'd23370,32'd23452,32'd23534,32'd23616,32'd23698,32'd23780,32'd23862,32'd23944,32'd24026,32'd24108,32'd24190,32'd24272,32'd24354,32'd24436,32'd24518,32'd24600,32'd24682,32'd24764,32'd24846,32'd24928,32'd25010,32'd25092,32'd25174,32'd25256,32'd25338,32'd25420,32'd25502,32'd25584,32'd25666,32'd25748,32'd25830,32'd25912,32'd25994,32'd26076,32'd26158,32'd26240,32'd26322,32'd26404,32'd26486,32'd26568,32'd26650,32'd26732,32'd26814,32'd26896,32'd26978,32'd27060,32'd27142,32'd27224,32'd27306,32'd27388,32'd27470,32'd27552,32'd27634,32'd27716,32'd27798,32'd27880,32'd27962,32'd28044,32'd28126,32'd28208,32'd28290,32'd28372,32'd28454,32'd28536,32'd28618,32'd28700,32'd28782,32'd28864,32'd28946,32'd29028,32'd29110,32'd29192,32'd29274,32'd29356,32'd29438,32'd29520,32'd29602,32'd29684,32'd29766,32'd29848,32'd29930,32'd30012,32'd30094,32'd30176,32'd30258,32'd30340,32'd30422,32'd30504,32'd30586,32'd30668,32'd30750,32'd30832,32'd30914,32'd30996,32'd31078,32'd31160,32'd31242,32'd31324,32'd31406,32'd31488,32'd31570,32'd31652,32'd31734,32'd31816,32'd31898,32'd31980,32'd32062,32'd32144,32'd32226,32'd32308,32'd32390,32'd32472,32'd32554,32'd32636,32'd32718 };matrix[83]='{32'd0,32'd83,32'd166,32'd249,32'd332,32'd415,32'd498,32'd581,32'd664,32'd747,32'd830,32'd913,32'd996,32'd1079,32'd1162,32'd1245,32'd1328,32'd1411,32'd1494,32'd1577,32'd1660,32'd1743,32'd1826,32'd1909,32'd1992,32'd2075,32'd2158,32'd2241,32'd2324,32'd2407,32'd2490,32'd2573,32'd2656,32'd2739,32'd2822,32'd2905,32'd2988,32'd3071,32'd3154,32'd3237,32'd3320,32'd3403,32'd3486,32'd3569,32'd3652,32'd3735,32'd3818,32'd3901,32'd3984,32'd4067,32'd4150,32'd4233,32'd4316,32'd4399,32'd4482,32'd4565,32'd4648,32'd4731,32'd4814,32'd4897,32'd4980,32'd5063,32'd5146,32'd5229,32'd5312,32'd5395,32'd5478,32'd5561,32'd5644,32'd5727,32'd5810,32'd5893,32'd5976,32'd6059,32'd6142,32'd6225,32'd6308,32'd6391,32'd6474,32'd6557,32'd6640,32'd6723,32'd6806,32'd6889,32'd6972,32'd7055,32'd7138,32'd7221,32'd7304,32'd7387,32'd7470,32'd7553,32'd7636,32'd7719,32'd7802,32'd7885,32'd7968,32'd8051,32'd8134,32'd8217,32'd8300,32'd8383,32'd8466,32'd8549,32'd8632,32'd8715,32'd8798,32'd8881,32'd8964,32'd9047,32'd9130,32'd9213,32'd9296,32'd9379,32'd9462,32'd9545,32'd9628,32'd9711,32'd9794,32'd9877,32'd9960,32'd10043,32'd10126,32'd10209,32'd10292,32'd10375,32'd10458,32'd10541,32'd10624,32'd10707,32'd10790,32'd10873,32'd10956,32'd11039,32'd11122,32'd11205,32'd11288,32'd11371,32'd11454,32'd11537,32'd11620,32'd11703,32'd11786,32'd11869,32'd11952,32'd12035,32'd12118,32'd12201,32'd12284,32'd12367,32'd12450,32'd12533,32'd12616,32'd12699,32'd12782,32'd12865,32'd12948,32'd13031,32'd13114,32'd13197,32'd13280,32'd13363,32'd13446,32'd13529,32'd13612,32'd13695,32'd13778,32'd13861,32'd13944,32'd14027,32'd14110,32'd14193,32'd14276,32'd14359,32'd14442,32'd14525,32'd14608,32'd14691,32'd14774,32'd14857,32'd14940,32'd15023,32'd15106,32'd15189,32'd15272,32'd15355,32'd15438,32'd15521,32'd15604,32'd15687,32'd15770,32'd15853,32'd15936,32'd16019,32'd16102,32'd16185,32'd16268,32'd16351,32'd16434,32'd16517,32'd16600,32'd16683,32'd16766,32'd16849,32'd16932,32'd17015,32'd17098,32'd17181,32'd17264,32'd17347,32'd17430,32'd17513,32'd17596,32'd17679,32'd17762,32'd17845,32'd17928,32'd18011,32'd18094,32'd18177,32'd18260,32'd18343,32'd18426,32'd18509,32'd18592,32'd18675,32'd18758,32'd18841,32'd18924,32'd19007,32'd19090,32'd19173,32'd19256,32'd19339,32'd19422,32'd19505,32'd19588,32'd19671,32'd19754,32'd19837,32'd19920,32'd20003,32'd20086,32'd20169,32'd20252,32'd20335,32'd20418,32'd20501,32'd20584,32'd20667,32'd20750,32'd20833,32'd20916,32'd20999,32'd21082,32'd21165,32'd21248,32'd21331,32'd21414,32'd21497,32'd21580,32'd21663,32'd21746,32'd21829,32'd21912,32'd21995,32'd22078,32'd22161,32'd22244,32'd22327,32'd22410,32'd22493,32'd22576,32'd22659,32'd22742,32'd22825,32'd22908,32'd22991,32'd23074,32'd23157,32'd23240,32'd23323,32'd23406,32'd23489,32'd23572,32'd23655,32'd23738,32'd23821,32'd23904,32'd23987,32'd24070,32'd24153,32'd24236,32'd24319,32'd24402,32'd24485,32'd24568,32'd24651,32'd24734,32'd24817,32'd24900,32'd24983,32'd25066,32'd25149,32'd25232,32'd25315,32'd25398,32'd25481,32'd25564,32'd25647,32'd25730,32'd25813,32'd25896,32'd25979,32'd26062,32'd26145,32'd26228,32'd26311,32'd26394,32'd26477,32'd26560,32'd26643,32'd26726,32'd26809,32'd26892,32'd26975,32'd27058,32'd27141,32'd27224,32'd27307,32'd27390,32'd27473,32'd27556,32'd27639,32'd27722,32'd27805,32'd27888,32'd27971,32'd28054,32'd28137,32'd28220,32'd28303,32'd28386,32'd28469,32'd28552,32'd28635,32'd28718,32'd28801,32'd28884,32'd28967,32'd29050,32'd29133,32'd29216,32'd29299,32'd29382,32'd29465,32'd29548,32'd29631,32'd29714,32'd29797,32'd29880,32'd29963,32'd30046,32'd30129,32'd30212,32'd30295,32'd30378,32'd30461,32'd30544,32'd30627,32'd30710,32'd30793,32'd30876,32'd30959,32'd31042,32'd31125,32'd31208,32'd31291,32'd31374,32'd31457,32'd31540,32'd31623,32'd31706,32'd31789,32'd31872,32'd31955,32'd32038,32'd32121,32'd32204,32'd32287,32'd32370,32'd32453,32'd32536,32'd32619,32'd32702,32'd32785,32'd32868,32'd32951,32'd33034,32'd33117 };matrix[84]='{32'd0,32'd84,32'd168,32'd252,32'd336,32'd420,32'd504,32'd588,32'd672,32'd756,32'd840,32'd924,32'd1008,32'd1092,32'd1176,32'd1260,32'd1344,32'd1428,32'd1512,32'd1596,32'd1680,32'd1764,32'd1848,32'd1932,32'd2016,32'd2100,32'd2184,32'd2268,32'd2352,32'd2436,32'd2520,32'd2604,32'd2688,32'd2772,32'd2856,32'd2940,32'd3024,32'd3108,32'd3192,32'd3276,32'd3360,32'd3444,32'd3528,32'd3612,32'd3696,32'd3780,32'd3864,32'd3948,32'd4032,32'd4116,32'd4200,32'd4284,32'd4368,32'd4452,32'd4536,32'd4620,32'd4704,32'd4788,32'd4872,32'd4956,32'd5040,32'd5124,32'd5208,32'd5292,32'd5376,32'd5460,32'd5544,32'd5628,32'd5712,32'd5796,32'd5880,32'd5964,32'd6048,32'd6132,32'd6216,32'd6300,32'd6384,32'd6468,32'd6552,32'd6636,32'd6720,32'd6804,32'd6888,32'd6972,32'd7056,32'd7140,32'd7224,32'd7308,32'd7392,32'd7476,32'd7560,32'd7644,32'd7728,32'd7812,32'd7896,32'd7980,32'd8064,32'd8148,32'd8232,32'd8316,32'd8400,32'd8484,32'd8568,32'd8652,32'd8736,32'd8820,32'd8904,32'd8988,32'd9072,32'd9156,32'd9240,32'd9324,32'd9408,32'd9492,32'd9576,32'd9660,32'd9744,32'd9828,32'd9912,32'd9996,32'd10080,32'd10164,32'd10248,32'd10332,32'd10416,32'd10500,32'd10584,32'd10668,32'd10752,32'd10836,32'd10920,32'd11004,32'd11088,32'd11172,32'd11256,32'd11340,32'd11424,32'd11508,32'd11592,32'd11676,32'd11760,32'd11844,32'd11928,32'd12012,32'd12096,32'd12180,32'd12264,32'd12348,32'd12432,32'd12516,32'd12600,32'd12684,32'd12768,32'd12852,32'd12936,32'd13020,32'd13104,32'd13188,32'd13272,32'd13356,32'd13440,32'd13524,32'd13608,32'd13692,32'd13776,32'd13860,32'd13944,32'd14028,32'd14112,32'd14196,32'd14280,32'd14364,32'd14448,32'd14532,32'd14616,32'd14700,32'd14784,32'd14868,32'd14952,32'd15036,32'd15120,32'd15204,32'd15288,32'd15372,32'd15456,32'd15540,32'd15624,32'd15708,32'd15792,32'd15876,32'd15960,32'd16044,32'd16128,32'd16212,32'd16296,32'd16380,32'd16464,32'd16548,32'd16632,32'd16716,32'd16800,32'd16884,32'd16968,32'd17052,32'd17136,32'd17220,32'd17304,32'd17388,32'd17472,32'd17556,32'd17640,32'd17724,32'd17808,32'd17892,32'd17976,32'd18060,32'd18144,32'd18228,32'd18312,32'd18396,32'd18480,32'd18564,32'd18648,32'd18732,32'd18816,32'd18900,32'd18984,32'd19068,32'd19152,32'd19236,32'd19320,32'd19404,32'd19488,32'd19572,32'd19656,32'd19740,32'd19824,32'd19908,32'd19992,32'd20076,32'd20160,32'd20244,32'd20328,32'd20412,32'd20496,32'd20580,32'd20664,32'd20748,32'd20832,32'd20916,32'd21000,32'd21084,32'd21168,32'd21252,32'd21336,32'd21420,32'd21504,32'd21588,32'd21672,32'd21756,32'd21840,32'd21924,32'd22008,32'd22092,32'd22176,32'd22260,32'd22344,32'd22428,32'd22512,32'd22596,32'd22680,32'd22764,32'd22848,32'd22932,32'd23016,32'd23100,32'd23184,32'd23268,32'd23352,32'd23436,32'd23520,32'd23604,32'd23688,32'd23772,32'd23856,32'd23940,32'd24024,32'd24108,32'd24192,32'd24276,32'd24360,32'd24444,32'd24528,32'd24612,32'd24696,32'd24780,32'd24864,32'd24948,32'd25032,32'd25116,32'd25200,32'd25284,32'd25368,32'd25452,32'd25536,32'd25620,32'd25704,32'd25788,32'd25872,32'd25956,32'd26040,32'd26124,32'd26208,32'd26292,32'd26376,32'd26460,32'd26544,32'd26628,32'd26712,32'd26796,32'd26880,32'd26964,32'd27048,32'd27132,32'd27216,32'd27300,32'd27384,32'd27468,32'd27552,32'd27636,32'd27720,32'd27804,32'd27888,32'd27972,32'd28056,32'd28140,32'd28224,32'd28308,32'd28392,32'd28476,32'd28560,32'd28644,32'd28728,32'd28812,32'd28896,32'd28980,32'd29064,32'd29148,32'd29232,32'd29316,32'd29400,32'd29484,32'd29568,32'd29652,32'd29736,32'd29820,32'd29904,32'd29988,32'd30072,32'd30156,32'd30240,32'd30324,32'd30408,32'd30492,32'd30576,32'd30660,32'd30744,32'd30828,32'd30912,32'd30996,32'd31080,32'd31164,32'd31248,32'd31332,32'd31416,32'd31500,32'd31584,32'd31668,32'd31752,32'd31836,32'd31920,32'd32004,32'd32088,32'd32172,32'd32256,32'd32340,32'd32424,32'd32508,32'd32592,32'd32676,32'd32760,32'd32844,32'd32928,32'd33012,32'd33096,32'd33180,32'd33264,32'd33348,32'd33432,32'd33516 };matrix[85]='{32'd0,32'd85,32'd170,32'd255,32'd340,32'd425,32'd510,32'd595,32'd680,32'd765,32'd850,32'd935,32'd1020,32'd1105,32'd1190,32'd1275,32'd1360,32'd1445,32'd1530,32'd1615,32'd1700,32'd1785,32'd1870,32'd1955,32'd2040,32'd2125,32'd2210,32'd2295,32'd2380,32'd2465,32'd2550,32'd2635,32'd2720,32'd2805,32'd2890,32'd2975,32'd3060,32'd3145,32'd3230,32'd3315,32'd3400,32'd3485,32'd3570,32'd3655,32'd3740,32'd3825,32'd3910,32'd3995,32'd4080,32'd4165,32'd4250,32'd4335,32'd4420,32'd4505,32'd4590,32'd4675,32'd4760,32'd4845,32'd4930,32'd5015,32'd5100,32'd5185,32'd5270,32'd5355,32'd5440,32'd5525,32'd5610,32'd5695,32'd5780,32'd5865,32'd5950,32'd6035,32'd6120,32'd6205,32'd6290,32'd6375,32'd6460,32'd6545,32'd6630,32'd6715,32'd6800,32'd6885,32'd6970,32'd7055,32'd7140,32'd7225,32'd7310,32'd7395,32'd7480,32'd7565,32'd7650,32'd7735,32'd7820,32'd7905,32'd7990,32'd8075,32'd8160,32'd8245,32'd8330,32'd8415,32'd8500,32'd8585,32'd8670,32'd8755,32'd8840,32'd8925,32'd9010,32'd9095,32'd9180,32'd9265,32'd9350,32'd9435,32'd9520,32'd9605,32'd9690,32'd9775,32'd9860,32'd9945,32'd10030,32'd10115,32'd10200,32'd10285,32'd10370,32'd10455,32'd10540,32'd10625,32'd10710,32'd10795,32'd10880,32'd10965,32'd11050,32'd11135,32'd11220,32'd11305,32'd11390,32'd11475,32'd11560,32'd11645,32'd11730,32'd11815,32'd11900,32'd11985,32'd12070,32'd12155,32'd12240,32'd12325,32'd12410,32'd12495,32'd12580,32'd12665,32'd12750,32'd12835,32'd12920,32'd13005,32'd13090,32'd13175,32'd13260,32'd13345,32'd13430,32'd13515,32'd13600,32'd13685,32'd13770,32'd13855,32'd13940,32'd14025,32'd14110,32'd14195,32'd14280,32'd14365,32'd14450,32'd14535,32'd14620,32'd14705,32'd14790,32'd14875,32'd14960,32'd15045,32'd15130,32'd15215,32'd15300,32'd15385,32'd15470,32'd15555,32'd15640,32'd15725,32'd15810,32'd15895,32'd15980,32'd16065,32'd16150,32'd16235,32'd16320,32'd16405,32'd16490,32'd16575,32'd16660,32'd16745,32'd16830,32'd16915,32'd17000,32'd17085,32'd17170,32'd17255,32'd17340,32'd17425,32'd17510,32'd17595,32'd17680,32'd17765,32'd17850,32'd17935,32'd18020,32'd18105,32'd18190,32'd18275,32'd18360,32'd18445,32'd18530,32'd18615,32'd18700,32'd18785,32'd18870,32'd18955,32'd19040,32'd19125,32'd19210,32'd19295,32'd19380,32'd19465,32'd19550,32'd19635,32'd19720,32'd19805,32'd19890,32'd19975,32'd20060,32'd20145,32'd20230,32'd20315,32'd20400,32'd20485,32'd20570,32'd20655,32'd20740,32'd20825,32'd20910,32'd20995,32'd21080,32'd21165,32'd21250,32'd21335,32'd21420,32'd21505,32'd21590,32'd21675,32'd21760,32'd21845,32'd21930,32'd22015,32'd22100,32'd22185,32'd22270,32'd22355,32'd22440,32'd22525,32'd22610,32'd22695,32'd22780,32'd22865,32'd22950,32'd23035,32'd23120,32'd23205,32'd23290,32'd23375,32'd23460,32'd23545,32'd23630,32'd23715,32'd23800,32'd23885,32'd23970,32'd24055,32'd24140,32'd24225,32'd24310,32'd24395,32'd24480,32'd24565,32'd24650,32'd24735,32'd24820,32'd24905,32'd24990,32'd25075,32'd25160,32'd25245,32'd25330,32'd25415,32'd25500,32'd25585,32'd25670,32'd25755,32'd25840,32'd25925,32'd26010,32'd26095,32'd26180,32'd26265,32'd26350,32'd26435,32'd26520,32'd26605,32'd26690,32'd26775,32'd26860,32'd26945,32'd27030,32'd27115,32'd27200,32'd27285,32'd27370,32'd27455,32'd27540,32'd27625,32'd27710,32'd27795,32'd27880,32'd27965,32'd28050,32'd28135,32'd28220,32'd28305,32'd28390,32'd28475,32'd28560,32'd28645,32'd28730,32'd28815,32'd28900,32'd28985,32'd29070,32'd29155,32'd29240,32'd29325,32'd29410,32'd29495,32'd29580,32'd29665,32'd29750,32'd29835,32'd29920,32'd30005,32'd30090,32'd30175,32'd30260,32'd30345,32'd30430,32'd30515,32'd30600,32'd30685,32'd30770,32'd30855,32'd30940,32'd31025,32'd31110,32'd31195,32'd31280,32'd31365,32'd31450,32'd31535,32'd31620,32'd31705,32'd31790,32'd31875,32'd31960,32'd32045,32'd32130,32'd32215,32'd32300,32'd32385,32'd32470,32'd32555,32'd32640,32'd32725,32'd32810,32'd32895,32'd32980,32'd33065,32'd33150,32'd33235,32'd33320,32'd33405,32'd33490,32'd33575,32'd33660,32'd33745,32'd33830,32'd33915 };matrix[86]='{32'd0,32'd86,32'd172,32'd258,32'd344,32'd430,32'd516,32'd602,32'd688,32'd774,32'd860,32'd946,32'd1032,32'd1118,32'd1204,32'd1290,32'd1376,32'd1462,32'd1548,32'd1634,32'd1720,32'd1806,32'd1892,32'd1978,32'd2064,32'd2150,32'd2236,32'd2322,32'd2408,32'd2494,32'd2580,32'd2666,32'd2752,32'd2838,32'd2924,32'd3010,32'd3096,32'd3182,32'd3268,32'd3354,32'd3440,32'd3526,32'd3612,32'd3698,32'd3784,32'd3870,32'd3956,32'd4042,32'd4128,32'd4214,32'd4300,32'd4386,32'd4472,32'd4558,32'd4644,32'd4730,32'd4816,32'd4902,32'd4988,32'd5074,32'd5160,32'd5246,32'd5332,32'd5418,32'd5504,32'd5590,32'd5676,32'd5762,32'd5848,32'd5934,32'd6020,32'd6106,32'd6192,32'd6278,32'd6364,32'd6450,32'd6536,32'd6622,32'd6708,32'd6794,32'd6880,32'd6966,32'd7052,32'd7138,32'd7224,32'd7310,32'd7396,32'd7482,32'd7568,32'd7654,32'd7740,32'd7826,32'd7912,32'd7998,32'd8084,32'd8170,32'd8256,32'd8342,32'd8428,32'd8514,32'd8600,32'd8686,32'd8772,32'd8858,32'd8944,32'd9030,32'd9116,32'd9202,32'd9288,32'd9374,32'd9460,32'd9546,32'd9632,32'd9718,32'd9804,32'd9890,32'd9976,32'd10062,32'd10148,32'd10234,32'd10320,32'd10406,32'd10492,32'd10578,32'd10664,32'd10750,32'd10836,32'd10922,32'd11008,32'd11094,32'd11180,32'd11266,32'd11352,32'd11438,32'd11524,32'd11610,32'd11696,32'd11782,32'd11868,32'd11954,32'd12040,32'd12126,32'd12212,32'd12298,32'd12384,32'd12470,32'd12556,32'd12642,32'd12728,32'd12814,32'd12900,32'd12986,32'd13072,32'd13158,32'd13244,32'd13330,32'd13416,32'd13502,32'd13588,32'd13674,32'd13760,32'd13846,32'd13932,32'd14018,32'd14104,32'd14190,32'd14276,32'd14362,32'd14448,32'd14534,32'd14620,32'd14706,32'd14792,32'd14878,32'd14964,32'd15050,32'd15136,32'd15222,32'd15308,32'd15394,32'd15480,32'd15566,32'd15652,32'd15738,32'd15824,32'd15910,32'd15996,32'd16082,32'd16168,32'd16254,32'd16340,32'd16426,32'd16512,32'd16598,32'd16684,32'd16770,32'd16856,32'd16942,32'd17028,32'd17114,32'd17200,32'd17286,32'd17372,32'd17458,32'd17544,32'd17630,32'd17716,32'd17802,32'd17888,32'd17974,32'd18060,32'd18146,32'd18232,32'd18318,32'd18404,32'd18490,32'd18576,32'd18662,32'd18748,32'd18834,32'd18920,32'd19006,32'd19092,32'd19178,32'd19264,32'd19350,32'd19436,32'd19522,32'd19608,32'd19694,32'd19780,32'd19866,32'd19952,32'd20038,32'd20124,32'd20210,32'd20296,32'd20382,32'd20468,32'd20554,32'd20640,32'd20726,32'd20812,32'd20898,32'd20984,32'd21070,32'd21156,32'd21242,32'd21328,32'd21414,32'd21500,32'd21586,32'd21672,32'd21758,32'd21844,32'd21930,32'd22016,32'd22102,32'd22188,32'd22274,32'd22360,32'd22446,32'd22532,32'd22618,32'd22704,32'd22790,32'd22876,32'd22962,32'd23048,32'd23134,32'd23220,32'd23306,32'd23392,32'd23478,32'd23564,32'd23650,32'd23736,32'd23822,32'd23908,32'd23994,32'd24080,32'd24166,32'd24252,32'd24338,32'd24424,32'd24510,32'd24596,32'd24682,32'd24768,32'd24854,32'd24940,32'd25026,32'd25112,32'd25198,32'd25284,32'd25370,32'd25456,32'd25542,32'd25628,32'd25714,32'd25800,32'd25886,32'd25972,32'd26058,32'd26144,32'd26230,32'd26316,32'd26402,32'd26488,32'd26574,32'd26660,32'd26746,32'd26832,32'd26918,32'd27004,32'd27090,32'd27176,32'd27262,32'd27348,32'd27434,32'd27520,32'd27606,32'd27692,32'd27778,32'd27864,32'd27950,32'd28036,32'd28122,32'd28208,32'd28294,32'd28380,32'd28466,32'd28552,32'd28638,32'd28724,32'd28810,32'd28896,32'd28982,32'd29068,32'd29154,32'd29240,32'd29326,32'd29412,32'd29498,32'd29584,32'd29670,32'd29756,32'd29842,32'd29928,32'd30014,32'd30100,32'd30186,32'd30272,32'd30358,32'd30444,32'd30530,32'd30616,32'd30702,32'd30788,32'd30874,32'd30960,32'd31046,32'd31132,32'd31218,32'd31304,32'd31390,32'd31476,32'd31562,32'd31648,32'd31734,32'd31820,32'd31906,32'd31992,32'd32078,32'd32164,32'd32250,32'd32336,32'd32422,32'd32508,32'd32594,32'd32680,32'd32766,32'd32852,32'd32938,32'd33024,32'd33110,32'd33196,32'd33282,32'd33368,32'd33454,32'd33540,32'd33626,32'd33712,32'd33798,32'd33884,32'd33970,32'd34056,32'd34142,32'd34228,32'd34314 };matrix[87]='{32'd0,32'd87,32'd174,32'd261,32'd348,32'd435,32'd522,32'd609,32'd696,32'd783,32'd870,32'd957,32'd1044,32'd1131,32'd1218,32'd1305,32'd1392,32'd1479,32'd1566,32'd1653,32'd1740,32'd1827,32'd1914,32'd2001,32'd2088,32'd2175,32'd2262,32'd2349,32'd2436,32'd2523,32'd2610,32'd2697,32'd2784,32'd2871,32'd2958,32'd3045,32'd3132,32'd3219,32'd3306,32'd3393,32'd3480,32'd3567,32'd3654,32'd3741,32'd3828,32'd3915,32'd4002,32'd4089,32'd4176,32'd4263,32'd4350,32'd4437,32'd4524,32'd4611,32'd4698,32'd4785,32'd4872,32'd4959,32'd5046,32'd5133,32'd5220,32'd5307,32'd5394,32'd5481,32'd5568,32'd5655,32'd5742,32'd5829,32'd5916,32'd6003,32'd6090,32'd6177,32'd6264,32'd6351,32'd6438,32'd6525,32'd6612,32'd6699,32'd6786,32'd6873,32'd6960,32'd7047,32'd7134,32'd7221,32'd7308,32'd7395,32'd7482,32'd7569,32'd7656,32'd7743,32'd7830,32'd7917,32'd8004,32'd8091,32'd8178,32'd8265,32'd8352,32'd8439,32'd8526,32'd8613,32'd8700,32'd8787,32'd8874,32'd8961,32'd9048,32'd9135,32'd9222,32'd9309,32'd9396,32'd9483,32'd9570,32'd9657,32'd9744,32'd9831,32'd9918,32'd10005,32'd10092,32'd10179,32'd10266,32'd10353,32'd10440,32'd10527,32'd10614,32'd10701,32'd10788,32'd10875,32'd10962,32'd11049,32'd11136,32'd11223,32'd11310,32'd11397,32'd11484,32'd11571,32'd11658,32'd11745,32'd11832,32'd11919,32'd12006,32'd12093,32'd12180,32'd12267,32'd12354,32'd12441,32'd12528,32'd12615,32'd12702,32'd12789,32'd12876,32'd12963,32'd13050,32'd13137,32'd13224,32'd13311,32'd13398,32'd13485,32'd13572,32'd13659,32'd13746,32'd13833,32'd13920,32'd14007,32'd14094,32'd14181,32'd14268,32'd14355,32'd14442,32'd14529,32'd14616,32'd14703,32'd14790,32'd14877,32'd14964,32'd15051,32'd15138,32'd15225,32'd15312,32'd15399,32'd15486,32'd15573,32'd15660,32'd15747,32'd15834,32'd15921,32'd16008,32'd16095,32'd16182,32'd16269,32'd16356,32'd16443,32'd16530,32'd16617,32'd16704,32'd16791,32'd16878,32'd16965,32'd17052,32'd17139,32'd17226,32'd17313,32'd17400,32'd17487,32'd17574,32'd17661,32'd17748,32'd17835,32'd17922,32'd18009,32'd18096,32'd18183,32'd18270,32'd18357,32'd18444,32'd18531,32'd18618,32'd18705,32'd18792,32'd18879,32'd18966,32'd19053,32'd19140,32'd19227,32'd19314,32'd19401,32'd19488,32'd19575,32'd19662,32'd19749,32'd19836,32'd19923,32'd20010,32'd20097,32'd20184,32'd20271,32'd20358,32'd20445,32'd20532,32'd20619,32'd20706,32'd20793,32'd20880,32'd20967,32'd21054,32'd21141,32'd21228,32'd21315,32'd21402,32'd21489,32'd21576,32'd21663,32'd21750,32'd21837,32'd21924,32'd22011,32'd22098,32'd22185,32'd22272,32'd22359,32'd22446,32'd22533,32'd22620,32'd22707,32'd22794,32'd22881,32'd22968,32'd23055,32'd23142,32'd23229,32'd23316,32'd23403,32'd23490,32'd23577,32'd23664,32'd23751,32'd23838,32'd23925,32'd24012,32'd24099,32'd24186,32'd24273,32'd24360,32'd24447,32'd24534,32'd24621,32'd24708,32'd24795,32'd24882,32'd24969,32'd25056,32'd25143,32'd25230,32'd25317,32'd25404,32'd25491,32'd25578,32'd25665,32'd25752,32'd25839,32'd25926,32'd26013,32'd26100,32'd26187,32'd26274,32'd26361,32'd26448,32'd26535,32'd26622,32'd26709,32'd26796,32'd26883,32'd26970,32'd27057,32'd27144,32'd27231,32'd27318,32'd27405,32'd27492,32'd27579,32'd27666,32'd27753,32'd27840,32'd27927,32'd28014,32'd28101,32'd28188,32'd28275,32'd28362,32'd28449,32'd28536,32'd28623,32'd28710,32'd28797,32'd28884,32'd28971,32'd29058,32'd29145,32'd29232,32'd29319,32'd29406,32'd29493,32'd29580,32'd29667,32'd29754,32'd29841,32'd29928,32'd30015,32'd30102,32'd30189,32'd30276,32'd30363,32'd30450,32'd30537,32'd30624,32'd30711,32'd30798,32'd30885,32'd30972,32'd31059,32'd31146,32'd31233,32'd31320,32'd31407,32'd31494,32'd31581,32'd31668,32'd31755,32'd31842,32'd31929,32'd32016,32'd32103,32'd32190,32'd32277,32'd32364,32'd32451,32'd32538,32'd32625,32'd32712,32'd32799,32'd32886,32'd32973,32'd33060,32'd33147,32'd33234,32'd33321,32'd33408,32'd33495,32'd33582,32'd33669,32'd33756,32'd33843,32'd33930,32'd34017,32'd34104,32'd34191,32'd34278,32'd34365,32'd34452,32'd34539,32'd34626,32'd34713 };matrix[88]='{32'd0,32'd88,32'd176,32'd264,32'd352,32'd440,32'd528,32'd616,32'd704,32'd792,32'd880,32'd968,32'd1056,32'd1144,32'd1232,32'd1320,32'd1408,32'd1496,32'd1584,32'd1672,32'd1760,32'd1848,32'd1936,32'd2024,32'd2112,32'd2200,32'd2288,32'd2376,32'd2464,32'd2552,32'd2640,32'd2728,32'd2816,32'd2904,32'd2992,32'd3080,32'd3168,32'd3256,32'd3344,32'd3432,32'd3520,32'd3608,32'd3696,32'd3784,32'd3872,32'd3960,32'd4048,32'd4136,32'd4224,32'd4312,32'd4400,32'd4488,32'd4576,32'd4664,32'd4752,32'd4840,32'd4928,32'd5016,32'd5104,32'd5192,32'd5280,32'd5368,32'd5456,32'd5544,32'd5632,32'd5720,32'd5808,32'd5896,32'd5984,32'd6072,32'd6160,32'd6248,32'd6336,32'd6424,32'd6512,32'd6600,32'd6688,32'd6776,32'd6864,32'd6952,32'd7040,32'd7128,32'd7216,32'd7304,32'd7392,32'd7480,32'd7568,32'd7656,32'd7744,32'd7832,32'd7920,32'd8008,32'd8096,32'd8184,32'd8272,32'd8360,32'd8448,32'd8536,32'd8624,32'd8712,32'd8800,32'd8888,32'd8976,32'd9064,32'd9152,32'd9240,32'd9328,32'd9416,32'd9504,32'd9592,32'd9680,32'd9768,32'd9856,32'd9944,32'd10032,32'd10120,32'd10208,32'd10296,32'd10384,32'd10472,32'd10560,32'd10648,32'd10736,32'd10824,32'd10912,32'd11000,32'd11088,32'd11176,32'd11264,32'd11352,32'd11440,32'd11528,32'd11616,32'd11704,32'd11792,32'd11880,32'd11968,32'd12056,32'd12144,32'd12232,32'd12320,32'd12408,32'd12496,32'd12584,32'd12672,32'd12760,32'd12848,32'd12936,32'd13024,32'd13112,32'd13200,32'd13288,32'd13376,32'd13464,32'd13552,32'd13640,32'd13728,32'd13816,32'd13904,32'd13992,32'd14080,32'd14168,32'd14256,32'd14344,32'd14432,32'd14520,32'd14608,32'd14696,32'd14784,32'd14872,32'd14960,32'd15048,32'd15136,32'd15224,32'd15312,32'd15400,32'd15488,32'd15576,32'd15664,32'd15752,32'd15840,32'd15928,32'd16016,32'd16104,32'd16192,32'd16280,32'd16368,32'd16456,32'd16544,32'd16632,32'd16720,32'd16808,32'd16896,32'd16984,32'd17072,32'd17160,32'd17248,32'd17336,32'd17424,32'd17512,32'd17600,32'd17688,32'd17776,32'd17864,32'd17952,32'd18040,32'd18128,32'd18216,32'd18304,32'd18392,32'd18480,32'd18568,32'd18656,32'd18744,32'd18832,32'd18920,32'd19008,32'd19096,32'd19184,32'd19272,32'd19360,32'd19448,32'd19536,32'd19624,32'd19712,32'd19800,32'd19888,32'd19976,32'd20064,32'd20152,32'd20240,32'd20328,32'd20416,32'd20504,32'd20592,32'd20680,32'd20768,32'd20856,32'd20944,32'd21032,32'd21120,32'd21208,32'd21296,32'd21384,32'd21472,32'd21560,32'd21648,32'd21736,32'd21824,32'd21912,32'd22000,32'd22088,32'd22176,32'd22264,32'd22352,32'd22440,32'd22528,32'd22616,32'd22704,32'd22792,32'd22880,32'd22968,32'd23056,32'd23144,32'd23232,32'd23320,32'd23408,32'd23496,32'd23584,32'd23672,32'd23760,32'd23848,32'd23936,32'd24024,32'd24112,32'd24200,32'd24288,32'd24376,32'd24464,32'd24552,32'd24640,32'd24728,32'd24816,32'd24904,32'd24992,32'd25080,32'd25168,32'd25256,32'd25344,32'd25432,32'd25520,32'd25608,32'd25696,32'd25784,32'd25872,32'd25960,32'd26048,32'd26136,32'd26224,32'd26312,32'd26400,32'd26488,32'd26576,32'd26664,32'd26752,32'd26840,32'd26928,32'd27016,32'd27104,32'd27192,32'd27280,32'd27368,32'd27456,32'd27544,32'd27632,32'd27720,32'd27808,32'd27896,32'd27984,32'd28072,32'd28160,32'd28248,32'd28336,32'd28424,32'd28512,32'd28600,32'd28688,32'd28776,32'd28864,32'd28952,32'd29040,32'd29128,32'd29216,32'd29304,32'd29392,32'd29480,32'd29568,32'd29656,32'd29744,32'd29832,32'd29920,32'd30008,32'd30096,32'd30184,32'd30272,32'd30360,32'd30448,32'd30536,32'd30624,32'd30712,32'd30800,32'd30888,32'd30976,32'd31064,32'd31152,32'd31240,32'd31328,32'd31416,32'd31504,32'd31592,32'd31680,32'd31768,32'd31856,32'd31944,32'd32032,32'd32120,32'd32208,32'd32296,32'd32384,32'd32472,32'd32560,32'd32648,32'd32736,32'd32824,32'd32912,32'd33000,32'd33088,32'd33176,32'd33264,32'd33352,32'd33440,32'd33528,32'd33616,32'd33704,32'd33792,32'd33880,32'd33968,32'd34056,32'd34144,32'd34232,32'd34320,32'd34408,32'd34496,32'd34584,32'd34672,32'd34760,32'd34848,32'd34936,32'd35024,32'd35112 };matrix[89]='{32'd0,32'd89,32'd178,32'd267,32'd356,32'd445,32'd534,32'd623,32'd712,32'd801,32'd890,32'd979,32'd1068,32'd1157,32'd1246,32'd1335,32'd1424,32'd1513,32'd1602,32'd1691,32'd1780,32'd1869,32'd1958,32'd2047,32'd2136,32'd2225,32'd2314,32'd2403,32'd2492,32'd2581,32'd2670,32'd2759,32'd2848,32'd2937,32'd3026,32'd3115,32'd3204,32'd3293,32'd3382,32'd3471,32'd3560,32'd3649,32'd3738,32'd3827,32'd3916,32'd4005,32'd4094,32'd4183,32'd4272,32'd4361,32'd4450,32'd4539,32'd4628,32'd4717,32'd4806,32'd4895,32'd4984,32'd5073,32'd5162,32'd5251,32'd5340,32'd5429,32'd5518,32'd5607,32'd5696,32'd5785,32'd5874,32'd5963,32'd6052,32'd6141,32'd6230,32'd6319,32'd6408,32'd6497,32'd6586,32'd6675,32'd6764,32'd6853,32'd6942,32'd7031,32'd7120,32'd7209,32'd7298,32'd7387,32'd7476,32'd7565,32'd7654,32'd7743,32'd7832,32'd7921,32'd8010,32'd8099,32'd8188,32'd8277,32'd8366,32'd8455,32'd8544,32'd8633,32'd8722,32'd8811,32'd8900,32'd8989,32'd9078,32'd9167,32'd9256,32'd9345,32'd9434,32'd9523,32'd9612,32'd9701,32'd9790,32'd9879,32'd9968,32'd10057,32'd10146,32'd10235,32'd10324,32'd10413,32'd10502,32'd10591,32'd10680,32'd10769,32'd10858,32'd10947,32'd11036,32'd11125,32'd11214,32'd11303,32'd11392,32'd11481,32'd11570,32'd11659,32'd11748,32'd11837,32'd11926,32'd12015,32'd12104,32'd12193,32'd12282,32'd12371,32'd12460,32'd12549,32'd12638,32'd12727,32'd12816,32'd12905,32'd12994,32'd13083,32'd13172,32'd13261,32'd13350,32'd13439,32'd13528,32'd13617,32'd13706,32'd13795,32'd13884,32'd13973,32'd14062,32'd14151,32'd14240,32'd14329,32'd14418,32'd14507,32'd14596,32'd14685,32'd14774,32'd14863,32'd14952,32'd15041,32'd15130,32'd15219,32'd15308,32'd15397,32'd15486,32'd15575,32'd15664,32'd15753,32'd15842,32'd15931,32'd16020,32'd16109,32'd16198,32'd16287,32'd16376,32'd16465,32'd16554,32'd16643,32'd16732,32'd16821,32'd16910,32'd16999,32'd17088,32'd17177,32'd17266,32'd17355,32'd17444,32'd17533,32'd17622,32'd17711,32'd17800,32'd17889,32'd17978,32'd18067,32'd18156,32'd18245,32'd18334,32'd18423,32'd18512,32'd18601,32'd18690,32'd18779,32'd18868,32'd18957,32'd19046,32'd19135,32'd19224,32'd19313,32'd19402,32'd19491,32'd19580,32'd19669,32'd19758,32'd19847,32'd19936,32'd20025,32'd20114,32'd20203,32'd20292,32'd20381,32'd20470,32'd20559,32'd20648,32'd20737,32'd20826,32'd20915,32'd21004,32'd21093,32'd21182,32'd21271,32'd21360,32'd21449,32'd21538,32'd21627,32'd21716,32'd21805,32'd21894,32'd21983,32'd22072,32'd22161,32'd22250,32'd22339,32'd22428,32'd22517,32'd22606,32'd22695,32'd22784,32'd22873,32'd22962,32'd23051,32'd23140,32'd23229,32'd23318,32'd23407,32'd23496,32'd23585,32'd23674,32'd23763,32'd23852,32'd23941,32'd24030,32'd24119,32'd24208,32'd24297,32'd24386,32'd24475,32'd24564,32'd24653,32'd24742,32'd24831,32'd24920,32'd25009,32'd25098,32'd25187,32'd25276,32'd25365,32'd25454,32'd25543,32'd25632,32'd25721,32'd25810,32'd25899,32'd25988,32'd26077,32'd26166,32'd26255,32'd26344,32'd26433,32'd26522,32'd26611,32'd26700,32'd26789,32'd26878,32'd26967,32'd27056,32'd27145,32'd27234,32'd27323,32'd27412,32'd27501,32'd27590,32'd27679,32'd27768,32'd27857,32'd27946,32'd28035,32'd28124,32'd28213,32'd28302,32'd28391,32'd28480,32'd28569,32'd28658,32'd28747,32'd28836,32'd28925,32'd29014,32'd29103,32'd29192,32'd29281,32'd29370,32'd29459,32'd29548,32'd29637,32'd29726,32'd29815,32'd29904,32'd29993,32'd30082,32'd30171,32'd30260,32'd30349,32'd30438,32'd30527,32'd30616,32'd30705,32'd30794,32'd30883,32'd30972,32'd31061,32'd31150,32'd31239,32'd31328,32'd31417,32'd31506,32'd31595,32'd31684,32'd31773,32'd31862,32'd31951,32'd32040,32'd32129,32'd32218,32'd32307,32'd32396,32'd32485,32'd32574,32'd32663,32'd32752,32'd32841,32'd32930,32'd33019,32'd33108,32'd33197,32'd33286,32'd33375,32'd33464,32'd33553,32'd33642,32'd33731,32'd33820,32'd33909,32'd33998,32'd34087,32'd34176,32'd34265,32'd34354,32'd34443,32'd34532,32'd34621,32'd34710,32'd34799,32'd34888,32'd34977,32'd35066,32'd35155,32'd35244,32'd35333,32'd35422,32'd35511 };matrix[90]='{32'd0,32'd90,32'd180,32'd270,32'd360,32'd450,32'd540,32'd630,32'd720,32'd810,32'd900,32'd990,32'd1080,32'd1170,32'd1260,32'd1350,32'd1440,32'd1530,32'd1620,32'd1710,32'd1800,32'd1890,32'd1980,32'd2070,32'd2160,32'd2250,32'd2340,32'd2430,32'd2520,32'd2610,32'd2700,32'd2790,32'd2880,32'd2970,32'd3060,32'd3150,32'd3240,32'd3330,32'd3420,32'd3510,32'd3600,32'd3690,32'd3780,32'd3870,32'd3960,32'd4050,32'd4140,32'd4230,32'd4320,32'd4410,32'd4500,32'd4590,32'd4680,32'd4770,32'd4860,32'd4950,32'd5040,32'd5130,32'd5220,32'd5310,32'd5400,32'd5490,32'd5580,32'd5670,32'd5760,32'd5850,32'd5940,32'd6030,32'd6120,32'd6210,32'd6300,32'd6390,32'd6480,32'd6570,32'd6660,32'd6750,32'd6840,32'd6930,32'd7020,32'd7110,32'd7200,32'd7290,32'd7380,32'd7470,32'd7560,32'd7650,32'd7740,32'd7830,32'd7920,32'd8010,32'd8100,32'd8190,32'd8280,32'd8370,32'd8460,32'd8550,32'd8640,32'd8730,32'd8820,32'd8910,32'd9000,32'd9090,32'd9180,32'd9270,32'd9360,32'd9450,32'd9540,32'd9630,32'd9720,32'd9810,32'd9900,32'd9990,32'd10080,32'd10170,32'd10260,32'd10350,32'd10440,32'd10530,32'd10620,32'd10710,32'd10800,32'd10890,32'd10980,32'd11070,32'd11160,32'd11250,32'd11340,32'd11430,32'd11520,32'd11610,32'd11700,32'd11790,32'd11880,32'd11970,32'd12060,32'd12150,32'd12240,32'd12330,32'd12420,32'd12510,32'd12600,32'd12690,32'd12780,32'd12870,32'd12960,32'd13050,32'd13140,32'd13230,32'd13320,32'd13410,32'd13500,32'd13590,32'd13680,32'd13770,32'd13860,32'd13950,32'd14040,32'd14130,32'd14220,32'd14310,32'd14400,32'd14490,32'd14580,32'd14670,32'd14760,32'd14850,32'd14940,32'd15030,32'd15120,32'd15210,32'd15300,32'd15390,32'd15480,32'd15570,32'd15660,32'd15750,32'd15840,32'd15930,32'd16020,32'd16110,32'd16200,32'd16290,32'd16380,32'd16470,32'd16560,32'd16650,32'd16740,32'd16830,32'd16920,32'd17010,32'd17100,32'd17190,32'd17280,32'd17370,32'd17460,32'd17550,32'd17640,32'd17730,32'd17820,32'd17910,32'd18000,32'd18090,32'd18180,32'd18270,32'd18360,32'd18450,32'd18540,32'd18630,32'd18720,32'd18810,32'd18900,32'd18990,32'd19080,32'd19170,32'd19260,32'd19350,32'd19440,32'd19530,32'd19620,32'd19710,32'd19800,32'd19890,32'd19980,32'd20070,32'd20160,32'd20250,32'd20340,32'd20430,32'd20520,32'd20610,32'd20700,32'd20790,32'd20880,32'd20970,32'd21060,32'd21150,32'd21240,32'd21330,32'd21420,32'd21510,32'd21600,32'd21690,32'd21780,32'd21870,32'd21960,32'd22050,32'd22140,32'd22230,32'd22320,32'd22410,32'd22500,32'd22590,32'd22680,32'd22770,32'd22860,32'd22950,32'd23040,32'd23130,32'd23220,32'd23310,32'd23400,32'd23490,32'd23580,32'd23670,32'd23760,32'd23850,32'd23940,32'd24030,32'd24120,32'd24210,32'd24300,32'd24390,32'd24480,32'd24570,32'd24660,32'd24750,32'd24840,32'd24930,32'd25020,32'd25110,32'd25200,32'd25290,32'd25380,32'd25470,32'd25560,32'd25650,32'd25740,32'd25830,32'd25920,32'd26010,32'd26100,32'd26190,32'd26280,32'd26370,32'd26460,32'd26550,32'd26640,32'd26730,32'd26820,32'd26910,32'd27000,32'd27090,32'd27180,32'd27270,32'd27360,32'd27450,32'd27540,32'd27630,32'd27720,32'd27810,32'd27900,32'd27990,32'd28080,32'd28170,32'd28260,32'd28350,32'd28440,32'd28530,32'd28620,32'd28710,32'd28800,32'd28890,32'd28980,32'd29070,32'd29160,32'd29250,32'd29340,32'd29430,32'd29520,32'd29610,32'd29700,32'd29790,32'd29880,32'd29970,32'd30060,32'd30150,32'd30240,32'd30330,32'd30420,32'd30510,32'd30600,32'd30690,32'd30780,32'd30870,32'd30960,32'd31050,32'd31140,32'd31230,32'd31320,32'd31410,32'd31500,32'd31590,32'd31680,32'd31770,32'd31860,32'd31950,32'd32040,32'd32130,32'd32220,32'd32310,32'd32400,32'd32490,32'd32580,32'd32670,32'd32760,32'd32850,32'd32940,32'd33030,32'd33120,32'd33210,32'd33300,32'd33390,32'd33480,32'd33570,32'd33660,32'd33750,32'd33840,32'd33930,32'd34020,32'd34110,32'd34200,32'd34290,32'd34380,32'd34470,32'd34560,32'd34650,32'd34740,32'd34830,32'd34920,32'd35010,32'd35100,32'd35190,32'd35280,32'd35370,32'd35460,32'd35550,32'd35640,32'd35730,32'd35820,32'd35910 };matrix[91]='{32'd0,32'd91,32'd182,32'd273,32'd364,32'd455,32'd546,32'd637,32'd728,32'd819,32'd910,32'd1001,32'd1092,32'd1183,32'd1274,32'd1365,32'd1456,32'd1547,32'd1638,32'd1729,32'd1820,32'd1911,32'd2002,32'd2093,32'd2184,32'd2275,32'd2366,32'd2457,32'd2548,32'd2639,32'd2730,32'd2821,32'd2912,32'd3003,32'd3094,32'd3185,32'd3276,32'd3367,32'd3458,32'd3549,32'd3640,32'd3731,32'd3822,32'd3913,32'd4004,32'd4095,32'd4186,32'd4277,32'd4368,32'd4459,32'd4550,32'd4641,32'd4732,32'd4823,32'd4914,32'd5005,32'd5096,32'd5187,32'd5278,32'd5369,32'd5460,32'd5551,32'd5642,32'd5733,32'd5824,32'd5915,32'd6006,32'd6097,32'd6188,32'd6279,32'd6370,32'd6461,32'd6552,32'd6643,32'd6734,32'd6825,32'd6916,32'd7007,32'd7098,32'd7189,32'd7280,32'd7371,32'd7462,32'd7553,32'd7644,32'd7735,32'd7826,32'd7917,32'd8008,32'd8099,32'd8190,32'd8281,32'd8372,32'd8463,32'd8554,32'd8645,32'd8736,32'd8827,32'd8918,32'd9009,32'd9100,32'd9191,32'd9282,32'd9373,32'd9464,32'd9555,32'd9646,32'd9737,32'd9828,32'd9919,32'd10010,32'd10101,32'd10192,32'd10283,32'd10374,32'd10465,32'd10556,32'd10647,32'd10738,32'd10829,32'd10920,32'd11011,32'd11102,32'd11193,32'd11284,32'd11375,32'd11466,32'd11557,32'd11648,32'd11739,32'd11830,32'd11921,32'd12012,32'd12103,32'd12194,32'd12285,32'd12376,32'd12467,32'd12558,32'd12649,32'd12740,32'd12831,32'd12922,32'd13013,32'd13104,32'd13195,32'd13286,32'd13377,32'd13468,32'd13559,32'd13650,32'd13741,32'd13832,32'd13923,32'd14014,32'd14105,32'd14196,32'd14287,32'd14378,32'd14469,32'd14560,32'd14651,32'd14742,32'd14833,32'd14924,32'd15015,32'd15106,32'd15197,32'd15288,32'd15379,32'd15470,32'd15561,32'd15652,32'd15743,32'd15834,32'd15925,32'd16016,32'd16107,32'd16198,32'd16289,32'd16380,32'd16471,32'd16562,32'd16653,32'd16744,32'd16835,32'd16926,32'd17017,32'd17108,32'd17199,32'd17290,32'd17381,32'd17472,32'd17563,32'd17654,32'd17745,32'd17836,32'd17927,32'd18018,32'd18109,32'd18200,32'd18291,32'd18382,32'd18473,32'd18564,32'd18655,32'd18746,32'd18837,32'd18928,32'd19019,32'd19110,32'd19201,32'd19292,32'd19383,32'd19474,32'd19565,32'd19656,32'd19747,32'd19838,32'd19929,32'd20020,32'd20111,32'd20202,32'd20293,32'd20384,32'd20475,32'd20566,32'd20657,32'd20748,32'd20839,32'd20930,32'd21021,32'd21112,32'd21203,32'd21294,32'd21385,32'd21476,32'd21567,32'd21658,32'd21749,32'd21840,32'd21931,32'd22022,32'd22113,32'd22204,32'd22295,32'd22386,32'd22477,32'd22568,32'd22659,32'd22750,32'd22841,32'd22932,32'd23023,32'd23114,32'd23205,32'd23296,32'd23387,32'd23478,32'd23569,32'd23660,32'd23751,32'd23842,32'd23933,32'd24024,32'd24115,32'd24206,32'd24297,32'd24388,32'd24479,32'd24570,32'd24661,32'd24752,32'd24843,32'd24934,32'd25025,32'd25116,32'd25207,32'd25298,32'd25389,32'd25480,32'd25571,32'd25662,32'd25753,32'd25844,32'd25935,32'd26026,32'd26117,32'd26208,32'd26299,32'd26390,32'd26481,32'd26572,32'd26663,32'd26754,32'd26845,32'd26936,32'd27027,32'd27118,32'd27209,32'd27300,32'd27391,32'd27482,32'd27573,32'd27664,32'd27755,32'd27846,32'd27937,32'd28028,32'd28119,32'd28210,32'd28301,32'd28392,32'd28483,32'd28574,32'd28665,32'd28756,32'd28847,32'd28938,32'd29029,32'd29120,32'd29211,32'd29302,32'd29393,32'd29484,32'd29575,32'd29666,32'd29757,32'd29848,32'd29939,32'd30030,32'd30121,32'd30212,32'd30303,32'd30394,32'd30485,32'd30576,32'd30667,32'd30758,32'd30849,32'd30940,32'd31031,32'd31122,32'd31213,32'd31304,32'd31395,32'd31486,32'd31577,32'd31668,32'd31759,32'd31850,32'd31941,32'd32032,32'd32123,32'd32214,32'd32305,32'd32396,32'd32487,32'd32578,32'd32669,32'd32760,32'd32851,32'd32942,32'd33033,32'd33124,32'd33215,32'd33306,32'd33397,32'd33488,32'd33579,32'd33670,32'd33761,32'd33852,32'd33943,32'd34034,32'd34125,32'd34216,32'd34307,32'd34398,32'd34489,32'd34580,32'd34671,32'd34762,32'd34853,32'd34944,32'd35035,32'd35126,32'd35217,32'd35308,32'd35399,32'd35490,32'd35581,32'd35672,32'd35763,32'd35854,32'd35945,32'd36036,32'd36127,32'd36218,32'd36309 };matrix[92]='{32'd0,32'd92,32'd184,32'd276,32'd368,32'd460,32'd552,32'd644,32'd736,32'd828,32'd920,32'd1012,32'd1104,32'd1196,32'd1288,32'd1380,32'd1472,32'd1564,32'd1656,32'd1748,32'd1840,32'd1932,32'd2024,32'd2116,32'd2208,32'd2300,32'd2392,32'd2484,32'd2576,32'd2668,32'd2760,32'd2852,32'd2944,32'd3036,32'd3128,32'd3220,32'd3312,32'd3404,32'd3496,32'd3588,32'd3680,32'd3772,32'd3864,32'd3956,32'd4048,32'd4140,32'd4232,32'd4324,32'd4416,32'd4508,32'd4600,32'd4692,32'd4784,32'd4876,32'd4968,32'd5060,32'd5152,32'd5244,32'd5336,32'd5428,32'd5520,32'd5612,32'd5704,32'd5796,32'd5888,32'd5980,32'd6072,32'd6164,32'd6256,32'd6348,32'd6440,32'd6532,32'd6624,32'd6716,32'd6808,32'd6900,32'd6992,32'd7084,32'd7176,32'd7268,32'd7360,32'd7452,32'd7544,32'd7636,32'd7728,32'd7820,32'd7912,32'd8004,32'd8096,32'd8188,32'd8280,32'd8372,32'd8464,32'd8556,32'd8648,32'd8740,32'd8832,32'd8924,32'd9016,32'd9108,32'd9200,32'd9292,32'd9384,32'd9476,32'd9568,32'd9660,32'd9752,32'd9844,32'd9936,32'd10028,32'd10120,32'd10212,32'd10304,32'd10396,32'd10488,32'd10580,32'd10672,32'd10764,32'd10856,32'd10948,32'd11040,32'd11132,32'd11224,32'd11316,32'd11408,32'd11500,32'd11592,32'd11684,32'd11776,32'd11868,32'd11960,32'd12052,32'd12144,32'd12236,32'd12328,32'd12420,32'd12512,32'd12604,32'd12696,32'd12788,32'd12880,32'd12972,32'd13064,32'd13156,32'd13248,32'd13340,32'd13432,32'd13524,32'd13616,32'd13708,32'd13800,32'd13892,32'd13984,32'd14076,32'd14168,32'd14260,32'd14352,32'd14444,32'd14536,32'd14628,32'd14720,32'd14812,32'd14904,32'd14996,32'd15088,32'd15180,32'd15272,32'd15364,32'd15456,32'd15548,32'd15640,32'd15732,32'd15824,32'd15916,32'd16008,32'd16100,32'd16192,32'd16284,32'd16376,32'd16468,32'd16560,32'd16652,32'd16744,32'd16836,32'd16928,32'd17020,32'd17112,32'd17204,32'd17296,32'd17388,32'd17480,32'd17572,32'd17664,32'd17756,32'd17848,32'd17940,32'd18032,32'd18124,32'd18216,32'd18308,32'd18400,32'd18492,32'd18584,32'd18676,32'd18768,32'd18860,32'd18952,32'd19044,32'd19136,32'd19228,32'd19320,32'd19412,32'd19504,32'd19596,32'd19688,32'd19780,32'd19872,32'd19964,32'd20056,32'd20148,32'd20240,32'd20332,32'd20424,32'd20516,32'd20608,32'd20700,32'd20792,32'd20884,32'd20976,32'd21068,32'd21160,32'd21252,32'd21344,32'd21436,32'd21528,32'd21620,32'd21712,32'd21804,32'd21896,32'd21988,32'd22080,32'd22172,32'd22264,32'd22356,32'd22448,32'd22540,32'd22632,32'd22724,32'd22816,32'd22908,32'd23000,32'd23092,32'd23184,32'd23276,32'd23368,32'd23460,32'd23552,32'd23644,32'd23736,32'd23828,32'd23920,32'd24012,32'd24104,32'd24196,32'd24288,32'd24380,32'd24472,32'd24564,32'd24656,32'd24748,32'd24840,32'd24932,32'd25024,32'd25116,32'd25208,32'd25300,32'd25392,32'd25484,32'd25576,32'd25668,32'd25760,32'd25852,32'd25944,32'd26036,32'd26128,32'd26220,32'd26312,32'd26404,32'd26496,32'd26588,32'd26680,32'd26772,32'd26864,32'd26956,32'd27048,32'd27140,32'd27232,32'd27324,32'd27416,32'd27508,32'd27600,32'd27692,32'd27784,32'd27876,32'd27968,32'd28060,32'd28152,32'd28244,32'd28336,32'd28428,32'd28520,32'd28612,32'd28704,32'd28796,32'd28888,32'd28980,32'd29072,32'd29164,32'd29256,32'd29348,32'd29440,32'd29532,32'd29624,32'd29716,32'd29808,32'd29900,32'd29992,32'd30084,32'd30176,32'd30268,32'd30360,32'd30452,32'd30544,32'd30636,32'd30728,32'd30820,32'd30912,32'd31004,32'd31096,32'd31188,32'd31280,32'd31372,32'd31464,32'd31556,32'd31648,32'd31740,32'd31832,32'd31924,32'd32016,32'd32108,32'd32200,32'd32292,32'd32384,32'd32476,32'd32568,32'd32660,32'd32752,32'd32844,32'd32936,32'd33028,32'd33120,32'd33212,32'd33304,32'd33396,32'd33488,32'd33580,32'd33672,32'd33764,32'd33856,32'd33948,32'd34040,32'd34132,32'd34224,32'd34316,32'd34408,32'd34500,32'd34592,32'd34684,32'd34776,32'd34868,32'd34960,32'd35052,32'd35144,32'd35236,32'd35328,32'd35420,32'd35512,32'd35604,32'd35696,32'd35788,32'd35880,32'd35972,32'd36064,32'd36156,32'd36248,32'd36340,32'd36432,32'd36524,32'd36616,32'd36708 };matrix[93]='{32'd0,32'd93,32'd186,32'd279,32'd372,32'd465,32'd558,32'd651,32'd744,32'd837,32'd930,32'd1023,32'd1116,32'd1209,32'd1302,32'd1395,32'd1488,32'd1581,32'd1674,32'd1767,32'd1860,32'd1953,32'd2046,32'd2139,32'd2232,32'd2325,32'd2418,32'd2511,32'd2604,32'd2697,32'd2790,32'd2883,32'd2976,32'd3069,32'd3162,32'd3255,32'd3348,32'd3441,32'd3534,32'd3627,32'd3720,32'd3813,32'd3906,32'd3999,32'd4092,32'd4185,32'd4278,32'd4371,32'd4464,32'd4557,32'd4650,32'd4743,32'd4836,32'd4929,32'd5022,32'd5115,32'd5208,32'd5301,32'd5394,32'd5487,32'd5580,32'd5673,32'd5766,32'd5859,32'd5952,32'd6045,32'd6138,32'd6231,32'd6324,32'd6417,32'd6510,32'd6603,32'd6696,32'd6789,32'd6882,32'd6975,32'd7068,32'd7161,32'd7254,32'd7347,32'd7440,32'd7533,32'd7626,32'd7719,32'd7812,32'd7905,32'd7998,32'd8091,32'd8184,32'd8277,32'd8370,32'd8463,32'd8556,32'd8649,32'd8742,32'd8835,32'd8928,32'd9021,32'd9114,32'd9207,32'd9300,32'd9393,32'd9486,32'd9579,32'd9672,32'd9765,32'd9858,32'd9951,32'd10044,32'd10137,32'd10230,32'd10323,32'd10416,32'd10509,32'd10602,32'd10695,32'd10788,32'd10881,32'd10974,32'd11067,32'd11160,32'd11253,32'd11346,32'd11439,32'd11532,32'd11625,32'd11718,32'd11811,32'd11904,32'd11997,32'd12090,32'd12183,32'd12276,32'd12369,32'd12462,32'd12555,32'd12648,32'd12741,32'd12834,32'd12927,32'd13020,32'd13113,32'd13206,32'd13299,32'd13392,32'd13485,32'd13578,32'd13671,32'd13764,32'd13857,32'd13950,32'd14043,32'd14136,32'd14229,32'd14322,32'd14415,32'd14508,32'd14601,32'd14694,32'd14787,32'd14880,32'd14973,32'd15066,32'd15159,32'd15252,32'd15345,32'd15438,32'd15531,32'd15624,32'd15717,32'd15810,32'd15903,32'd15996,32'd16089,32'd16182,32'd16275,32'd16368,32'd16461,32'd16554,32'd16647,32'd16740,32'd16833,32'd16926,32'd17019,32'd17112,32'd17205,32'd17298,32'd17391,32'd17484,32'd17577,32'd17670,32'd17763,32'd17856,32'd17949,32'd18042,32'd18135,32'd18228,32'd18321,32'd18414,32'd18507,32'd18600,32'd18693,32'd18786,32'd18879,32'd18972,32'd19065,32'd19158,32'd19251,32'd19344,32'd19437,32'd19530,32'd19623,32'd19716,32'd19809,32'd19902,32'd19995,32'd20088,32'd20181,32'd20274,32'd20367,32'd20460,32'd20553,32'd20646,32'd20739,32'd20832,32'd20925,32'd21018,32'd21111,32'd21204,32'd21297,32'd21390,32'd21483,32'd21576,32'd21669,32'd21762,32'd21855,32'd21948,32'd22041,32'd22134,32'd22227,32'd22320,32'd22413,32'd22506,32'd22599,32'd22692,32'd22785,32'd22878,32'd22971,32'd23064,32'd23157,32'd23250,32'd23343,32'd23436,32'd23529,32'd23622,32'd23715,32'd23808,32'd23901,32'd23994,32'd24087,32'd24180,32'd24273,32'd24366,32'd24459,32'd24552,32'd24645,32'd24738,32'd24831,32'd24924,32'd25017,32'd25110,32'd25203,32'd25296,32'd25389,32'd25482,32'd25575,32'd25668,32'd25761,32'd25854,32'd25947,32'd26040,32'd26133,32'd26226,32'd26319,32'd26412,32'd26505,32'd26598,32'd26691,32'd26784,32'd26877,32'd26970,32'd27063,32'd27156,32'd27249,32'd27342,32'd27435,32'd27528,32'd27621,32'd27714,32'd27807,32'd27900,32'd27993,32'd28086,32'd28179,32'd28272,32'd28365,32'd28458,32'd28551,32'd28644,32'd28737,32'd28830,32'd28923,32'd29016,32'd29109,32'd29202,32'd29295,32'd29388,32'd29481,32'd29574,32'd29667,32'd29760,32'd29853,32'd29946,32'd30039,32'd30132,32'd30225,32'd30318,32'd30411,32'd30504,32'd30597,32'd30690,32'd30783,32'd30876,32'd30969,32'd31062,32'd31155,32'd31248,32'd31341,32'd31434,32'd31527,32'd31620,32'd31713,32'd31806,32'd31899,32'd31992,32'd32085,32'd32178,32'd32271,32'd32364,32'd32457,32'd32550,32'd32643,32'd32736,32'd32829,32'd32922,32'd33015,32'd33108,32'd33201,32'd33294,32'd33387,32'd33480,32'd33573,32'd33666,32'd33759,32'd33852,32'd33945,32'd34038,32'd34131,32'd34224,32'd34317,32'd34410,32'd34503,32'd34596,32'd34689,32'd34782,32'd34875,32'd34968,32'd35061,32'd35154,32'd35247,32'd35340,32'd35433,32'd35526,32'd35619,32'd35712,32'd35805,32'd35898,32'd35991,32'd36084,32'd36177,32'd36270,32'd36363,32'd36456,32'd36549,32'd36642,32'd36735,32'd36828,32'd36921,32'd37014,32'd37107 };matrix[94]='{32'd0,32'd94,32'd188,32'd282,32'd376,32'd470,32'd564,32'd658,32'd752,32'd846,32'd940,32'd1034,32'd1128,32'd1222,32'd1316,32'd1410,32'd1504,32'd1598,32'd1692,32'd1786,32'd1880,32'd1974,32'd2068,32'd2162,32'd2256,32'd2350,32'd2444,32'd2538,32'd2632,32'd2726,32'd2820,32'd2914,32'd3008,32'd3102,32'd3196,32'd3290,32'd3384,32'd3478,32'd3572,32'd3666,32'd3760,32'd3854,32'd3948,32'd4042,32'd4136,32'd4230,32'd4324,32'd4418,32'd4512,32'd4606,32'd4700,32'd4794,32'd4888,32'd4982,32'd5076,32'd5170,32'd5264,32'd5358,32'd5452,32'd5546,32'd5640,32'd5734,32'd5828,32'd5922,32'd6016,32'd6110,32'd6204,32'd6298,32'd6392,32'd6486,32'd6580,32'd6674,32'd6768,32'd6862,32'd6956,32'd7050,32'd7144,32'd7238,32'd7332,32'd7426,32'd7520,32'd7614,32'd7708,32'd7802,32'd7896,32'd7990,32'd8084,32'd8178,32'd8272,32'd8366,32'd8460,32'd8554,32'd8648,32'd8742,32'd8836,32'd8930,32'd9024,32'd9118,32'd9212,32'd9306,32'd9400,32'd9494,32'd9588,32'd9682,32'd9776,32'd9870,32'd9964,32'd10058,32'd10152,32'd10246,32'd10340,32'd10434,32'd10528,32'd10622,32'd10716,32'd10810,32'd10904,32'd10998,32'd11092,32'd11186,32'd11280,32'd11374,32'd11468,32'd11562,32'd11656,32'd11750,32'd11844,32'd11938,32'd12032,32'd12126,32'd12220,32'd12314,32'd12408,32'd12502,32'd12596,32'd12690,32'd12784,32'd12878,32'd12972,32'd13066,32'd13160,32'd13254,32'd13348,32'd13442,32'd13536,32'd13630,32'd13724,32'd13818,32'd13912,32'd14006,32'd14100,32'd14194,32'd14288,32'd14382,32'd14476,32'd14570,32'd14664,32'd14758,32'd14852,32'd14946,32'd15040,32'd15134,32'd15228,32'd15322,32'd15416,32'd15510,32'd15604,32'd15698,32'd15792,32'd15886,32'd15980,32'd16074,32'd16168,32'd16262,32'd16356,32'd16450,32'd16544,32'd16638,32'd16732,32'd16826,32'd16920,32'd17014,32'd17108,32'd17202,32'd17296,32'd17390,32'd17484,32'd17578,32'd17672,32'd17766,32'd17860,32'd17954,32'd18048,32'd18142,32'd18236,32'd18330,32'd18424,32'd18518,32'd18612,32'd18706,32'd18800,32'd18894,32'd18988,32'd19082,32'd19176,32'd19270,32'd19364,32'd19458,32'd19552,32'd19646,32'd19740,32'd19834,32'd19928,32'd20022,32'd20116,32'd20210,32'd20304,32'd20398,32'd20492,32'd20586,32'd20680,32'd20774,32'd20868,32'd20962,32'd21056,32'd21150,32'd21244,32'd21338,32'd21432,32'd21526,32'd21620,32'd21714,32'd21808,32'd21902,32'd21996,32'd22090,32'd22184,32'd22278,32'd22372,32'd22466,32'd22560,32'd22654,32'd22748,32'd22842,32'd22936,32'd23030,32'd23124,32'd23218,32'd23312,32'd23406,32'd23500,32'd23594,32'd23688,32'd23782,32'd23876,32'd23970,32'd24064,32'd24158,32'd24252,32'd24346,32'd24440,32'd24534,32'd24628,32'd24722,32'd24816,32'd24910,32'd25004,32'd25098,32'd25192,32'd25286,32'd25380,32'd25474,32'd25568,32'd25662,32'd25756,32'd25850,32'd25944,32'd26038,32'd26132,32'd26226,32'd26320,32'd26414,32'd26508,32'd26602,32'd26696,32'd26790,32'd26884,32'd26978,32'd27072,32'd27166,32'd27260,32'd27354,32'd27448,32'd27542,32'd27636,32'd27730,32'd27824,32'd27918,32'd28012,32'd28106,32'd28200,32'd28294,32'd28388,32'd28482,32'd28576,32'd28670,32'd28764,32'd28858,32'd28952,32'd29046,32'd29140,32'd29234,32'd29328,32'd29422,32'd29516,32'd29610,32'd29704,32'd29798,32'd29892,32'd29986,32'd30080,32'd30174,32'd30268,32'd30362,32'd30456,32'd30550,32'd30644,32'd30738,32'd30832,32'd30926,32'd31020,32'd31114,32'd31208,32'd31302,32'd31396,32'd31490,32'd31584,32'd31678,32'd31772,32'd31866,32'd31960,32'd32054,32'd32148,32'd32242,32'd32336,32'd32430,32'd32524,32'd32618,32'd32712,32'd32806,32'd32900,32'd32994,32'd33088,32'd33182,32'd33276,32'd33370,32'd33464,32'd33558,32'd33652,32'd33746,32'd33840,32'd33934,32'd34028,32'd34122,32'd34216,32'd34310,32'd34404,32'd34498,32'd34592,32'd34686,32'd34780,32'd34874,32'd34968,32'd35062,32'd35156,32'd35250,32'd35344,32'd35438,32'd35532,32'd35626,32'd35720,32'd35814,32'd35908,32'd36002,32'd36096,32'd36190,32'd36284,32'd36378,32'd36472,32'd36566,32'd36660,32'd36754,32'd36848,32'd36942,32'd37036,32'd37130,32'd37224,32'd37318,32'd37412,32'd37506 };matrix[95]='{32'd0,32'd95,32'd190,32'd285,32'd380,32'd475,32'd570,32'd665,32'd760,32'd855,32'd950,32'd1045,32'd1140,32'd1235,32'd1330,32'd1425,32'd1520,32'd1615,32'd1710,32'd1805,32'd1900,32'd1995,32'd2090,32'd2185,32'd2280,32'd2375,32'd2470,32'd2565,32'd2660,32'd2755,32'd2850,32'd2945,32'd3040,32'd3135,32'd3230,32'd3325,32'd3420,32'd3515,32'd3610,32'd3705,32'd3800,32'd3895,32'd3990,32'd4085,32'd4180,32'd4275,32'd4370,32'd4465,32'd4560,32'd4655,32'd4750,32'd4845,32'd4940,32'd5035,32'd5130,32'd5225,32'd5320,32'd5415,32'd5510,32'd5605,32'd5700,32'd5795,32'd5890,32'd5985,32'd6080,32'd6175,32'd6270,32'd6365,32'd6460,32'd6555,32'd6650,32'd6745,32'd6840,32'd6935,32'd7030,32'd7125,32'd7220,32'd7315,32'd7410,32'd7505,32'd7600,32'd7695,32'd7790,32'd7885,32'd7980,32'd8075,32'd8170,32'd8265,32'd8360,32'd8455,32'd8550,32'd8645,32'd8740,32'd8835,32'd8930,32'd9025,32'd9120,32'd9215,32'd9310,32'd9405,32'd9500,32'd9595,32'd9690,32'd9785,32'd9880,32'd9975,32'd10070,32'd10165,32'd10260,32'd10355,32'd10450,32'd10545,32'd10640,32'd10735,32'd10830,32'd10925,32'd11020,32'd11115,32'd11210,32'd11305,32'd11400,32'd11495,32'd11590,32'd11685,32'd11780,32'd11875,32'd11970,32'd12065,32'd12160,32'd12255,32'd12350,32'd12445,32'd12540,32'd12635,32'd12730,32'd12825,32'd12920,32'd13015,32'd13110,32'd13205,32'd13300,32'd13395,32'd13490,32'd13585,32'd13680,32'd13775,32'd13870,32'd13965,32'd14060,32'd14155,32'd14250,32'd14345,32'd14440,32'd14535,32'd14630,32'd14725,32'd14820,32'd14915,32'd15010,32'd15105,32'd15200,32'd15295,32'd15390,32'd15485,32'd15580,32'd15675,32'd15770,32'd15865,32'd15960,32'd16055,32'd16150,32'd16245,32'd16340,32'd16435,32'd16530,32'd16625,32'd16720,32'd16815,32'd16910,32'd17005,32'd17100,32'd17195,32'd17290,32'd17385,32'd17480,32'd17575,32'd17670,32'd17765,32'd17860,32'd17955,32'd18050,32'd18145,32'd18240,32'd18335,32'd18430,32'd18525,32'd18620,32'd18715,32'd18810,32'd18905,32'd19000,32'd19095,32'd19190,32'd19285,32'd19380,32'd19475,32'd19570,32'd19665,32'd19760,32'd19855,32'd19950,32'd20045,32'd20140,32'd20235,32'd20330,32'd20425,32'd20520,32'd20615,32'd20710,32'd20805,32'd20900,32'd20995,32'd21090,32'd21185,32'd21280,32'd21375,32'd21470,32'd21565,32'd21660,32'd21755,32'd21850,32'd21945,32'd22040,32'd22135,32'd22230,32'd22325,32'd22420,32'd22515,32'd22610,32'd22705,32'd22800,32'd22895,32'd22990,32'd23085,32'd23180,32'd23275,32'd23370,32'd23465,32'd23560,32'd23655,32'd23750,32'd23845,32'd23940,32'd24035,32'd24130,32'd24225,32'd24320,32'd24415,32'd24510,32'd24605,32'd24700,32'd24795,32'd24890,32'd24985,32'd25080,32'd25175,32'd25270,32'd25365,32'd25460,32'd25555,32'd25650,32'd25745,32'd25840,32'd25935,32'd26030,32'd26125,32'd26220,32'd26315,32'd26410,32'd26505,32'd26600,32'd26695,32'd26790,32'd26885,32'd26980,32'd27075,32'd27170,32'd27265,32'd27360,32'd27455,32'd27550,32'd27645,32'd27740,32'd27835,32'd27930,32'd28025,32'd28120,32'd28215,32'd28310,32'd28405,32'd28500,32'd28595,32'd28690,32'd28785,32'd28880,32'd28975,32'd29070,32'd29165,32'd29260,32'd29355,32'd29450,32'd29545,32'd29640,32'd29735,32'd29830,32'd29925,32'd30020,32'd30115,32'd30210,32'd30305,32'd30400,32'd30495,32'd30590,32'd30685,32'd30780,32'd30875,32'd30970,32'd31065,32'd31160,32'd31255,32'd31350,32'd31445,32'd31540,32'd31635,32'd31730,32'd31825,32'd31920,32'd32015,32'd32110,32'd32205,32'd32300,32'd32395,32'd32490,32'd32585,32'd32680,32'd32775,32'd32870,32'd32965,32'd33060,32'd33155,32'd33250,32'd33345,32'd33440,32'd33535,32'd33630,32'd33725,32'd33820,32'd33915,32'd34010,32'd34105,32'd34200,32'd34295,32'd34390,32'd34485,32'd34580,32'd34675,32'd34770,32'd34865,32'd34960,32'd35055,32'd35150,32'd35245,32'd35340,32'd35435,32'd35530,32'd35625,32'd35720,32'd35815,32'd35910,32'd36005,32'd36100,32'd36195,32'd36290,32'd36385,32'd36480,32'd36575,32'd36670,32'd36765,32'd36860,32'd36955,32'd37050,32'd37145,32'd37240,32'd37335,32'd37430,32'd37525,32'd37620,32'd37715,32'd37810,32'd37905 };matrix[96]='{32'd0,32'd96,32'd192,32'd288,32'd384,32'd480,32'd576,32'd672,32'd768,32'd864,32'd960,32'd1056,32'd1152,32'd1248,32'd1344,32'd1440,32'd1536,32'd1632,32'd1728,32'd1824,32'd1920,32'd2016,32'd2112,32'd2208,32'd2304,32'd2400,32'd2496,32'd2592,32'd2688,32'd2784,32'd2880,32'd2976,32'd3072,32'd3168,32'd3264,32'd3360,32'd3456,32'd3552,32'd3648,32'd3744,32'd3840,32'd3936,32'd4032,32'd4128,32'd4224,32'd4320,32'd4416,32'd4512,32'd4608,32'd4704,32'd4800,32'd4896,32'd4992,32'd5088,32'd5184,32'd5280,32'd5376,32'd5472,32'd5568,32'd5664,32'd5760,32'd5856,32'd5952,32'd6048,32'd6144,32'd6240,32'd6336,32'd6432,32'd6528,32'd6624,32'd6720,32'd6816,32'd6912,32'd7008,32'd7104,32'd7200,32'd7296,32'd7392,32'd7488,32'd7584,32'd7680,32'd7776,32'd7872,32'd7968,32'd8064,32'd8160,32'd8256,32'd8352,32'd8448,32'd8544,32'd8640,32'd8736,32'd8832,32'd8928,32'd9024,32'd9120,32'd9216,32'd9312,32'd9408,32'd9504,32'd9600,32'd9696,32'd9792,32'd9888,32'd9984,32'd10080,32'd10176,32'd10272,32'd10368,32'd10464,32'd10560,32'd10656,32'd10752,32'd10848,32'd10944,32'd11040,32'd11136,32'd11232,32'd11328,32'd11424,32'd11520,32'd11616,32'd11712,32'd11808,32'd11904,32'd12000,32'd12096,32'd12192,32'd12288,32'd12384,32'd12480,32'd12576,32'd12672,32'd12768,32'd12864,32'd12960,32'd13056,32'd13152,32'd13248,32'd13344,32'd13440,32'd13536,32'd13632,32'd13728,32'd13824,32'd13920,32'd14016,32'd14112,32'd14208,32'd14304,32'd14400,32'd14496,32'd14592,32'd14688,32'd14784,32'd14880,32'd14976,32'd15072,32'd15168,32'd15264,32'd15360,32'd15456,32'd15552,32'd15648,32'd15744,32'd15840,32'd15936,32'd16032,32'd16128,32'd16224,32'd16320,32'd16416,32'd16512,32'd16608,32'd16704,32'd16800,32'd16896,32'd16992,32'd17088,32'd17184,32'd17280,32'd17376,32'd17472,32'd17568,32'd17664,32'd17760,32'd17856,32'd17952,32'd18048,32'd18144,32'd18240,32'd18336,32'd18432,32'd18528,32'd18624,32'd18720,32'd18816,32'd18912,32'd19008,32'd19104,32'd19200,32'd19296,32'd19392,32'd19488,32'd19584,32'd19680,32'd19776,32'd19872,32'd19968,32'd20064,32'd20160,32'd20256,32'd20352,32'd20448,32'd20544,32'd20640,32'd20736,32'd20832,32'd20928,32'd21024,32'd21120,32'd21216,32'd21312,32'd21408,32'd21504,32'd21600,32'd21696,32'd21792,32'd21888,32'd21984,32'd22080,32'd22176,32'd22272,32'd22368,32'd22464,32'd22560,32'd22656,32'd22752,32'd22848,32'd22944,32'd23040,32'd23136,32'd23232,32'd23328,32'd23424,32'd23520,32'd23616,32'd23712,32'd23808,32'd23904,32'd24000,32'd24096,32'd24192,32'd24288,32'd24384,32'd24480,32'd24576,32'd24672,32'd24768,32'd24864,32'd24960,32'd25056,32'd25152,32'd25248,32'd25344,32'd25440,32'd25536,32'd25632,32'd25728,32'd25824,32'd25920,32'd26016,32'd26112,32'd26208,32'd26304,32'd26400,32'd26496,32'd26592,32'd26688,32'd26784,32'd26880,32'd26976,32'd27072,32'd27168,32'd27264,32'd27360,32'd27456,32'd27552,32'd27648,32'd27744,32'd27840,32'd27936,32'd28032,32'd28128,32'd28224,32'd28320,32'd28416,32'd28512,32'd28608,32'd28704,32'd28800,32'd28896,32'd28992,32'd29088,32'd29184,32'd29280,32'd29376,32'd29472,32'd29568,32'd29664,32'd29760,32'd29856,32'd29952,32'd30048,32'd30144,32'd30240,32'd30336,32'd30432,32'd30528,32'd30624,32'd30720,32'd30816,32'd30912,32'd31008,32'd31104,32'd31200,32'd31296,32'd31392,32'd31488,32'd31584,32'd31680,32'd31776,32'd31872,32'd31968,32'd32064,32'd32160,32'd32256,32'd32352,32'd32448,32'd32544,32'd32640,32'd32736,32'd32832,32'd32928,32'd33024,32'd33120,32'd33216,32'd33312,32'd33408,32'd33504,32'd33600,32'd33696,32'd33792,32'd33888,32'd33984,32'd34080,32'd34176,32'd34272,32'd34368,32'd34464,32'd34560,32'd34656,32'd34752,32'd34848,32'd34944,32'd35040,32'd35136,32'd35232,32'd35328,32'd35424,32'd35520,32'd35616,32'd35712,32'd35808,32'd35904,32'd36000,32'd36096,32'd36192,32'd36288,32'd36384,32'd36480,32'd36576,32'd36672,32'd36768,32'd36864,32'd36960,32'd37056,32'd37152,32'd37248,32'd37344,32'd37440,32'd37536,32'd37632,32'd37728,32'd37824,32'd37920,32'd38016,32'd38112,32'd38208,32'd38304 };matrix[97]='{32'd0,32'd97,32'd194,32'd291,32'd388,32'd485,32'd582,32'd679,32'd776,32'd873,32'd970,32'd1067,32'd1164,32'd1261,32'd1358,32'd1455,32'd1552,32'd1649,32'd1746,32'd1843,32'd1940,32'd2037,32'd2134,32'd2231,32'd2328,32'd2425,32'd2522,32'd2619,32'd2716,32'd2813,32'd2910,32'd3007,32'd3104,32'd3201,32'd3298,32'd3395,32'd3492,32'd3589,32'd3686,32'd3783,32'd3880,32'd3977,32'd4074,32'd4171,32'd4268,32'd4365,32'd4462,32'd4559,32'd4656,32'd4753,32'd4850,32'd4947,32'd5044,32'd5141,32'd5238,32'd5335,32'd5432,32'd5529,32'd5626,32'd5723,32'd5820,32'd5917,32'd6014,32'd6111,32'd6208,32'd6305,32'd6402,32'd6499,32'd6596,32'd6693,32'd6790,32'd6887,32'd6984,32'd7081,32'd7178,32'd7275,32'd7372,32'd7469,32'd7566,32'd7663,32'd7760,32'd7857,32'd7954,32'd8051,32'd8148,32'd8245,32'd8342,32'd8439,32'd8536,32'd8633,32'd8730,32'd8827,32'd8924,32'd9021,32'd9118,32'd9215,32'd9312,32'd9409,32'd9506,32'd9603,32'd9700,32'd9797,32'd9894,32'd9991,32'd10088,32'd10185,32'd10282,32'd10379,32'd10476,32'd10573,32'd10670,32'd10767,32'd10864,32'd10961,32'd11058,32'd11155,32'd11252,32'd11349,32'd11446,32'd11543,32'd11640,32'd11737,32'd11834,32'd11931,32'd12028,32'd12125,32'd12222,32'd12319,32'd12416,32'd12513,32'd12610,32'd12707,32'd12804,32'd12901,32'd12998,32'd13095,32'd13192,32'd13289,32'd13386,32'd13483,32'd13580,32'd13677,32'd13774,32'd13871,32'd13968,32'd14065,32'd14162,32'd14259,32'd14356,32'd14453,32'd14550,32'd14647,32'd14744,32'd14841,32'd14938,32'd15035,32'd15132,32'd15229,32'd15326,32'd15423,32'd15520,32'd15617,32'd15714,32'd15811,32'd15908,32'd16005,32'd16102,32'd16199,32'd16296,32'd16393,32'd16490,32'd16587,32'd16684,32'd16781,32'd16878,32'd16975,32'd17072,32'd17169,32'd17266,32'd17363,32'd17460,32'd17557,32'd17654,32'd17751,32'd17848,32'd17945,32'd18042,32'd18139,32'd18236,32'd18333,32'd18430,32'd18527,32'd18624,32'd18721,32'd18818,32'd18915,32'd19012,32'd19109,32'd19206,32'd19303,32'd19400,32'd19497,32'd19594,32'd19691,32'd19788,32'd19885,32'd19982,32'd20079,32'd20176,32'd20273,32'd20370,32'd20467,32'd20564,32'd20661,32'd20758,32'd20855,32'd20952,32'd21049,32'd21146,32'd21243,32'd21340,32'd21437,32'd21534,32'd21631,32'd21728,32'd21825,32'd21922,32'd22019,32'd22116,32'd22213,32'd22310,32'd22407,32'd22504,32'd22601,32'd22698,32'd22795,32'd22892,32'd22989,32'd23086,32'd23183,32'd23280,32'd23377,32'd23474,32'd23571,32'd23668,32'd23765,32'd23862,32'd23959,32'd24056,32'd24153,32'd24250,32'd24347,32'd24444,32'd24541,32'd24638,32'd24735,32'd24832,32'd24929,32'd25026,32'd25123,32'd25220,32'd25317,32'd25414,32'd25511,32'd25608,32'd25705,32'd25802,32'd25899,32'd25996,32'd26093,32'd26190,32'd26287,32'd26384,32'd26481,32'd26578,32'd26675,32'd26772,32'd26869,32'd26966,32'd27063,32'd27160,32'd27257,32'd27354,32'd27451,32'd27548,32'd27645,32'd27742,32'd27839,32'd27936,32'd28033,32'd28130,32'd28227,32'd28324,32'd28421,32'd28518,32'd28615,32'd28712,32'd28809,32'd28906,32'd29003,32'd29100,32'd29197,32'd29294,32'd29391,32'd29488,32'd29585,32'd29682,32'd29779,32'd29876,32'd29973,32'd30070,32'd30167,32'd30264,32'd30361,32'd30458,32'd30555,32'd30652,32'd30749,32'd30846,32'd30943,32'd31040,32'd31137,32'd31234,32'd31331,32'd31428,32'd31525,32'd31622,32'd31719,32'd31816,32'd31913,32'd32010,32'd32107,32'd32204,32'd32301,32'd32398,32'd32495,32'd32592,32'd32689,32'd32786,32'd32883,32'd32980,32'd33077,32'd33174,32'd33271,32'd33368,32'd33465,32'd33562,32'd33659,32'd33756,32'd33853,32'd33950,32'd34047,32'd34144,32'd34241,32'd34338,32'd34435,32'd34532,32'd34629,32'd34726,32'd34823,32'd34920,32'd35017,32'd35114,32'd35211,32'd35308,32'd35405,32'd35502,32'd35599,32'd35696,32'd35793,32'd35890,32'd35987,32'd36084,32'd36181,32'd36278,32'd36375,32'd36472,32'd36569,32'd36666,32'd36763,32'd36860,32'd36957,32'd37054,32'd37151,32'd37248,32'd37345,32'd37442,32'd37539,32'd37636,32'd37733,32'd37830,32'd37927,32'd38024,32'd38121,32'd38218,32'd38315,32'd38412,32'd38509,32'd38606,32'd38703 };matrix[98]='{32'd0,32'd98,32'd196,32'd294,32'd392,32'd490,32'd588,32'd686,32'd784,32'd882,32'd980,32'd1078,32'd1176,32'd1274,32'd1372,32'd1470,32'd1568,32'd1666,32'd1764,32'd1862,32'd1960,32'd2058,32'd2156,32'd2254,32'd2352,32'd2450,32'd2548,32'd2646,32'd2744,32'd2842,32'd2940,32'd3038,32'd3136,32'd3234,32'd3332,32'd3430,32'd3528,32'd3626,32'd3724,32'd3822,32'd3920,32'd4018,32'd4116,32'd4214,32'd4312,32'd4410,32'd4508,32'd4606,32'd4704,32'd4802,32'd4900,32'd4998,32'd5096,32'd5194,32'd5292,32'd5390,32'd5488,32'd5586,32'd5684,32'd5782,32'd5880,32'd5978,32'd6076,32'd6174,32'd6272,32'd6370,32'd6468,32'd6566,32'd6664,32'd6762,32'd6860,32'd6958,32'd7056,32'd7154,32'd7252,32'd7350,32'd7448,32'd7546,32'd7644,32'd7742,32'd7840,32'd7938,32'd8036,32'd8134,32'd8232,32'd8330,32'd8428,32'd8526,32'd8624,32'd8722,32'd8820,32'd8918,32'd9016,32'd9114,32'd9212,32'd9310,32'd9408,32'd9506,32'd9604,32'd9702,32'd9800,32'd9898,32'd9996,32'd10094,32'd10192,32'd10290,32'd10388,32'd10486,32'd10584,32'd10682,32'd10780,32'd10878,32'd10976,32'd11074,32'd11172,32'd11270,32'd11368,32'd11466,32'd11564,32'd11662,32'd11760,32'd11858,32'd11956,32'd12054,32'd12152,32'd12250,32'd12348,32'd12446,32'd12544,32'd12642,32'd12740,32'd12838,32'd12936,32'd13034,32'd13132,32'd13230,32'd13328,32'd13426,32'd13524,32'd13622,32'd13720,32'd13818,32'd13916,32'd14014,32'd14112,32'd14210,32'd14308,32'd14406,32'd14504,32'd14602,32'd14700,32'd14798,32'd14896,32'd14994,32'd15092,32'd15190,32'd15288,32'd15386,32'd15484,32'd15582,32'd15680,32'd15778,32'd15876,32'd15974,32'd16072,32'd16170,32'd16268,32'd16366,32'd16464,32'd16562,32'd16660,32'd16758,32'd16856,32'd16954,32'd17052,32'd17150,32'd17248,32'd17346,32'd17444,32'd17542,32'd17640,32'd17738,32'd17836,32'd17934,32'd18032,32'd18130,32'd18228,32'd18326,32'd18424,32'd18522,32'd18620,32'd18718,32'd18816,32'd18914,32'd19012,32'd19110,32'd19208,32'd19306,32'd19404,32'd19502,32'd19600,32'd19698,32'd19796,32'd19894,32'd19992,32'd20090,32'd20188,32'd20286,32'd20384,32'd20482,32'd20580,32'd20678,32'd20776,32'd20874,32'd20972,32'd21070,32'd21168,32'd21266,32'd21364,32'd21462,32'd21560,32'd21658,32'd21756,32'd21854,32'd21952,32'd22050,32'd22148,32'd22246,32'd22344,32'd22442,32'd22540,32'd22638,32'd22736,32'd22834,32'd22932,32'd23030,32'd23128,32'd23226,32'd23324,32'd23422,32'd23520,32'd23618,32'd23716,32'd23814,32'd23912,32'd24010,32'd24108,32'd24206,32'd24304,32'd24402,32'd24500,32'd24598,32'd24696,32'd24794,32'd24892,32'd24990,32'd25088,32'd25186,32'd25284,32'd25382,32'd25480,32'd25578,32'd25676,32'd25774,32'd25872,32'd25970,32'd26068,32'd26166,32'd26264,32'd26362,32'd26460,32'd26558,32'd26656,32'd26754,32'd26852,32'd26950,32'd27048,32'd27146,32'd27244,32'd27342,32'd27440,32'd27538,32'd27636,32'd27734,32'd27832,32'd27930,32'd28028,32'd28126,32'd28224,32'd28322,32'd28420,32'd28518,32'd28616,32'd28714,32'd28812,32'd28910,32'd29008,32'd29106,32'd29204,32'd29302,32'd29400,32'd29498,32'd29596,32'd29694,32'd29792,32'd29890,32'd29988,32'd30086,32'd30184,32'd30282,32'd30380,32'd30478,32'd30576,32'd30674,32'd30772,32'd30870,32'd30968,32'd31066,32'd31164,32'd31262,32'd31360,32'd31458,32'd31556,32'd31654,32'd31752,32'd31850,32'd31948,32'd32046,32'd32144,32'd32242,32'd32340,32'd32438,32'd32536,32'd32634,32'd32732,32'd32830,32'd32928,32'd33026,32'd33124,32'd33222,32'd33320,32'd33418,32'd33516,32'd33614,32'd33712,32'd33810,32'd33908,32'd34006,32'd34104,32'd34202,32'd34300,32'd34398,32'd34496,32'd34594,32'd34692,32'd34790,32'd34888,32'd34986,32'd35084,32'd35182,32'd35280,32'd35378,32'd35476,32'd35574,32'd35672,32'd35770,32'd35868,32'd35966,32'd36064,32'd36162,32'd36260,32'd36358,32'd36456,32'd36554,32'd36652,32'd36750,32'd36848,32'd36946,32'd37044,32'd37142,32'd37240,32'd37338,32'd37436,32'd37534,32'd37632,32'd37730,32'd37828,32'd37926,32'd38024,32'd38122,32'd38220,32'd38318,32'd38416,32'd38514,32'd38612,32'd38710,32'd38808,32'd38906,32'd39004,32'd39102 };matrix[99]='{32'd0,32'd99,32'd198,32'd297,32'd396,32'd495,32'd594,32'd693,32'd792,32'd891,32'd990,32'd1089,32'd1188,32'd1287,32'd1386,32'd1485,32'd1584,32'd1683,32'd1782,32'd1881,32'd1980,32'd2079,32'd2178,32'd2277,32'd2376,32'd2475,32'd2574,32'd2673,32'd2772,32'd2871,32'd2970,32'd3069,32'd3168,32'd3267,32'd3366,32'd3465,32'd3564,32'd3663,32'd3762,32'd3861,32'd3960,32'd4059,32'd4158,32'd4257,32'd4356,32'd4455,32'd4554,32'd4653,32'd4752,32'd4851,32'd4950,32'd5049,32'd5148,32'd5247,32'd5346,32'd5445,32'd5544,32'd5643,32'd5742,32'd5841,32'd5940,32'd6039,32'd6138,32'd6237,32'd6336,32'd6435,32'd6534,32'd6633,32'd6732,32'd6831,32'd6930,32'd7029,32'd7128,32'd7227,32'd7326,32'd7425,32'd7524,32'd7623,32'd7722,32'd7821,32'd7920,32'd8019,32'd8118,32'd8217,32'd8316,32'd8415,32'd8514,32'd8613,32'd8712,32'd8811,32'd8910,32'd9009,32'd9108,32'd9207,32'd9306,32'd9405,32'd9504,32'd9603,32'd9702,32'd9801,32'd9900,32'd9999,32'd10098,32'd10197,32'd10296,32'd10395,32'd10494,32'd10593,32'd10692,32'd10791,32'd10890,32'd10989,32'd11088,32'd11187,32'd11286,32'd11385,32'd11484,32'd11583,32'd11682,32'd11781,32'd11880,32'd11979,32'd12078,32'd12177,32'd12276,32'd12375,32'd12474,32'd12573,32'd12672,32'd12771,32'd12870,32'd12969,32'd13068,32'd13167,32'd13266,32'd13365,32'd13464,32'd13563,32'd13662,32'd13761,32'd13860,32'd13959,32'd14058,32'd14157,32'd14256,32'd14355,32'd14454,32'd14553,32'd14652,32'd14751,32'd14850,32'd14949,32'd15048,32'd15147,32'd15246,32'd15345,32'd15444,32'd15543,32'd15642,32'd15741,32'd15840,32'd15939,32'd16038,32'd16137,32'd16236,32'd16335,32'd16434,32'd16533,32'd16632,32'd16731,32'd16830,32'd16929,32'd17028,32'd17127,32'd17226,32'd17325,32'd17424,32'd17523,32'd17622,32'd17721,32'd17820,32'd17919,32'd18018,32'd18117,32'd18216,32'd18315,32'd18414,32'd18513,32'd18612,32'd18711,32'd18810,32'd18909,32'd19008,32'd19107,32'd19206,32'd19305,32'd19404,32'd19503,32'd19602,32'd19701,32'd19800,32'd19899,32'd19998,32'd20097,32'd20196,32'd20295,32'd20394,32'd20493,32'd20592,32'd20691,32'd20790,32'd20889,32'd20988,32'd21087,32'd21186,32'd21285,32'd21384,32'd21483,32'd21582,32'd21681,32'd21780,32'd21879,32'd21978,32'd22077,32'd22176,32'd22275,32'd22374,32'd22473,32'd22572,32'd22671,32'd22770,32'd22869,32'd22968,32'd23067,32'd23166,32'd23265,32'd23364,32'd23463,32'd23562,32'd23661,32'd23760,32'd23859,32'd23958,32'd24057,32'd24156,32'd24255,32'd24354,32'd24453,32'd24552,32'd24651,32'd24750,32'd24849,32'd24948,32'd25047,32'd25146,32'd25245,32'd25344,32'd25443,32'd25542,32'd25641,32'd25740,32'd25839,32'd25938,32'd26037,32'd26136,32'd26235,32'd26334,32'd26433,32'd26532,32'd26631,32'd26730,32'd26829,32'd26928,32'd27027,32'd27126,32'd27225,32'd27324,32'd27423,32'd27522,32'd27621,32'd27720,32'd27819,32'd27918,32'd28017,32'd28116,32'd28215,32'd28314,32'd28413,32'd28512,32'd28611,32'd28710,32'd28809,32'd28908,32'd29007,32'd29106,32'd29205,32'd29304,32'd29403,32'd29502,32'd29601,32'd29700,32'd29799,32'd29898,32'd29997,32'd30096,32'd30195,32'd30294,32'd30393,32'd30492,32'd30591,32'd30690,32'd30789,32'd30888,32'd30987,32'd31086,32'd31185,32'd31284,32'd31383,32'd31482,32'd31581,32'd31680,32'd31779,32'd31878,32'd31977,32'd32076,32'd32175,32'd32274,32'd32373,32'd32472,32'd32571,32'd32670,32'd32769,32'd32868,32'd32967,32'd33066,32'd33165,32'd33264,32'd33363,32'd33462,32'd33561,32'd33660,32'd33759,32'd33858,32'd33957,32'd34056,32'd34155,32'd34254,32'd34353,32'd34452,32'd34551,32'd34650,32'd34749,32'd34848,32'd34947,32'd35046,32'd35145,32'd35244,32'd35343,32'd35442,32'd35541,32'd35640,32'd35739,32'd35838,32'd35937,32'd36036,32'd36135,32'd36234,32'd36333,32'd36432,32'd36531,32'd36630,32'd36729,32'd36828,32'd36927,32'd37026,32'd37125,32'd37224,32'd37323,32'd37422,32'd37521,32'd37620,32'd37719,32'd37818,32'd37917,32'd38016,32'd38115,32'd38214,32'd38313,32'd38412,32'd38511,32'd38610,32'd38709,32'd38808,32'd38907,32'd39006,32'd39105,32'd39204,32'd39303,32'd39402,32'd39501 };
    vector='{32'd0,32'd1,32'd2,32'd3,32'd4,32'd5,32'd6,32'd7,32'd8,32'd9,32'd10,32'd11,32'd12,32'd13,32'd14,32'd15,32'd16,32'd17,32'd18,32'd19,32'd20,32'd21,32'd22,32'd23,32'd24,32'd25,32'd26,32'd27,32'd28,32'd29,32'd30,32'd31,32'd32,32'd33,32'd34,32'd35,32'd36,32'd37,32'd38,32'd39,32'd40,32'd41,32'd42,32'd43,32'd44,32'd45,32'd46,32'd47,32'd48,32'd49,32'd50,32'd51,32'd52,32'd53,32'd54,32'd55,32'd56,32'd57,32'd58,32'd59,32'd60,32'd61,32'd62,32'd63,32'd64,32'd65,32'd66,32'd67,32'd68,32'd69,32'd70,32'd71,32'd72,32'd73,32'd74,32'd75,32'd76,32'd77,32'd78,32'd79,32'd80,32'd81,32'd82,32'd83,32'd84,32'd85,32'd86,32'd87,32'd88,32'd89,32'd90,32'd91,32'd92,32'd93,32'd94,32'd95,32'd96,32'd97,32'd98,32'd99 };
    //======================================
    
    // Apply stimulus
    #10;
    
    // Display the result
    $display("Result: %d", result);
    
    // End simulation
    #10$finish;
  end
  
endmodule
