`include "vmvmb.sv"

    //========== this a testbench driven by 6 data in a group from python gen txt =========
    module tb;
    logic signed [31:0] x[0:99];
    logic signed [31:0] Wx[0:99][0:399];
    logic signed [31:0] h_prev[0:99];
    logic signed [31:0] Wh[0:99][0:399];
    logic signed [31:0] b[0:399];
    logic signed [31:0] A[0:399];
    vmvmb dut(
        x,Wx,h_prev,Wh,b,A
    );
    initial begin
        $fsdbDumpfile("tb_6data.fsdb");
        $fsdbDumpvars("+all");
    end
    initial begin
    #10;
    x='{32'd2330,32'd2047,32'd-49,32'd-2961,32'd-54,32'd480,32'd-1728,32'd-1111,32'd2214,32'd-9575,32'd993,32'd4052,32'd-3518,32'd-3215,32'd430,32'd2386,32'd-1245,32'd1867,32'd330,32'd1953,32'd-4775,32'd3457,32'd-2783,32'd1555,32'd2954,32'd-2602,32'd-1588,32'd2763,32'd-4379,32'd6376,32'd-815,32'd3034,32'd-2458,32'd-523,32'd-392,32'd-2536,32'd-1047,32'd-1115,32'd516,32'd-577,32'd12,32'd4538,32'd-1199,32'd2971,32'd-2912,32'd3154,32'd4538,32'd2980,32'd-897,32'd1973,32'd-2158,32'd1784,32'd4509,32'd-113,32'd-3269,32'd-2697,32'd-4052,32'd-2844,32'd-5234,32'd-1096,32'd-203,32'd1050,32'd3071,32'd4003,32'd-777,32'd2778,32'd1890,32'd298,32'd178,32'd-4899,32'd1799,32'd-2454,32'd5170,32'd-3618,32'd-5302,32'd-1679,32'd-123,32'd3493,32'd3388,32'd5361,32'd-754,32'd3559,32'd-3815,32'd4370,32'd-1448,32'd-4143,32'd-720,32'd-1811,32'd1986,32'd-2951,32'd563,32'd1052,32'd745,32'd2186,32'd4262,32'd-846,32'd-1157,32'd262,32'd249,32'd-4721};
    h_prev='{32'd0,32'd7531,32'd-31,32'd536,32'd5,32'd-11,32'd-345,32'd-3206,32'd655,32'd1300,32'd-150,32'd-1578,32'd545,32'd3005,32'd0,32'd1619,32'd6694,32'd1093,32'd-451,32'd43,32'd49,32'd5,32'd-690,32'd2,32'd0,32'd-3087,32'd0,32'd4420,32'd-297,32'd-634,32'd386,32'd6774,32'd253,32'd-4078,32'd43,32'd-16,32'd8,32'd596,32'd-6244,32'd-5694,32'd-124,32'd6721,32'd-6314,32'd-7489,32'd-4378,32'd7047,32'd1937,32'd576,32'd-345,32'd-1097,32'd7322,32'd-7510,32'd443,32'd6400,32'd-310,32'd-1839,32'd-3803,32'd-35,32'd-647,32'd6255,32'd615,32'd-26,32'd-3230,32'd398,32'd-848,32'd0,32'd-2154,32'd7441,32'd-576,32'd-57,32'd257,32'd-7257,32'd-25,32'd-5635,32'd1,32'd-56,32'd-7604,32'd5018,32'd873,32'd-4056,32'd9,32'd7315,32'd-107,32'd-7266,32'd0,32'd5227,32'd-53,32'd1492,32'd-638,32'd6954,32'd-2,32'd-978,32'd-278,32'd4962,32'd926,32'd-3516,32'd628,32'd41,32'd86,32'd-5108};
    b='{32'd2325,32'd-16591,32'd-5761,32'd-12939,32'd-2268,32'd8706,32'd-14824,32'd-7407,32'd1971,32'd-6577,32'd-8862,32'd3022,32'd1065,32'd-15878,32'd-7822,32'd-8212,32'd-12353,32'd13,32'd-2687,32'd-8769,32'd816,32'd-7163,32'd-5839,32'd-8320,32'd-1706,32'd-406,32'd-5483,32'd-1447,32'd-5449,32'd-2780,32'd-4860,32'd-11816,32'd-14082,32'd-8930,32'd30156,32'd-7968,32'd13271,32'd-3193,32'd-9770,32'd-15302,32'd1127,32'd-25781,32'd23574,32'd-13740,32'd-2033,32'd-680,32'd-20019,32'd2381,32'd-14257,32'd33281,32'd-10078,32'd-16669,32'd5009,32'd13349,32'd5454,32'd16015,32'd-8173,32'd911,32'd-10722,32'd16494,32'd-1926,32'd-9931,32'd-13828,32'd1466,32'd-125,32'd-4362,32'd3579,32'd-21718,32'd42,32'd-3796,32'd25058,32'd-19199,32'd-13105,32'd-16464,32'd-3146,32'd-6401,32'd-6411,32'd-9160,32'd36113,32'd1428,32'd-5668,32'd-23535,32'd-12744,32'd-22968,32'd2939,32'd-15312,32'd-1862,32'd-7666,32'd8647,32'd1607,32'd-6269,32'd-16708,32'd-11044,32'd-22578,32'd-25273,32'd-7495,32'd2443,32'd-21816,32'd-8652,32'd-11708,32'd-2158,32'd5581,32'd-11201,32'd4299,32'd5498,32'd-12734,32'd-22167,32'd-13652,32'd12119,32'd-9165,32'd-7456,32'd2143,32'd875,32'd1092,32'd-1405,32'd11923,32'd-6508,32'd-10478,32'd-10673,32'd3737,32'd15556,32'd4450,32'd-2470,32'd-2175,32'd-7202,32'd9233,32'd-4433,32'd-5571,32'd1979,32'd-5434,32'd-6669,32'd-9204,32'd10234,32'd9111,32'd35332,32'd15410,32'd14570,32'd8989,32'd5957,32'd-7246,32'd-5693,32'd-621,32'd3356,32'd15781,32'd-6186,32'd2531,32'd22500,32'd10458,32'd2587,32'd-2441,32'd-10810,32'd-20,32'd9965,32'd-4663,32'd-13378,32'd-7387,32'd13769,32'd-17402,32'd-12050,32'd10888,32'd-11406,32'd-7739,32'd2778,32'd-18427,32'd4763,32'd-8984,32'd-13447,32'd-11982,32'd-18017,32'd16992,32'd5170,32'd-9428,32'd5800,32'd-10996,32'd10546,32'd2462,32'd-520,32'd2225,32'd6923,32'd18095,32'd13564,32'd18623,32'd-12714,32'd5654,32'd15625,32'd909,32'd-14062,32'd7416,32'd-11494,32'd21191,32'd-10449,32'd-3354,32'd-5722,32'd28671,32'd19765,32'd-7260,32'd12441,32'd921,32'd13,32'd4580,32'd-3010,32'd11337,32'd-35,32'd-582,32'd-1089,32'd4050,32'd5527,32'd7456,32'd-5185,32'd-2135,32'd9526,32'd-8574,32'd-12910,32'd12626,32'd9956,32'd-7827,32'd-3574,32'd637,32'd-10634,32'd-10566,32'd481,32'd-3547,32'd-9575,32'd-3740,32'd-5263,32'd-5961,32'd-8510,32'd581,32'd3078,32'd-10800,32'd-6459,32'd6196,32'd13212,32'd6865,32'd-20234,32'd-5776,32'd-22832,32'd-262,32'd14921,32'd12695,32'd-2697,32'd11035,32'd-8994,32'd12646,32'd-1105,32'd5795,32'd4804,32'd-3356,32'd-643,32'd-25292,32'd16640,32'd10166,32'd-4919,32'd-7661,32'd-15009,32'd-7006,32'd-5561,32'd-1893,32'd-1473,32'd-23085,32'd-15087,32'd-5205,32'd24472,32'd-3608,32'd7495,32'd-12607,32'd-6894,32'd5776,32'd1760,32'd-3903,32'd-26796,32'd3188,32'd-6088,32'd8295,32'd-4401,32'd5615,32'd612,32'd11337,32'd-27773,32'd-4133,32'd-6674,32'd9150,32'd-2237,32'd21113,32'd-863,32'd8994,32'd-5307,32'd4187,32'd-18476,32'd103,32'd-16796,32'd25820,32'd1778,32'd7016,32'd8984,32'd930,32'd-6279,32'd12656,32'd-8710,32'd13720,32'd-15244,32'd26035,32'd-34160,32'd2376,32'd-1462,32'd-34628,32'd-2639,32'd10302,32'd2487,32'd-7680,32'd8588,32'd-2191,32'd-16396,32'd15078,32'd18701,32'd15185,32'd23945,32'd-715,32'd-7021,32'd-25820,32'd-26542,32'd-5571,32'd-11767,32'd-4133,32'd-7934,32'd-3090,32'd-1916,32'd-7265,32'd4565,32'd6542,32'd-9467,32'd18251,32'd11855,32'd15849,32'd8735,32'd-8808,32'd6689,32'd-10859,32'd13847,32'd16093,32'd4677,32'd20195,32'd6220,32'd4038,32'd11347,32'd7685,32'd26074,32'd3815,32'd-10781,32'd12343,32'd22519,32'd20742,32'd-2722,32'd12509,32'd-6474,32'd14277,32'd-896,32'd-34160,32'd6064,32'd-659,32'd-14785,32'd6728,32'd12919,32'd7866,32'd16679,32'd-25976,32'd-11464,32'd22382,32'd-20390,32'd-21054,32'd2895,32'd343,32'd-11220,32'd13896,32'd-15517,32'd8417,32'd16220,32'd10205,32'd22402,32'd-1508,32'd-4157,32'd27792,32'd-2673,32'd24042,32'd-6416,32'd17197,32'd-10869,32'd-672,32'd-3002,32'd-35761,32'd-6186,32'd6982,32'd9575,32'd-20820,32'd16318,32'd2413,32'd-4609,32'd27324,32'd-9907,32'd15625};
    Wx[0]='{32'd1748,32'd-2391,32'd-84,32'd-2595,32'd-209,32'd1027,32'd-4772,32'd-1782,32'd-413,32'd-1520,32'd45,32'd-1872,32'd-1966,32'd-1979,32'd-526,32'd5195,32'd2395,32'd-995,32'd3034,32'd159,32'd374,32'd-450,32'd-1140,32'd861,32'd698,32'd3110,32'd509,32'd560,32'd-3002,32'd-2878,32'd124,32'd-6796,32'd813,32'd3708,32'd-253,32'd-2749,32'd548,32'd1571,32'd1977,32'd-2110,32'd273,32'd4450,32'd2651,32'd4565,32'd8852,32'd-3347,32'd-1206,32'd3969,32'd-1697,32'd1602,32'd-2812,32'd558,32'd-1474,32'd4772,32'd1049,32'd-2697,32'd-2244,32'd4650,32'd-5063,32'd1347,32'd3984,32'd-2482,32'd-862,32'd-337,32'd-4309,32'd-708,32'd-5053,32'd12568,32'd1018,32'd-1983,32'd-3234,32'd-3654,32'd2120,32'd-8930,32'd2741,32'd2115,32'd1712,32'd-1268,32'd-3627,32'd-4992,32'd1536,32'd-3159,32'd-319,32'd935,32'd109,32'd-3535,32'd426,32'd-294,32'd182,32'd-2978,32'd-2978,32'd2917,32'd-2316,32'd-1596,32'd870,32'd-1390,32'd-2846,32'd-197,32'd1804,32'd-326,32'd1583,32'd6962,32'd-1955,32'd2944,32'd4387,32'd-2283,32'd4411,32'd-5000,32'd3989,32'd2934,32'd1784,32'd-5107,32'd228,32'd-5942,32'd-8730,32'd9541,32'd-2150,32'd6176,32'd2575,32'd2617,32'd-3586,32'd-5991,32'd-4536,32'd5209,32'd-143,32'd7387,32'd-4245,32'd3369,32'd-14296,32'd-2315,32'd3391,32'd-17060,32'd7104,32'd10263,32'd-8037,32'd1678,32'd-416,32'd-1987,32'd28105,32'd3261,32'd3913,32'd5102,32'd9169,32'd-9174,32'd2028,32'd2015,32'd-6606,32'd2050,32'd-2495,32'd3811,32'd9936,32'd1859,32'd2335,32'd4294,32'd565,32'd-4707,32'd-539,32'd-2788,32'd-9370,32'd-4548,32'd-3381,32'd1191,32'd-20722,32'd3979,32'd-2504,32'd1778,32'd2271,32'd-474,32'd2880,32'd1074,32'd-3071,32'd-8071,32'd-2854,32'd2395,32'd2292,32'd-733,32'd-841,32'd-7021,32'd-4082,32'd1253,32'd435,32'd8632,32'd4997,32'd-12705,32'd-972,32'd6191,32'd-2617,32'd2043,32'd1710,32'd-581,32'd1738,32'd14316,32'd-1013,32'd297,32'd-5737,32'd6621,32'd-5258,32'd1318,32'd6606,32'd2980,32'd-1444,32'd-1418,32'd-916,32'd1661,32'd1507,32'd-93,32'd-5585,32'd-5903,32'd-288,32'd-548,32'd-3378,32'd-5424,32'd-5219,32'd-5625,32'd8593,32'd6660,32'd-1472,32'd-5000,32'd-3410,32'd-4416,32'd2408,32'd433,32'd-590,32'd-541,32'd-3034,32'd-3247,32'd-9838,32'd-407,32'd-10341,32'd6596,32'd-441,32'd-3569,32'd2214,32'd1781,32'd1525,32'd-3254,32'd-3762,32'd1170,32'd-3942,32'd-2453,32'd-182,32'd2249,32'd-3850,32'd-3728,32'd6162,32'd-2399,32'd-2829,32'd-3703,32'd272,32'd-522,32'd-4211,32'd1148,32'd-3193,32'd2199,32'd-3359,32'd-2219,32'd-6923,32'd438,32'd342,32'd2124,32'd336,32'd-3952,32'd-686,32'd166,32'd-11054,32'd-650,32'd-6704,32'd422,32'd3620,32'd-2998,32'd3195,32'd1872,32'd-1497,32'd-1053,32'd169,32'd-6333,32'd4965,32'd-3796,32'd-5019,32'd2269,32'd-1610,32'd8442,32'd497,32'd-4912,32'd-5034,32'd-2641,32'd1246,32'd-2156,32'd2364,32'd-1135,32'd-4892,32'd376,32'd4299,32'd2954,32'd1356,32'd3378,32'd-1019,32'd-5283,32'd-485,32'd323,32'd-2773,32'd15,32'd2834,32'd-2497,32'd520,32'd-6713,32'd-7416,32'd2053,32'd5898,32'd78,32'd-6425,32'd-3461,32'd-1616,32'd-4121,32'd385,32'd4965,32'd1895,32'd-9873,32'd1890,32'd137,32'd180,32'd-1066,32'd242,32'd-2509,32'd-4313,32'd514,32'd-5942,32'd1334,32'd-2377,32'd1319,32'd442,32'd-3041,32'd-2205,32'd1828,32'd6313,32'd-5771,32'd4162,32'd7934,32'd2741,32'd-9667,32'd3291,32'd-3044,32'd-5097,32'd-990,32'd-620,32'd-2073,32'd4191,32'd2719,32'd2023,32'd-1494,32'd-6391,32'd-2124,32'd-3437,32'd130,32'd413,32'd-6918,32'd-6210,32'd6098,32'd-2575,32'd6240,32'd2470,32'd-4121,32'd759,32'd4123,32'd-1907,32'd-4995,32'd-8745,32'd1820,32'd-1737,32'd-9316,32'd-3542,32'd-3884,32'd5810,32'd-10664,32'd3352,32'd1601,32'd1304,32'd-4602,32'd1939,32'd4042,32'd2287,32'd1691,32'd6450,32'd-4123,32'd-4870,32'd-1944,32'd2680,32'd-955,32'd2553,32'd12402,32'd-4328,32'd-3818,32'd-3901,32'd13681,32'd-2954,32'd5732,32'd-4650,32'd5253,32'd-911,32'd391};
    Wx[1]='{32'd-2021,32'd792,32'd-446,32'd-1254,32'd3015,32'd2592,32'd-2670,32'd-2197,32'd895,32'd-872,32'd5546,32'd1298,32'd-979,32'd-1141,32'd155,32'd5888,32'd8510,32'd2963,32'd-1262,32'd-963,32'd1883,32'd4477,32'd-2131,32'd2548,32'd3872,32'd3259,32'd1389,32'd1835,32'd-2279,32'd4406,32'd17,32'd3405,32'd-950,32'd2327,32'd-745,32'd1199,32'd-1387,32'd563,32'd-1486,32'd-419,32'd496,32'd-636,32'd-720,32'd5898,32'd-2249,32'd2795,32'd1356,32'd-3088,32'd2056,32'd-2056,32'd-7431,32'd5249,32'd-164,32'd-3552,32'd2687,32'd8447,32'd-5312,32'd422,32'd3210,32'd66,32'd6196,32'd-5874,32'd2478,32'd718,32'd3750,32'd833,32'd1325,32'd-2285,32'd-1298,32'd1722,32'd-1585,32'd-42,32'd-418,32'd777,32'd-995,32'd3562,32'd5908,32'd2109,32'd-882,32'd1676,32'd-1661,32'd-778,32'd5903,32'd3464,32'd-875,32'd1605,32'd1285,32'd4020,32'd3762,32'd-385,32'd-935,32'd5019,32'd2602,32'd-1090,32'd-1021,32'd297,32'd-2384,32'd2312,32'd-1245,32'd6396,32'd-3503,32'd3107,32'd-190,32'd1981,32'd1885,32'd-832,32'd1749,32'd1257,32'd-3190,32'd-6499,32'd4633,32'd1876,32'd-229,32'd142,32'd8466,32'd-2770,32'd3012,32'd1375,32'd-2010,32'd-549,32'd-1965,32'd5166,32'd2604,32'd3222,32'd4072,32'd-2392,32'd-1826,32'd50,32'd-2203,32'd-3081,32'd5249,32'd22226,32'd5556,32'd1284,32'd-1746,32'd1431,32'd2382,32'd-7675,32'd-8666,32'd5214,32'd-1248,32'd-11318,32'd-9062,32'd4724,32'd3200,32'd-7836,32'd15537,32'd-11865,32'd-5478,32'd4738,32'd-7329,32'd-5522,32'd5263,32'd-9487,32'd2330,32'd-12861,32'd-374,32'd2102,32'd4245,32'd3220,32'd1607,32'd-7065,32'd-16474,32'd-2941,32'd9692,32'd11,32'd-3347,32'd7983,32'd1732,32'd-3784,32'd-1051,32'd1297,32'd-2604,32'd-3515,32'd3391,32'd-1973,32'd-15302,32'd-8378,32'd-2105,32'd6596,32'd6220,32'd15576,32'd2475,32'd-4357,32'd-1325,32'd-3288,32'd1268,32'd-7397,32'd-1754,32'd-1472,32'd2266,32'd-8457,32'd4267,32'd1472,32'd9252,32'd1516,32'd1409,32'd-553,32'd-4443,32'd-5703,32'd739,32'd-10156,32'd1785,32'd94,32'd1374,32'd-690,32'd-898,32'd-2218,32'd-10400,32'd978,32'd-8500,32'd-1187,32'd1237,32'd1070,32'd-5078,32'd-4675,32'd-13300,32'd7060,32'd4013,32'd1518,32'd2719,32'd894,32'd9194,32'd100,32'd-3120,32'd-2329,32'd5366,32'd-3132,32'd-7001,32'd-2293,32'd-605,32'd-4895,32'd3251,32'd-1917,32'd6298,32'd228,32'd-4052,32'd870,32'd-4765,32'd-8183,32'd1215,32'd364,32'd2303,32'd-2277,32'd-75,32'd-1030,32'd-3066,32'd4345,32'd-294,32'd-6401,32'd-304,32'd2834,32'd-31,32'd-6416,32'd-2117,32'd-3637,32'd3088,32'd4890,32'd-9697,32'd586,32'd1417,32'd-3977,32'd3666,32'd-1117,32'd-309,32'd-793,32'd1115,32'd-7539,32'd888,32'd-1911,32'd-4365,32'd-6132,32'd515,32'd-1495,32'd-430,32'd2724,32'd-3422,32'd1096,32'd-2556,32'd2008,32'd5507,32'd1337,32'd-782,32'd-5327,32'd-3828,32'd-4113,32'd-4008,32'd3022,32'd-7719,32'd-1665,32'd5292,32'd-5698,32'd-2814,32'd593,32'd5439,32'd-5908,32'd3576,32'd-13242,32'd4179,32'd-6132,32'd5737,32'd-6044,32'd-4899,32'd1315,32'd7763,32'd-1192,32'd1078,32'd27,32'd-4416,32'd7861,32'd-579,32'd-847,32'd3249,32'd891,32'd-2332,32'd-4953,32'd-3508,32'd6127,32'd-3166,32'd-1361,32'd129,32'd672,32'd5971,32'd4274,32'd6464,32'd-3962,32'd519,32'd-1973,32'd2169,32'd1781,32'd-567,32'd-3020,32'd-11279,32'd-6552,32'd3303,32'd-3452,32'd247,32'd1834,32'd-8803,32'd-13613,32'd4926,32'd1600,32'd-3669,32'd-6113,32'd-80,32'd-6196,32'd2248,32'd-842,32'd484,32'd-4118,32'd-5087,32'd-444,32'd-6093,32'd-2341,32'd-6567,32'd-276,32'd-2138,32'd6889,32'd-5424,32'd8012,32'd4926,32'd-8168,32'd208,32'd-2314,32'd3068,32'd8227,32'd1760,32'd2575,32'd4440,32'd634,32'd-3950,32'd475,32'd-133,32'd245,32'd4145,32'd-9858,32'd6806,32'd-3410,32'd-4670,32'd620,32'd5307,32'd-1348,32'd-2932,32'd-6074,32'd8315,32'd3569,32'd115,32'd-4050,32'd17,32'd8076,32'd260,32'd-10585,32'd-3166,32'd6669,32'd-13056,32'd-269,32'd2232,32'd10468,32'd6459,32'd-3510};
    Wx[2]='{32'd-2290,32'd5834,32'd-2166,32'd-440,32'd833,32'd-1110,32'd3168,32'd5678,32'd-485,32'd-415,32'd3071,32'd-838,32'd6782,32'd-2108,32'd4978,32'd3525,32'd-8276,32'd4807,32'd2937,32'd2111,32'd1343,32'd1026,32'd-4538,32'd3178,32'd-138,32'd1131,32'd-487,32'd1563,32'd2829,32'd8876,32'd-2069,32'd8051,32'd1767,32'd1799,32'd-3918,32'd-1702,32'd4411,32'd3222,32'd869,32'd2025,32'd3349,32'd-2124,32'd-185,32'd2006,32'd-252,32'd-538,32'd-2990,32'd2185,32'd3715,32'd665,32'd3513,32'd10585,32'd1539,32'd1430,32'd2192,32'd-251,32'd4829,32'd-1114,32'd3605,32'd2968,32'd4682,32'd1182,32'd557,32'd308,32'd-292,32'd-3881,32'd-632,32'd7373,32'd906,32'd221,32'd-244,32'd3442,32'd515,32'd6728,32'd1580,32'd-930,32'd-3356,32'd1623,32'd-1708,32'd-519,32'd2061,32'd2727,32'd3024,32'd-2180,32'd-1903,32'd5922,32'd-3,32'd2474,32'd-1386,32'd799,32'd3984,32'd3173,32'd-4641,32'd-345,32'd3649,32'd2763,32'd3300,32'd5034,32'd3615,32'd3964,32'd-555,32'd-8715,32'd151,32'd535,32'd-3776,32'd578,32'd10400,32'd-6596,32'd-4194,32'd-1437,32'd6889,32'd-8388,32'd3774,32'd-5229,32'd-3168,32'd-5537,32'd2464,32'd2568,32'd-1842,32'd5932,32'd479,32'd-144,32'd2440,32'd-6772,32'd-4191,32'd5112,32'd-5405,32'd-1348,32'd-6533,32'd12021,32'd-235,32'd13652,32'd3164,32'd-7055,32'd580,32'd-5629,32'd-1439,32'd7929,32'd-2988,32'd-9238,32'd4506,32'd718,32'd-15126,32'd-3625,32'd-7993,32'd-2722,32'd9311,32'd-1068,32'd1965,32'd-5830,32'd1086,32'd-7885,32'd-6147,32'd-10537,32'd-999,32'd-997,32'd-8012,32'd-1826,32'd-7270,32'd1997,32'd-5468,32'd828,32'd-18730,32'd2934,32'd2498,32'd341,32'd8408,32'd-12744,32'd-1989,32'd64,32'd-834,32'd-1106,32'd-242,32'd-12509,32'd1473,32'd-6748,32'd-1668,32'd12675,32'd6235,32'd1617,32'd735,32'd-131,32'd-9379,32'd-11376,32'd7543,32'd1028,32'd-4384,32'd-4885,32'd-3337,32'd-6665,32'd3220,32'd10820,32'd1198,32'd3732,32'd-4594,32'd6250,32'd1644,32'd-1787,32'd-9589,32'd-5815,32'd-3078,32'd-17617,32'd-2973,32'd-838,32'd4348,32'd-79,32'd-8383,32'd1903,32'd3754,32'd874,32'd-5268,32'd2390,32'd2006,32'd-419,32'd-2656,32'd-7290,32'd-6718,32'd-533,32'd-384,32'd4052,32'd-1183,32'd-2144,32'd702,32'd5053,32'd-1557,32'd-6967,32'd1210,32'd600,32'd-8071,32'd1557,32'd2036,32'd7934,32'd-12822,32'd-1376,32'd-1237,32'd-4863,32'd-3986,32'd913,32'd-5961,32'd-3244,32'd152,32'd-12929,32'd1765,32'd-996,32'd-3713,32'd2239,32'd1749,32'd-2374,32'd-3466,32'd-1414,32'd7622,32'd1099,32'd-1239,32'd-5830,32'd-307,32'd-4350,32'd-6176,32'd838,32'd-10175,32'd-3862,32'd-2832,32'd-5146,32'd-1585,32'd3793,32'd1702,32'd-8242,32'd-1738,32'd-6992,32'd-527,32'd-2473,32'd44,32'd-3898,32'd-2780,32'd-9721,32'd88,32'd-350,32'd-227,32'd-7856,32'd1391,32'd1082,32'd2507,32'd-9360,32'd-1857,32'd4621,32'd-3215,32'd-9311,32'd-1309,32'd761,32'd-6108,32'd120,32'd-2604,32'd-2064,32'd-4020,32'd-4794,32'd-17773,32'd-3459,32'd-797,32'd-3776,32'd1861,32'd-3403,32'd1766,32'd-4902,32'd9990,32'd-878,32'd2479,32'd-151,32'd-5449,32'd-1232,32'd464,32'd6171,32'd675,32'd-5903,32'd6801,32'd-4367,32'd7290,32'd-3701,32'd-8261,32'd-5825,32'd6083,32'd-2106,32'd1777,32'd-2727,32'd1304,32'd3916,32'd3127,32'd-5400,32'd-6708,32'd5249,32'd-2724,32'd-92,32'd778,32'd12324,32'd-3564,32'd-6103,32'd-10361,32'd-4892,32'd-3940,32'd-1065,32'd2061,32'd-4770,32'd2156,32'd-9023,32'd2624,32'd2204,32'd-2396,32'd-1202,32'd-753,32'd-7001,32'd7915,32'd-503,32'd-1875,32'd4790,32'd3154,32'd1801,32'd-1816,32'd-2880,32'd-357,32'd-9736,32'd-2359,32'd2052,32'd-533,32'd-1429,32'd-1816,32'd7246,32'd-2995,32'd-4455,32'd1160,32'd-6845,32'd9760,32'd-864,32'd-460,32'd6435,32'd-1812,32'd-4079,32'd4460,32'd617,32'd-3920,32'd-2885,32'd-6206,32'd-5073,32'd1684,32'd-248,32'd-6362,32'd-1962,32'd5004,32'd-1857,32'd7065,32'd-6186,32'd-661,32'd2082,32'd-2907,32'd-3293,32'd-3813,32'd15185,32'd845,32'd-2905,32'd-2841,32'd4204,32'd-1400,32'd4619};
    Wx[3]='{32'd-1378,32'd-2309,32'd-282,32'd2299,32'd-298,32'd-214,32'd1143,32'd-1861,32'd-3410,32'd-574,32'd2142,32'd3945,32'd-971,32'd-3937,32'd5864,32'd3054,32'd-1604,32'd2622,32'd2875,32'd842,32'd2017,32'd2160,32'd1865,32'd1461,32'd-1249,32'd-507,32'd2336,32'd-164,32'd-841,32'd-3747,32'd-1455,32'd242,32'd1093,32'd26,32'd6474,32'd2692,32'd-655,32'd-2164,32'd1408,32'd1848,32'd3530,32'd3967,32'd-2656,32'd2299,32'd-6035,32'd1715,32'd184,32'd1267,32'd-22,32'd-454,32'd-8232,32'd2966,32'd3361,32'd-1784,32'd-633,32'd2434,32'd-583,32'd4980,32'd-4274,32'd-3503,32'd2331,32'd3771,32'd-2758,32'd944,32'd2758,32'd1129,32'd-3142,32'd5898,32'd-4025,32'd429,32'd-892,32'd-741,32'd2352,32'd-1569,32'd466,32'd6523,32'd2731,32'd3815,32'd-167,32'd255,32'd402,32'd4348,32'd-1184,32'd2971,32'd1939,32'd4001,32'd878,32'd-2250,32'd1079,32'd7675,32'd2631,32'd1065,32'd1727,32'd-3020,32'd3574,32'd-3078,32'd-4484,32'd4213,32'd-106,32'd3627,32'd-977,32'd-11533,32'd917,32'd-199,32'd-3879,32'd919,32'd-8740,32'd-1040,32'd-4504,32'd-2614,32'd3798,32'd5678,32'd5615,32'd16455,32'd265,32'd7768,32'd-10937,32'd-8652,32'd4731,32'd1784,32'd-1571,32'd6074,32'd-1126,32'd5966,32'd-429,32'd-2094,32'd2299,32'd-6909,32'd-11572,32'd-2819,32'd207,32'd8466,32'd-6728,32'd2392,32'd3859,32'd6884,32'd-3774,32'd5258,32'd9414,32'd-9355,32'd1990,32'd-12490,32'd-4589,32'd7426,32'd7246,32'd-969,32'd16123,32'd-567,32'd-1239,32'd2091,32'd-2093,32'd-8925,32'd5874,32'd-3840,32'd1618,32'd1334,32'd7709,32'd-3981,32'd3562,32'd1700,32'd-1507,32'd15136,32'd-4377,32'd-1738,32'd1712,32'd-3020,32'd4909,32'd5429,32'd4680,32'd-1998,32'd2575,32'd-12119,32'd-3278,32'd2478,32'd614,32'd-10009,32'd14658,32'd-9428,32'd-12324,32'd6982,32'd-4682,32'd-344,32'd-5795,32'd-2330,32'd819,32'd9960,32'd-5073,32'd-1693,32'd401,32'd4995,32'd-2392,32'd-3208,32'd-10673,32'd-1693,32'd244,32'd693,32'd-4008,32'd4121,32'd-4582,32'd3312,32'd687,32'd8798,32'd1505,32'd3642,32'd4589,32'd1597,32'd6000,32'd181,32'd-4316,32'd467,32'd-1317,32'd-2719,32'd-775,32'd2868,32'd4702,32'd-1191,32'd-9990,32'd7128,32'd617,32'd2866,32'd2081,32'd-1832,32'd-1967,32'd2434,32'd2714,32'd4262,32'd-1191,32'd2905,32'd-70,32'd2261,32'd5830,32'd-4865,32'd10878,32'd403,32'd1455,32'd-3217,32'd-3886,32'd249,32'd-5600,32'd-2423,32'd7465,32'd2846,32'd2054,32'd12011,32'd-7626,32'd-6494,32'd-6635,32'd-885,32'd-1210,32'd2330,32'd1209,32'd-4750,32'd6240,32'd1488,32'd3095,32'd2639,32'd-5209,32'd3142,32'd5112,32'd792,32'd-4550,32'd4970,32'd-3093,32'd634,32'd2978,32'd-600,32'd-4750,32'd-3237,32'd-1166,32'd-2897,32'd1100,32'd2778,32'd-850,32'd391,32'd1134,32'd-1589,32'd-2644,32'd-3828,32'd-7973,32'd-2980,32'd1318,32'd-8920,32'd-75,32'd-6538,32'd3288,32'd-1279,32'd7,32'd6254,32'd-1126,32'd-411,32'd-2946,32'd3977,32'd2563,32'd-1843,32'd-7255,32'd6333,32'd-8564,32'd502,32'd4045,32'd-2570,32'd989,32'd11152,32'd-2812,32'd199,32'd4062,32'd-6044,32'd10908,32'd-512,32'd-1544,32'd215,32'd1069,32'd69,32'd2286,32'd555,32'd4768,32'd-10849,32'd-389,32'd3298,32'd1457,32'd3679,32'd881,32'd-722,32'd4484,32'd7626,32'd2153,32'd8413,32'd3662,32'd2683,32'd4055,32'd4438,32'd1677,32'd-654,32'd13173,32'd2078,32'd3303,32'd-5566,32'd-2412,32'd-1442,32'd903,32'd3842,32'd6289,32'd2648,32'd-72,32'd5888,32'd-3652,32'd-4721,32'd3127,32'd-3146,32'd-6640,32'd-219,32'd1203,32'd-3115,32'd2379,32'd-8500,32'd8056,32'd1806,32'd-2761,32'd-1246,32'd7773,32'd414,32'd561,32'd-2094,32'd-3776,32'd2238,32'd5400,32'd-3522,32'd-7993,32'd-428,32'd-6718,32'd1594,32'd-5874,32'd604,32'd4692,32'd1888,32'd4423,32'd4973,32'd8798,32'd-487,32'd-5922,32'd-1259,32'd-351,32'd-1043,32'd6914,32'd-4313,32'd5400,32'd-1370,32'd4870,32'd3085,32'd-1842,32'd4897,32'd-4536,32'd2425,32'd-60,32'd919,32'd-3164,32'd693,32'd-6621,32'd3945,32'd7241,32'd-10283};
    Wx[4]='{32'd-2120,32'd1262,32'd-1751,32'd-261,32'd-1295,32'd485,32'd2841,32'd-2780,32'd-6284,32'd2010,32'd3139,32'd-184,32'd-10283,32'd802,32'd-1137,32'd-526,32'd-6420,32'd-871,32'd-979,32'd-1685,32'd283,32'd-1663,32'd358,32'd-1470,32'd-5834,32'd-240,32'd2242,32'd-3981,32'd-583,32'd-2949,32'd-144,32'd-2261,32'd-442,32'd-3454,32'd-9301,32'd956,32'd-3791,32'd-1911,32'd-1442,32'd4643,32'd57,32'd1027,32'd-7158,32'd2902,32'd-2575,32'd-4560,32'd-4985,32'd2219,32'd-4907,32'd444,32'd4348,32'd-451,32'd-1375,32'd-1580,32'd-892,32'd-7788,32'd859,32'd-1555,32'd-220,32'd-3784,32'd-2548,32'd-2465,32'd-758,32'd-5336,32'd-758,32'd990,32'd-2415,32'd3879,32'd-471,32'd-889,32'd-3083,32'd3105,32'd-4816,32'd2653,32'd-4172,32'd-8715,32'd337,32'd1502,32'd-3498,32'd-6289,32'd-2471,32'd1137,32'd-900,32'd-3461,32'd-28,32'd-8354,32'd460,32'd-508,32'd-3251,32'd-1368,32'd648,32'd8701,32'd515,32'd2626,32'd-2976,32'd-2495,32'd-3339,32'd1925,32'd-2067,32'd-385,32'd1574,32'd5048,32'd385,32'd3757,32'd-4018,32'd-267,32'd-7280,32'd-5039,32'd4467,32'd4294,32'd-3935,32'd-2946,32'd-858,32'd4577,32'd-21406,32'd3498,32'd-5439,32'd1093,32'd1303,32'd-1646,32'd2800,32'd5532,32'd3469,32'd-613,32'd-5239,32'd-2152,32'd-578,32'd823,32'd1278,32'd3103,32'd2391,32'd19951,32'd12841,32'd-4777,32'd-3305,32'd6528,32'd-5473,32'd2297,32'd-3918,32'd-7158,32'd-3688,32'd-8398,32'd-3833,32'd-3344,32'd-9331,32'd2949,32'd-5014,32'd6850,32'd-9658,32'd-4838,32'd-6196,32'd-10839,32'd3894,32'd15087,32'd-1883,32'd-9208,32'd-1602,32'd-4160,32'd5581,32'd1441,32'd-2257,32'd9536,32'd4421,32'd12255,32'd-2644,32'd2954,32'd4982,32'd-17255,32'd369,32'd-3820,32'd-6362,32'd-3591,32'd498,32'd2836,32'd-804,32'd-9252,32'd454,32'd-4160,32'd11484,32'd-5229,32'd-3164,32'd1368,32'd-1318,32'd-5878,32'd-7807,32'd-409,32'd159,32'd-975,32'd-4018,32'd-2570,32'd-14941,32'd-4301,32'd-5732,32'd-3225,32'd-1145,32'd-8183,32'd-1695,32'd2641,32'd2161,32'd4665,32'd-4921,32'd8496,32'd1102,32'd-2985,32'd2017,32'd1074,32'd-4084,32'd-8027,32'd712,32'd396,32'd-2939,32'd1063,32'd-6479,32'd-6391,32'd-3332,32'd1160,32'd13486,32'd4567,32'd-764,32'd-1018,32'd4960,32'd-1652,32'd-4833,32'd2663,32'd3911,32'd-246,32'd-24,32'd2133,32'd748,32'd-398,32'd484,32'd-3125,32'd1468,32'd-9257,32'd849,32'd-3305,32'd-2207,32'd2856,32'd-26,32'd-279,32'd-3425,32'd5810,32'd4621,32'd9951,32'd862,32'd109,32'd-9965,32'd-4572,32'd-3710,32'd-403,32'd-1494,32'd-5634,32'd-4584,32'd2724,32'd-2291,32'd1324,32'd-2004,32'd4899,32'd-3334,32'd8276,32'd-1549,32'd-1044,32'd-223,32'd-11367,32'd3020,32'd1086,32'd-2072,32'd2736,32'd995,32'd1845,32'd940,32'd792,32'd-5048,32'd-7368,32'd-4809,32'd-3005,32'd-8027,32'd-256,32'd1879,32'd-47,32'd-2122,32'd4931,32'd23,32'd-164,32'd-1016,32'd278,32'd-2260,32'd-4858,32'd1860,32'd3347,32'd-2722,32'd2719,32'd-4531,32'd-958,32'd-6513,32'd-858,32'd-9047,32'd-3210,32'd-8051,32'd8857,32'd-3657,32'd4035,32'd1549,32'd1693,32'd-1374,32'd-922,32'd-3452,32'd-13193,32'd-4104,32'd-1779,32'd-126,32'd-5195,32'd-13984,32'd373,32'd-411,32'd3422,32'd6499,32'd207,32'd1627,32'd-4685,32'd1172,32'd-5283,32'd-2731,32'd3786,32'd-1486,32'd3366,32'd1727,32'd647,32'd1159,32'd640,32'd2990,32'd-6645,32'd3317,32'd-804,32'd2082,32'd-6035,32'd-6850,32'd2349,32'd4848,32'd518,32'd2734,32'd6279,32'd1583,32'd6083,32'd191,32'd-139,32'd-10556,32'd-3989,32'd3637,32'd431,32'd9545,32'd-2221,32'd-6728,32'd-8442,32'd5405,32'd-7568,32'd-3491,32'd-9067,32'd3437,32'd-1970,32'd-1343,32'd-450,32'd-6962,32'd-3940,32'd4262,32'd2978,32'd-8164,32'd10566,32'd-1456,32'd-11884,32'd-3278,32'd-1367,32'd-3295,32'd-1588,32'd-3208,32'd-10410,32'd-708,32'd-1604,32'd-1754,32'd-2836,32'd-2695,32'd9638,32'd2010,32'd-696,32'd-6469,32'd-5322,32'd1120,32'd-4228,32'd-2744,32'd-431,32'd3315,32'd-9755,32'd-3637,32'd6376,32'd-2648,32'd-324,32'd-8842,32'd-2800,32'd-4729,32'd6552};
    Wx[5]='{32'd155,32'd2254,32'd368,32'd-125,32'd-80,32'd-1270,32'd3820,32'd2248,32'd3728,32'd-449,32'd4257,32'd1976,32'd1739,32'd-1855,32'd3935,32'd-3686,32'd-7739,32'd9492,32'd2644,32'd2005,32'd-153,32'd1569,32'd573,32'd-713,32'd2048,32'd-1510,32'd-3676,32'd2230,32'd2175,32'd135,32'd-793,32'd943,32'd2517,32'd0,32'd742,32'd-1204,32'd-2374,32'd291,32'd-367,32'd-786,32'd-354,32'd2200,32'd-1906,32'd339,32'd214,32'd-183,32'd-3432,32'd-275,32'd2961,32'd-3801,32'd-5019,32'd802,32'd-957,32'd4282,32'd1129,32'd3461,32'd3337,32'd-991,32'd1687,32'd2536,32'd2854,32'd2073,32'd6850,32'd-3120,32'd-190,32'd-2651,32'd-123,32'd-2927,32'd903,32'd-561,32'd-6767,32'd4199,32'd-3103,32'd1376,32'd-1268,32'd-590,32'd6088,32'd877,32'd-5336,32'd2133,32'd-30,32'd-6660,32'd2026,32'd3212,32'd-1882,32'd3347,32'd-30,32'd-1730,32'd44,32'd-1605,32'd-750,32'd-4113,32'd5224,32'd-2946,32'd-3823,32'd-1096,32'd4470,32'd4968,32'd1403,32'd609,32'd1684,32'd14921,32'd1478,32'd-6494,32'd3996,32'd4631,32'd-11328,32'd-12714,32'd3291,32'd-3388,32'd11250,32'd1951,32'd-3222,32'd3913,32'd6782,32'd6518,32'd6127,32'd-5834,32'd-3022,32'd-2583,32'd2207,32'd5795,32'd5488,32'd9628,32'd2067,32'd4025,32'd2482,32'd2944,32'd5390,32'd646,32'd-3952,32'd17382,32'd5986,32'd1138,32'd3469,32'd4233,32'd6171,32'd2004,32'd-8261,32'd-6201,32'd-1975,32'd-3610,32'd-17304,32'd8486,32'd3442,32'd-7441,32'd14873,32'd2663,32'd3530,32'd-12021,32'd11552,32'd-13437,32'd650,32'd-10175,32'd4614,32'd-1190,32'd8330,32'd2415,32'd-4377,32'd101,32'd-1479,32'd-3718,32'd4477,32'd-5668,32'd9350,32'd922,32'd2690,32'd-8608,32'd-570,32'd-5112,32'd-139,32'd-12343,32'd-3547,32'd-10312,32'd-1286,32'd17128,32'd-7539,32'd-10126,32'd-2102,32'd-6328,32'd3640,32'd429,32'd-7602,32'd-1029,32'd177,32'd-10468,32'd6030,32'd5805,32'd988,32'd-5102,32'd153,32'd-4628,32'd-4345,32'd-1459,32'd9189,32'd-2124,32'd-4084,32'd8125,32'd9443,32'd6875,32'd-3449,32'd3986,32'd-339,32'd2340,32'd-1699,32'd-3437,32'd-7099,32'd-5380,32'd-3210,32'd5224,32'd2136,32'd2059,32'd629,32'd-10615,32'd-5029,32'd-7436,32'd-8750,32'd-2783,32'd-1756,32'd824,32'd-827,32'd1,32'd3708,32'd-7221,32'd-1063,32'd-2946,32'd-4057,32'd-244,32'd-1145,32'd-2221,32'd-2294,32'd-6010,32'd-6938,32'd-8256,32'd-1331,32'd-3576,32'd-8520,32'd-8715,32'd2116,32'd-6386,32'd1397,32'd-10312,32'd1397,32'd-7753,32'd4919,32'd-5625,32'd5917,32'd-2154,32'd1916,32'd-1881,32'd-8110,32'd6269,32'd-2778,32'd-2819,32'd3222,32'd-3596,32'd-1741,32'd-876,32'd5429,32'd1823,32'd2617,32'd-6240,32'd-5083,32'd2358,32'd-4616,32'd-6699,32'd-1828,32'd-1079,32'd4038,32'd1080,32'd5151,32'd-1613,32'd-1571,32'd2849,32'd-1506,32'd-951,32'd4707,32'd-8369,32'd-2119,32'd60,32'd-2646,32'd-4350,32'd-127,32'd-1131,32'd-4140,32'd-4819,32'd-79,32'd1057,32'd-1354,32'd-1596,32'd-1992,32'd-783,32'd-4436,32'd-2310,32'd-3066,32'd-7612,32'd-4360,32'd-3569,32'd6884,32'd-2430,32'd-7050,32'd5473,32'd4965,32'd1818,32'd-2159,32'd-5043,32'd4384,32'd-5698,32'd-4074,32'd5185,32'd-4216,32'd6743,32'd-3034,32'd-10947,32'd-4902,32'd-3205,32'd-4929,32'd-2175,32'd-674,32'd3637,32'd-3132,32'd-3879,32'd1383,32'd-3005,32'd-3212,32'd-1976,32'd-1947,32'd-1768,32'd-1472,32'd-1082,32'd-913,32'd-10185,32'd-6650,32'd-1499,32'd1417,32'd-1768,32'd-5566,32'd-3251,32'd-3063,32'd-4179,32'd4904,32'd-3461,32'd-1470,32'd-4133,32'd6679,32'd-2462,32'd7646,32'd-4023,32'd-939,32'd-5400,32'd-1183,32'd1331,32'd-345,32'd-5947,32'd8022,32'd5341,32'd-3610,32'd-3037,32'd3442,32'd1485,32'd619,32'd1318,32'd-8779,32'd390,32'd-4104,32'd-4016,32'd1898,32'd-10107,32'd1475,32'd5449,32'd-3122,32'd5556,32'd-236,32'd-2824,32'd5102,32'd-5371,32'd-2281,32'd-6088,32'd3234,32'd2318,32'd-1575,32'd1502,32'd2695,32'd7539,32'd-104,32'd-5019,32'd3718,32'd913,32'd-655,32'd1527,32'd-3334,32'd-6855,32'd-5825,32'd17861,32'd-4079,32'd-8432,32'd2614,32'd2714,32'd3271,32'd-3728};
    Wx[6]='{32'd-1413,32'd2678,32'd3400,32'd-1433,32'd1183,32'd2570,32'd4470,32'd4216,32'd-1572,32'd-1800,32'd-1971,32'd1004,32'd-307,32'd2934,32'd1525,32'd7988,32'd1459,32'd2305,32'd3645,32'd-3310,32'd-3156,32'd-2663,32'd2312,32'd-330,32'd3869,32'd11,32'd1812,32'd-1346,32'd4763,32'd1206,32'd506,32'd-1147,32'd5957,32'd1628,32'd-3999,32'd-284,32'd1291,32'd-2031,32'd167,32'd5502,32'd548,32'd-466,32'd6455,32'd919,32'd6884,32'd-2177,32'd3703,32'd1334,32'd1989,32'd1062,32'd2185,32'd1505,32'd2829,32'd535,32'd-875,32'd3935,32'd-640,32'd-5410,32'd3869,32'd-1784,32'd-2369,32'd-3908,32'd704,32'd-1066,32'd4707,32'd-2800,32'd201,32'd5502,32'd1161,32'd-2142,32'd1047,32'd2500,32'd4501,32'd311,32'd-4489,32'd-1826,32'd4804,32'd1489,32'd698,32'd6381,32'd1369,32'd1243,32'd-4929,32'd2329,32'd2631,32'd8491,32'd-161,32'd4025,32'd-823,32'd-4204,32'd3044,32'd-1796,32'd-1244,32'd2091,32'd-4050,32'd-884,32'd2401,32'd140,32'd294,32'd-4421,32'd-1602,32'd-3527,32'd-3413,32'd9282,32'd-1024,32'd-520,32'd7832,32'd5234,32'd9960,32'd-990,32'd721,32'd-4672,32'd-7797,32'd14755,32'd-5166,32'd-5375,32'd-2281,32'd-2685,32'd-7749,32'd-2805,32'd-3356,32'd6044,32'd-631,32'd2229,32'd3525,32'd6508,32'd1273,32'd3789,32'd8002,32'd-1594,32'd-3449,32'd14482,32'd9370,32'd1241,32'd2172,32'd7700,32'd-914,32'd340,32'd-10048,32'd-9282,32'd677,32'd-7011,32'd-8764,32'd13251,32'd1677,32'd4384,32'd1389,32'd-9663,32'd-4755,32'd3593,32'd-6259,32'd-5209,32'd2187,32'd6875,32'd-561,32'd8041,32'd-718,32'd3598,32'd11904,32'd128,32'd3342,32'd564,32'd10957,32'd1477,32'd15351,32'd-164,32'd2333,32'd-349,32'd-1729,32'd-5219,32'd-8442,32'd5717,32'd-4865,32'd3833,32'd3012,32'd10888,32'd724,32'd-19013,32'd-5415,32'd-2880,32'd1263,32'd7192,32'd9970,32'd-2236,32'd-916,32'd-2944,32'd-3137,32'd1966,32'd3913,32'd-3920,32'd-1317,32'd4543,32'd63,32'd568,32'd1469,32'd7187,32'd6562,32'd2142,32'd-4477,32'd1036,32'd1005,32'd2425,32'd8637,32'd430,32'd4677,32'd-795,32'd-4733,32'd1865,32'd570,32'd-846,32'd7890,32'd1085,32'd-251,32'd984,32'd361,32'd-2570,32'd10839,32'd-4382,32'd3066,32'd-1813,32'd-2407,32'd2011,32'd343,32'd-40,32'd5473,32'd-458,32'd708,32'd3728,32'd-14208,32'd-9433,32'd-2186,32'd9726,32'd2766,32'd3364,32'd2005,32'd2108,32'd-892,32'd-189,32'd-466,32'd-8173,32'd-2668,32'd8530,32'd-5317,32'd5996,32'd10546,32'd1523,32'd-1689,32'd-2353,32'd-3232,32'd1480,32'd-787,32'd4279,32'd-157,32'd-1291,32'd5312,32'd4045,32'd620,32'd1916,32'd-1477,32'd-3085,32'd1141,32'd9331,32'd-87,32'd2514,32'd-2641,32'd-121,32'd-446,32'd-2322,32'd1351,32'd-2333,32'd-1676,32'd-4589,32'd451,32'd5097,32'd-371,32'd8974,32'd659,32'd429,32'd-2993,32'd6928,32'd6508,32'd6557,32'd-2551,32'd1030,32'd-897,32'd6328,32'd3964,32'd-3046,32'd1945,32'd-997,32'd-2080,32'd2221,32'd-1040,32'd6279,32'd-7138,32'd320,32'd-1374,32'd8164,32'd-2695,32'd-3740,32'd-2580,32'd211,32'd5263,32'd172,32'd5317,32'd-184,32'd-15068,32'd-11113,32'd-6313,32'd1472,32'd3310,32'd-2766,32'd-3803,32'd-4697,32'd3300,32'd3432,32'd-539,32'd1881,32'd-2958,32'd-1442,32'd-1644,32'd-432,32'd2607,32'd-282,32'd6171,32'd676,32'd1220,32'd2308,32'd-11103,32'd-1807,32'd-6284,32'd-566,32'd4914,32'd510,32'd4494,32'd-2204,32'd1854,32'd2343,32'd1420,32'd-989,32'd1188,32'd-4133,32'd4868,32'd4313,32'd-1330,32'd71,32'd-461,32'd-6015,32'd2120,32'd-3002,32'd4028,32'd-4125,32'd-1216,32'd-444,32'd12470,32'd6826,32'd-5502,32'd-838,32'd3476,32'd-6821,32'd-5351,32'd-686,32'd-3405,32'd-113,32'd5317,32'd-2846,32'd307,32'd5961,32'd-1562,32'd-7446,32'd-736,32'd-9531,32'd-5551,32'd10078,32'd3173,32'd-217,32'd-1606,32'd-3884,32'd-5258,32'd6308,32'd8793,32'd7939,32'd1733,32'd8837,32'd-1541,32'd3481,32'd2485,32'd-2641,32'd-3957,32'd-6406,32'd-2553,32'd8339,32'd-1165,32'd14755,32'd-10478,32'd-2651,32'd6035,32'd6406,32'd5961,32'd-5327};
    Wx[7]='{32'd-2200,32'd5971,32'd1126,32'd56,32'd462,32'd266,32'd6035,32'd4860,32'd3225,32'd2675,32'd-1798,32'd-4223,32'd3271,32'd2678,32'd507,32'd-2067,32'd1276,32'd1165,32'd-3298,32'd8,32'd-1811,32'd2648,32'd110,32'd1350,32'd-1173,32'd-5214,32'd1523,32'd-1113,32'd6269,32'd-145,32'd1372,32'd7841,32'd1260,32'd-945,32'd-2944,32'd-1324,32'd-3156,32'd2739,32'd2403,32'd1420,32'd3620,32'd6406,32'd-2980,32'd2656,32'd1862,32'd-201,32'd-10546,32'd1702,32'd-4328,32'd-2573,32'd5556,32'd503,32'd-3867,32'd1372,32'd-1170,32'd2312,32'd-1494,32'd-6777,32'd3808,32'd-431,32'd853,32'd720,32'd3520,32'd2305,32'd2355,32'd-1209,32'd1800,32'd358,32'd-2932,32'd-4587,32'd-3105,32'd311,32'd-3681,32'd81,32'd-1606,32'd4816,32'd5844,32'd193,32'd-3522,32'd614,32'd2387,32'd-2812,32'd667,32'd-3950,32'd-1231,32'd902,32'd-2081,32'd21,32'd379,32'd-282,32'd-363,32'd3208,32'd4719,32'd-1402,32'd6821,32'd490,32'd5136,32'd10634,32'd-3808,32'd-242,32'd-1693,32'd5341,32'd988,32'd-1838,32'd-1341,32'd0,32'd-6357,32'd96,32'd-5488,32'd-4572,32'd1320,32'd3000,32'd5839,32'd7680,32'd-12519,32'd15136,32'd9687,32'd382,32'd-303,32'd-1611,32'd4179,32'd-5073,32'd1051,32'd-8447,32'd1407,32'd-962,32'd2829,32'd-2792,32'd20488,32'd-2376,32'd-562,32'd-5351,32'd789,32'd-292,32'd5097,32'd-4775,32'd2770,32'd4228,32'd-4797,32'd-874,32'd4680,32'd2883,32'd-6884,32'd-8759,32'd-7197,32'd4094,32'd2094,32'd-8583,32'd20,32'd-4951,32'd-13134,32'd2988,32'd-1385,32'd565,32'd-4787,32'd6333,32'd-1676,32'd2119,32'd-16787,32'd6225,32'd6523,32'd10058,32'd-6899,32'd2331,32'd-7617,32'd-2052,32'd196,32'd-797,32'd-2548,32'd-1061,32'd7045,32'd12910,32'd1459,32'd1215,32'd-1016,32'd4287,32'd9536,32'd-7329,32'd-883,32'd-1243,32'd6850,32'd6035,32'd-9008,32'd14169,32'd-1843,32'd-1240,32'd4555,32'd-2768,32'd-2910,32'd-309,32'd-8447,32'd-7460,32'd3676,32'd-962,32'd489,32'd-5004,32'd2866,32'd18974,32'd2348,32'd5346,32'd3552,32'd-12304,32'd1318,32'd6542,32'd1761,32'd2971,32'd-28,32'd-9541,32'd387,32'd-428,32'd2646,32'd1799,32'd1717,32'd7832,32'd-12763,32'd9072,32'd-1934,32'd1134,32'd1074,32'd-1953,32'd-1878,32'd1253,32'd-1328,32'd2369,32'd-4714,32'd-1867,32'd-2846,32'd2126,32'd-1813,32'd2558,32'd2670,32'd4023,32'd-4887,32'd-620,32'd-2072,32'd-4536,32'd-836,32'd-2211,32'd1510,32'd1944,32'd-1334,32'd-3225,32'd9223,32'd-4880,32'd-508,32'd4692,32'd5507,32'd258,32'd4865,32'd6069,32'd3276,32'd12314,32'd-550,32'd9536,32'd823,32'd-1938,32'd4157,32'd-5761,32'd3867,32'd4006,32'd2113,32'd-2259,32'd1890,32'd-1081,32'd2320,32'd-617,32'd3691,32'd-4365,32'd1197,32'd-5249,32'd1645,32'd1245,32'd5180,32'd1331,32'd477,32'd1306,32'd-426,32'd-4924,32'd2583,32'd-195,32'd-2480,32'd-1481,32'd9296,32'd5532,32'd-5366,32'd1102,32'd2583,32'd-235,32'd2973,32'd4274,32'd3205,32'd-2004,32'd-5488,32'd4626,32'd-866,32'd-2941,32'd1530,32'd5400,32'd-4062,32'd334,32'd-1662,32'd6650,32'd2067,32'd8828,32'd-1290,32'd-7290,32'd-8354,32'd-11132,32'd2824,32'd80,32'd2690,32'd6030,32'd-554,32'd3005,32'd-5424,32'd7641,32'd-2275,32'd9130,32'd2583,32'd-2912,32'd-13525,32'd4912,32'd993,32'd2290,32'd-7924,32'd-203,32'd-2773,32'd-243,32'd2009,32'd-7539,32'd-2614,32'd8090,32'd-2227,32'd1110,32'd-237,32'd-5034,32'd-4624,32'd1298,32'd-3063,32'd3051,32'd1639,32'd1574,32'd3176,32'd1746,32'd681,32'd8930,32'd585,32'd-1240,32'd-1739,32'd-1156,32'd385,32'd10195,32'd-123,32'd4541,32'd853,32'd297,32'd-1582,32'd-8432,32'd5273,32'd-2410,32'd-4543,32'd150,32'd621,32'd-175,32'd8217,32'd-2822,32'd8828,32'd-11972,32'd5405,32'd29,32'd-2357,32'd-121,32'd828,32'd3820,32'd-9008,32'd-1634,32'd114,32'd3208,32'd-5903,32'd2091,32'd-1215,32'd5170,32'd9472,32'd248,32'd-11972,32'd6796,32'd5039,32'd4416,32'd4033,32'd-3391,32'd127,32'd3046,32'd-424,32'd-2719,32'd2426,32'd-6357,32'd4453,32'd-47,32'd3151,32'd3654};
    Wx[8]='{32'd512,32'd1589,32'd1065,32'd1262,32'd1115,32'd-743,32'd-2854,32'd-4377,32'd1734,32'd164,32'd-3076,32'd739,32'd-131,32'd-1416,32'd3159,32'd2155,32'd10156,32'd1095,32'd-161,32'd1115,32'd2103,32'd-221,32'd-2951,32'd897,32'd1058,32'd-2152,32'd4836,32'd524,32'd-5581,32'd-1788,32'd2893,32'd-5156,32'd-8178,32'd-4033,32'd-410,32'd432,32'd-201,32'd2573,32'd-1513,32'd-4443,32'd-1478,32'd-3864,32'd-2927,32'd3083,32'd-4699,32'd817,32'd10878,32'd4541,32'd-2993,32'd-1497,32'd6147,32'd-6181,32'd-92,32'd3498,32'd-1768,32'd5229,32'd646,32'd1679,32'd-3486,32'd-2126,32'd-2705,32'd-3479,32'd-1066,32'd593,32'd-760,32'd1652,32'd3618,32'd-3034,32'd520,32'd1223,32'd718,32'd-9750,32'd2132,32'd1885,32'd2479,32'd-2807,32'd-2849,32'd1362,32'd2025,32'd2922,32'd1133,32'd4428,32'd2380,32'd-1512,32'd2961,32'd-4506,32'd1864,32'd837,32'd1246,32'd-281,32'd4931,32'd-6948,32'd-3981,32'd-4704,32'd-7138,32'd-1739,32'd-1966,32'd-2156,32'd368,32'd2476,32'd-1523,32'd-12792,32'd1381,32'd-4416,32'd2072,32'd-1270,32'd1207,32'd-5878,32'd2531,32'd-3015,32'd1927,32'd838,32'd1846,32'd6894,32'd-15771,32'd-11523,32'd-6621,32'd4172,32'd-1489,32'd650,32'd1425,32'd-2802,32'd-2590,32'd-4514,32'd-2186,32'd-5107,32'd122,32'd-1328,32'd-11748,32'd-5947,32'd931,32'd24160,32'd2207,32'd-4252,32'd362,32'd4121,32'd2700,32'd1431,32'd3845,32'd-5004,32'd2340,32'd-4472,32'd-13105,32'd-745,32'd13623,32'd-549,32'd3957,32'd-7485,32'd-1098,32'd5117,32'd-1165,32'd-9838,32'd3774,32'd-924,32'd7260,32'd8520,32'd-9370,32'd1060,32'd1100,32'd2839,32'd1138,32'd-4042,32'd-5048,32'd-4328,32'd-6035,32'd-442,32'd-3137,32'd-7929,32'd-351,32'd1252,32'd-5732,32'd-11796,32'd-6391,32'd-8154,32'd3745,32'd260,32'd-7412,32'd-8955,32'd-9438,32'd-1798,32'd-2084,32'd1887,32'd1396,32'd14228,32'd6240,32'd4499,32'd3686,32'd-2573,32'd-1680,32'd3881,32'd2529,32'd11367,32'd-6225,32'd-492,32'd-12080,32'd8339,32'd4235,32'd5288,32'd-2727,32'd-760,32'd550,32'd2915,32'd2663,32'd-482,32'd249,32'd734,32'd5795,32'd-102,32'd-4353,32'd1549,32'd-3156,32'd2147,32'd-346,32'd-1010,32'd5371,32'd321,32'd751,32'd6401,32'd4899,32'd842,32'd1475,32'd1445,32'd2076,32'd3762,32'd1433,32'd5214,32'd733,32'd1412,32'd-1173,32'd-1205,32'd2507,32'd1112,32'd2055,32'd-2824,32'd-10156,32'd-1228,32'd1542,32'd2558,32'd-6689,32'd-2851,32'd-2271,32'd-1199,32'd-7529,32'd2661,32'd-5629,32'd-5747,32'd-8159,32'd1750,32'd-4887,32'd-4694,32'd-6997,32'd6586,32'd3815,32'd-5239,32'd-4106,32'd-1723,32'd-4228,32'd5571,32'd-795,32'd-4682,32'd1231,32'd-1267,32'd2761,32'd-1323,32'd-2580,32'd2702,32'd5053,32'd-4072,32'd-212,32'd-1888,32'd2028,32'd3820,32'd-743,32'd-4331,32'd2612,32'd136,32'd4440,32'd3183,32'd-2700,32'd1702,32'd2255,32'd-1148,32'd1470,32'd-5366,32'd-3881,32'd99,32'd-108,32'd1850,32'd-8271,32'd1076,32'd-5913,32'd-145,32'd-1967,32'd616,32'd-34,32'd3732,32'd6298,32'd239,32'd3625,32'd-1459,32'd-1300,32'd2143,32'd3034,32'd2966,32'd-1208,32'd2205,32'd4477,32'd227,32'd-5004,32'd-2243,32'd-4331,32'd-2149,32'd-6293,32'd-3085,32'd2873,32'd-1491,32'd-1514,32'd3466,32'd-2003,32'd-849,32'd-2656,32'd1555,32'd-2509,32'd7431,32'd3710,32'd-2763,32'd2253,32'd6958,32'd-2617,32'd-547,32'd1513,32'd-1176,32'd-6572,32'd-983,32'd5205,32'd542,32'd6523,32'd1702,32'd531,32'd-4016,32'd-2705,32'd3562,32'd-3117,32'd-1652,32'd-6655,32'd-10966,32'd-1034,32'd3488,32'd1781,32'd-4335,32'd2148,32'd1340,32'd693,32'd-9291,32'd270,32'd-1230,32'd-3684,32'd2539,32'd3125,32'd-1677,32'd3229,32'd-3049,32'd-2043,32'd-5888,32'd2487,32'd3073,32'd8510,32'd1249,32'd7416,32'd-1949,32'd1204,32'd722,32'd5634,32'd2119,32'd9697,32'd161,32'd7519,32'd2961,32'd-2465,32'd-3432,32'd7543,32'd1385,32'd3088,32'd1373,32'd1715,32'd-4687,32'd-511,32'd2059,32'd-5600,32'd7480,32'd1156,32'd-9912,32'd-2221,32'd4733,32'd-4484,32'd7348,32'd9360,32'd-2597,32'd7045,32'd-1613};
    Wx[9]='{32'd1690,32'd2399,32'd1552,32'd-796,32'd3037,32'd759,32'd6308,32'd1051,32'd6289,32'd791,32'd424,32'd1627,32'd3354,32'd1691,32'd-830,32'd6474,32'd-2092,32'd-1599,32'd2351,32'd1685,32'd-2026,32'd1364,32'd-1158,32'd3222,32'd-687,32'd4741,32'd905,32'd1348,32'd2424,32'd45,32'd3813,32'd465,32'd-728,32'd256,32'd2097,32'd792,32'd6787,32'd598,32'd-2457,32'd-172,32'd-351,32'd-1011,32'd1875,32'd-1350,32'd8735,32'd2590,32'd8579,32'd412,32'd855,32'd331,32'd2705,32'd3276,32'd1148,32'd2427,32'd320,32'd-1724,32'd-1826,32'd5400,32'd306,32'd159,32'd-1478,32'd3649,32'd-3522,32'd5971,32'd9248,32'd-2430,32'd-4179,32'd-3105,32'd-642,32'd256,32'd786,32'd1958,32'd657,32'd6450,32'd2758,32'd-90,32'd-334,32'd-1019,32'd4755,32'd2171,32'd2291,32'd4860,32'd6269,32'd-182,32'd3947,32'd6103,32'd2232,32'd4829,32'd3908,32'd-2756,32'd2153,32'd7749,32'd3249,32'd-2670,32'd-6865,32'd-545,32'd3796,32'd-1386,32'd1268,32'd1752,32'd-3256,32'd1364,32'd2467,32'd-3811,32'd-2932,32'd-407,32'd8759,32'd1520,32'd3933,32'd8115,32'd-3964,32'd-3935,32'd-1445,32'd14375,32'd-5112,32'd-2294,32'd3913,32'd10009,32'd-4169,32'd4270,32'd692,32'd1481,32'd5419,32'd12158,32'd-481,32'd-8813,32'd1362,32'd764,32'd-200,32'd332,32'd689,32'd-4086,32'd-10283,32'd-16162,32'd3808,32'd-6728,32'd-291,32'd-6669,32'd1910,32'd-15771,32'd3945,32'd853,32'd-7890,32'd-6328,32'd-2570,32'd-3725,32'd205,32'd4675,32'd-4475,32'd3452,32'd1486,32'd9492,32'd1556,32'd-857,32'd2315,32'd13515,32'd-7841,32'd-5625,32'd4389,32'd2521,32'd-2064,32'd4689,32'd17119,32'd-1467,32'd-2095,32'd3093,32'd7050,32'd21953,32'd-3229,32'd-1520,32'd-3906,32'd8989,32'd-4167,32'd519,32'd-3420,32'd-3967,32'd-10478,32'd-12431,32'd89,32'd5014,32'd-715,32'd6103,32'd9877,32'd-5014,32'd892,32'd-73,32'd-2283,32'd4638,32'd5161,32'd473,32'd5219,32'd-1706,32'd-4831,32'd-1978,32'd-5541,32'd-2308,32'd-123,32'd-1634,32'd-3608,32'd-10449,32'd403,32'd1801,32'd102,32'd521,32'd320,32'd-1307,32'd5732,32'd-6650,32'd-3557,32'd-6215,32'd2226,32'd3186,32'd-3562,32'd8759,32'd3410,32'd-11298,32'd-9033,32'd3818,32'd4787,32'd1437,32'd-1064,32'd-2241,32'd-182,32'd-7016,32'd-4069,32'd1840,32'd-411,32'd-6,32'd-3520,32'd652,32'd-501,32'd5219,32'd8134,32'd645,32'd1793,32'd-98,32'd-7216,32'd3156,32'd1907,32'd-5336,32'd3593,32'd91,32'd-10849,32'd4992,32'd9057,32'd670,32'd5366,32'd4069,32'd1883,32'd-2092,32'd-2180,32'd7573,32'd2194,32'd-924,32'd-5449,32'd-7153,32'd4460,32'd1545,32'd-668,32'd-3156,32'd2265,32'd-3225,32'd6127,32'd3159,32'd6020,32'd-2423,32'd361,32'd7509,32'd469,32'd-1562,32'd-3388,32'd-5458,32'd-1394,32'd-300,32'd-113,32'd-2971,32'd10009,32'd2592,32'd-505,32'd4230,32'd-1429,32'd6992,32'd-4265,32'd-3281,32'd-1478,32'd-5737,32'd-841,32'd2612,32'd-3020,32'd-587,32'd-2651,32'd-2583,32'd1122,32'd1058,32'd11132,32'd-769,32'd9809,32'd-2597,32'd879,32'd3452,32'd-4465,32'd-3347,32'd-6967,32'd2413,32'd1685,32'd-7021,32'd2181,32'd-3828,32'd3544,32'd-3430,32'd1978,32'd4787,32'd1442,32'd3471,32'd2624,32'd-1684,32'd-11435,32'd-399,32'd-542,32'd2893,32'd-8520,32'd-1154,32'd3041,32'd-1889,32'd-2161,32'd2675,32'd-3618,32'd806,32'd2163,32'd5341,32'd4841,32'd5986,32'd2083,32'd780,32'd-8149,32'd-502,32'd-1697,32'd-2702,32'd5068,32'd-7211,32'd-598,32'd12910,32'd-2008,32'd7250,32'd3579,32'd-2493,32'd7368,32'd3847,32'd3015,32'd-4023,32'd215,32'd1822,32'd545,32'd5708,32'd-7851,32'd-6518,32'd-3981,32'd4174,32'd-5102,32'd1444,32'd5517,32'd1781,32'd11074,32'd-3378,32'd6494,32'd-3210,32'd-6708,32'd3366,32'd9511,32'd-532,32'd-4960,32'd1988,32'd-528,32'd852,32'd-5473,32'd-1284,32'd12500,32'd2385,32'd1381,32'd3947,32'd2927,32'd4897,32'd-117,32'd6040,32'd3347,32'd6635,32'd1936,32'd3571,32'd1234,32'd16884,32'd-2683,32'd-606,32'd1782,32'd3208,32'd4497,32'd-1173,32'd4904,32'd87,32'd2756,32'd5786};
    Wx[10]='{32'd1484,32'd4936,32'd-1878,32'd-189,32'd1380,32'd5444,32'd-132,32'd-1140,32'd-2003,32'd-319,32'd-6005,32'd-608,32'd-670,32'd6684,32'd-3054,32'd7548,32'd7153,32'd-5327,32'd854,32'd-2221,32'd-3513,32'd-4450,32'd-1843,32'd-3603,32'd68,32'd-2409,32'd830,32'd223,32'd2061,32'd1546,32'd558,32'd-4165,32'd3295,32'd-5483,32'd1159,32'd-2626,32'd-1405,32'd719,32'd5400,32'd1738,32'd-122,32'd1573,32'd7128,32'd-574,32'd4953,32'd-432,32'd-9213,32'd-612,32'd-847,32'd-1024,32'd1235,32'd-276,32'd-323,32'd-121,32'd4831,32'd4025,32'd1481,32'd-102,32'd3723,32'd3891,32'd2536,32'd168,32'd3662,32'd3012,32'd-2929,32'd-4113,32'd269,32'd-1525,32'd2258,32'd-1724,32'd-673,32'd1583,32'd6425,32'd3708,32'd-1917,32'd-1186,32'd5024,32'd4333,32'd-1406,32'd-1838,32'd-1087,32'd-398,32'd-290,32'd-5874,32'd903,32'd4291,32'd3386,32'd-517,32'd-448,32'd1855,32'd627,32'd3320,32'd-2812,32'd414,32'd-5869,32'd2044,32'd4792,32'd-1511,32'd-502,32'd-3090,32'd-6440,32'd12851,32'd-682,32'd5991,32'd4553,32'd-1195,32'd-226,32'd6816,32'd9350,32'd3256,32'd9106,32'd-12744,32'd-6201,32'd-8720,32'd6000,32'd3234,32'd21562,32'd473,32'd-3623,32'd46,32'd-4099,32'd-10517,32'd-978,32'd-6679,32'd-2103,32'd-403,32'd-35,32'd6333,32'd-2829,32'd-9575,32'd4499,32'd-5239,32'd16044,32'd-17041,32'd-4841,32'd-8041,32'd2082,32'd-149,32'd2308,32'd12460,32'd1506,32'd10576,32'd7148,32'd-15644,32'd10273,32'd-6982,32'd1964,32'd6728,32'd1342,32'd4763,32'd14755,32'd-3671,32'd-1486,32'd6713,32'd-1096,32'd-1368,32'd-662,32'd1676,32'd-839,32'd-2727,32'd888,32'd774,32'd-19042,32'd9379,32'd-14619,32'd2309,32'd-68,32'd-2531,32'd-45,32'd848,32'd286,32'd-2980,32'd3129,32'd11181,32'd2951,32'd5063,32'd783,32'd207,32'd6552,32'd-1582,32'd11347,32'd-1457,32'd15703,32'd-2127,32'd3874,32'd-6865,32'd-3801,32'd4008,32'd5014,32'd-873,32'd-5673,32'd1363,32'd1965,32'd5317,32'd-12109,32'd-5673,32'd677,32'd15751,32'd9482,32'd-17089,32'd-997,32'd-528,32'd-1557,32'd1218,32'd-1370,32'd-425,32'd-4426,32'd-5166,32'd-2241,32'd2180,32'd1781,32'd-3012,32'd-925,32'd798,32'd-1341,32'd3273,32'd11591,32'd-7861,32'd872,32'd-1113,32'd-2012,32'd-312,32'd-2978,32'd-3156,32'd-2575,32'd3005,32'd-14296,32'd-3232,32'd-4572,32'd-9975,32'd-4853,32'd2531,32'd-4526,32'd4970,32'd-4013,32'd-6948,32'd-5092,32'd-2951,32'd-1384,32'd-3764,32'd-7578,32'd3115,32'd2609,32'd-6748,32'd-13867,32'd-9213,32'd-4877,32'd-7392,32'd-3730,32'd4833,32'd-5795,32'd5825,32'd-2937,32'd-2504,32'd3508,32'd-6147,32'd-1673,32'd-2037,32'd-7133,32'd624,32'd1905,32'd1024,32'd1337,32'd-4194,32'd-4094,32'd-3347,32'd-3159,32'd-3112,32'd2255,32'd782,32'd2048,32'd7822,32'd1096,32'd2854,32'd-1860,32'd2088,32'd6796,32'd-1682,32'd5463,32'd6601,32'd-6098,32'd3811,32'd3637,32'd-279,32'd-6630,32'd1973,32'd-314,32'd-2514,32'd-1045,32'd-988,32'd-10507,32'd2753,32'd-1069,32'd-2177,32'd-2741,32'd-4592,32'd-6713,32'd160,32'd-7490,32'd137,32'd-4792,32'd2575,32'd-218,32'd-2041,32'd-469,32'd4353,32'd-15078,32'd-2443,32'd-7446,32'd-4235,32'd-483,32'd-1077,32'd-1147,32'd2199,32'd-114,32'd10234,32'd5917,32'd-6269,32'd-5981,32'd-8168,32'd1318,32'd-3012,32'd-1564,32'd-3796,32'd-3593,32'd4619,32'd-5654,32'd5087,32'd-5214,32'd-7104,32'd-462,32'd-2590,32'd-1184,32'd-3669,32'd-509,32'd-2976,32'd3659,32'd4860,32'd-4130,32'd-7192,32'd-910,32'd-5571,32'd5224,32'd-4694,32'd-5034,32'd-7919,32'd-10654,32'd-789,32'd-530,32'd957,32'd-8369,32'd2521,32'd-4509,32'd708,32'd4104,32'd1848,32'd-2717,32'd75,32'd-5092,32'd14736,32'd-4326,32'd-2526,32'd-10976,32'd-386,32'd4694,32'd-6181,32'd6992,32'd11425,32'd-7460,32'd-9541,32'd4731,32'd-4501,32'd4680,32'd-1771,32'd-5776,32'd388,32'd10078,32'd-3132,32'd2866,32'd10898,32'd-5693,32'd4860,32'd-6264,32'd2683,32'd14238,32'd4375,32'd31,32'd-1802,32'd229,32'd-1674,32'd-4987,32'd-903,32'd167,32'd5678,32'd-9326,32'd-4467,32'd4577,32'd-1669,32'd-5825,32'd-4819};
    Wx[11]='{32'd4357,32'd557,32'd2822,32'd1516,32'd-1109,32'd853,32'd2675,32'd-6962,32'd-1116,32'd-3830,32'd-1463,32'd-1154,32'd5825,32'd-831,32'd806,32'd7797,32'd301,32'd981,32'd-470,32'd3259,32'd-370,32'd-1463,32'd-4040,32'd906,32'd-377,32'd2374,32'd1541,32'd-882,32'd2459,32'd-177,32'd883,32'd480,32'd4526,32'd-2729,32'd7426,32'd872,32'd2980,32'd1082,32'd4978,32'd4350,32'd72,32'd618,32'd-3698,32'd1018,32'd1590,32'd3090,32'd-3823,32'd3483,32'd7470,32'd-903,32'd4941,32'd-2670,32'd-2322,32'd5659,32'd-1246,32'd6333,32'd1527,32'd-143,32'd-2463,32'd4697,32'd-826,32'd4487,32'd-1345,32'd3037,32'd-3164,32'd103,32'd3330,32'd-4023,32'd-2956,32'd-911,32'd114,32'd4592,32'd-5688,32'd2575,32'd4111,32'd4082,32'd9194,32'd-378,32'd128,32'd274,32'd947,32'd7236,32'd365,32'd-2824,32'd1051,32'd3811,32'd-1489,32'd105,32'd3830,32'd2202,32'd-1787,32'd-2203,32'd-883,32'd218,32'd-1986,32'd278,32'd276,32'd-5244,32'd-2312,32'd-1730,32'd-34,32'd-6918,32'd1457,32'd540,32'd-4467,32'd310,32'd1920,32'd-7827,32'd4616,32'd-104,32'd6040,32'd-1290,32'd-2817,32'd8247,32'd3342,32'd-7895,32'd3684,32'd8579,32'd4199,32'd3703,32'd-3828,32'd-3923,32'd8022,32'd-3723,32'd-2291,32'd3293,32'd2946,32'd-4541,32'd1658,32'd-4152,32'd3601,32'd-5,32'd-2111,32'd11035,32'd378,32'd4255,32'd6015,32'd-4030,32'd14121,32'd4475,32'd2673,32'd-3732,32'd-1838,32'd-2575,32'd6987,32'd4196,32'd-6616,32'd-5957,32'd3828,32'd4028,32'd9184,32'd-12861,32'd-1071,32'd-1361,32'd2159,32'd6918,32'd-3715,32'd-350,32'd960,32'd1257,32'd-3806,32'd-2218,32'd2109,32'd-2469,32'd-3762,32'd511,32'd-6977,32'd1506,32'd-1334,32'd1246,32'd7705,32'd12324,32'd-1906,32'd-10009,32'd6020,32'd-5805,32'd-2475,32'd-1125,32'd-1693,32'd-2443,32'd-1057,32'd-6416,32'd7138,32'd2978,32'd2792,32'd-9804,32'd459,32'd-7280,32'd9472,32'd-581,32'd10107,32'd7172,32'd15419,32'd-1649,32'd-11611,32'd-703,32'd1915,32'd-17880,32'd4079,32'd-4924,32'd942,32'd9843,32'd2274,32'd1329,32'd896,32'd433,32'd4680,32'd-6518,32'd-5371,32'd-279,32'd-1927,32'd1503,32'd-4123,32'd4699,32'd8618,32'd6704,32'd3991,32'd-4106,32'd-900,32'd1936,32'd-470,32'd-2839,32'd-3615,32'd149,32'd905,32'd-3735,32'd972,32'd-1394,32'd-868,32'd834,32'd798,32'd4284,32'd1857,32'd-3593,32'd-1547,32'd2211,32'd-1868,32'd-1855,32'd-5366,32'd-7836,32'd2159,32'd9208,32'd-1419,32'd1524,32'd12773,32'd118,32'd6547,32'd1738,32'd-1876,32'd2458,32'd-5600,32'd-8471,32'd-431,32'd1907,32'd-5820,32'd-6406,32'd-2293,32'd4494,32'd2727,32'd-9897,32'd1319,32'd1613,32'd-2181,32'd-6635,32'd10742,32'd-4716,32'd6665,32'd-13203,32'd-2707,32'd-3583,32'd-3869,32'd3969,32'd-3,32'd839,32'd5263,32'd278,32'd2165,32'd1997,32'd-1849,32'd-2060,32'd2143,32'd-1741,32'd-3859,32'd1083,32'd6699,32'd4152,32'd1239,32'd-4995,32'd-857,32'd-1163,32'd6914,32'd2011,32'd-3249,32'd-3452,32'd9516,32'd-376,32'd4641,32'd-554,32'd5239,32'd-1036,32'd-2144,32'd3769,32'd4157,32'd3115,32'd5004,32'd1080,32'd718,32'd-6044,32'd-7280,32'd-566,32'd-1396,32'd610,32'd740,32'd-737,32'd6611,32'd-875,32'd-2839,32'd437,32'd-5913,32'd3132,32'd1994,32'd449,32'd-1060,32'd1712,32'd5375,32'd-2773,32'd-530,32'd-7265,32'd-359,32'd-4838,32'd2204,32'd557,32'd-4108,32'd-4301,32'd2301,32'd6977,32'd4414,32'd278,32'd1589,32'd3029,32'd-4453,32'd712,32'd1060,32'd4924,32'd10761,32'd-4047,32'd2104,32'd3815,32'd6059,32'd885,32'd-1907,32'd-9345,32'd1340,32'd332,32'd-12001,32'd-3432,32'd-7534,32'd-2349,32'd-4699,32'd1427,32'd3288,32'd-301,32'd-1,32'd1486,32'd5346,32'd1047,32'd4924,32'd-2319,32'd-5947,32'd3210,32'd-3774,32'd-2812,32'd-2546,32'd283,32'd1807,32'd2188,32'd6552,32'd-3364,32'd-186,32'd-6396,32'd8671,32'd-9218,32'd-10898,32'd8876,32'd10751,32'd-148,32'd-3825,32'd-700,32'd1044,32'd3459,32'd2023,32'd-1007,32'd-213,32'd-3635,32'd8818,32'd4187,32'd6948,32'd704,32'd5488,32'd-560};
    Wx[12]='{32'd1596,32'd3435,32'd3120,32'd1920,32'd-694,32'd870,32'd1702,32'd-43,32'd2150,32'd-773,32'd-2768,32'd-1557,32'd-293,32'd1868,32'd2934,32'd11250,32'd-467,32'd-686,32'd-1103,32'd1023,32'd-1882,32'd-286,32'd-2470,32'd734,32'd-598,32'd-3518,32'd1994,32'd-1896,32'd9,32'd1778,32'd-44,32'd2656,32'd6689,32'd1749,32'd-1066,32'd2322,32'd3310,32'd9843,32'd811,32'd4941,32'd2749,32'd5131,32'd95,32'd5297,32'd-1646,32'd1229,32'd4775,32'd1506,32'd2526,32'd-756,32'd351,32'd888,32'd-1519,32'd1226,32'd4365,32'd358,32'd-62,32'd-2215,32'd3039,32'd1623,32'd-4118,32'd477,32'd2359,32'd-916,32'd-248,32'd-4687,32'd515,32'd1539,32'd-1789,32'd-5229,32'd-1011,32'd1739,32'd2208,32'd-939,32'd979,32'd194,32'd1926,32'd2980,32'd-1783,32'd-4475,32'd-2578,32'd-2055,32'd8574,32'd4858,32'd-5585,32'd6225,32'd16,32'd-305,32'd-1783,32'd4267,32'd370,32'd4123,32'd-2095,32'd-5185,32'd3037,32'd-34,32'd5170,32'd2595,32'd-2656,32'd938,32'd4997,32'd-17138,32'd-3720,32'd4465,32'd-3764,32'd1630,32'd-3210,32'd-14228,32'd-5449,32'd-2487,32'd-560,32'd-1590,32'd-6113,32'd8354,32'd8911,32'd6372,32'd6923,32'd4648,32'd-707,32'd-3200,32'd1095,32'd1600,32'd8427,32'd2770,32'd-3876,32'd8315,32'd569,32'd5449,32'd-1837,32'd642,32'd6054,32'd14755,32'd-19677,32'd14150,32'd5239,32'd-6396,32'd-873,32'd6748,32'd-125,32'd2067,32'd-5869,32'd10419,32'd-8164,32'd-4709,32'd-1613,32'd3129,32'd-8984,32'd-8559,32'd3312,32'd429,32'd18564,32'd-6894,32'd-609,32'd-2269,32'd-2993,32'd7885,32'd-528,32'd788,32'd-2349,32'd2692,32'd-3017,32'd1156,32'd-2534,32'd8315,32'd2534,32'd1201,32'd1798,32'd14638,32'd-3107,32'd-2402,32'd5078,32'd9262,32'd9736,32'd-1538,32'd89,32'd6625,32'd9111,32'd-2218,32'd1932,32'd3371,32'd-2917,32'd9345,32'd6166,32'd-8134,32'd-1983,32'd-20507,32'd-3266,32'd9023,32'd4204,32'd1717,32'd1319,32'd-3393,32'd3125,32'd637,32'd-12675,32'd-98,32'd-4030,32'd-9682,32'd-5966,32'd756,32'd-4326,32'd-4201,32'd3188,32'd4562,32'd3190,32'd-1352,32'd-8740,32'd-5737,32'd-1104,32'd-3356,32'd1356,32'd-1102,32'd3735,32'd6367,32'd-7788,32'd-4323,32'd2299,32'd-8017,32'd99,32'd-1556,32'd1395,32'd-153,32'd-3759,32'd-2668,32'd-4035,32'd-201,32'd-1361,32'd2109,32'd9418,32'd-568,32'd1213,32'd5073,32'd-5659,32'd-9560,32'd-1055,32'd1763,32'd-2558,32'd2485,32'd1925,32'd-5302,32'd-3049,32'd-3173,32'd187,32'd-287,32'd378,32'd6899,32'd2998,32'd855,32'd2756,32'd-2568,32'd4545,32'd6196,32'd-614,32'd4970,32'd2214,32'd-5229,32'd4748,32'd-3666,32'd94,32'd-4702,32'd5937,32'd-4213,32'd1616,32'd1402,32'd-3515,32'd-3005,32'd-3059,32'd1440,32'd-1990,32'd-941,32'd-1373,32'd7519,32'd5068,32'd2165,32'd1276,32'd598,32'd4970,32'd-7460,32'd3435,32'd5249,32'd2924,32'd5664,32'd8740,32'd1080,32'd-2856,32'd-9155,32'd1138,32'd-216,32'd1094,32'd1135,32'd8364,32'd11220,32'd-4499,32'd-4819,32'd-5839,32'd-1635,32'd-2133,32'd867,32'd-2275,32'd-6220,32'd-410,32'd-1600,32'd6157,32'd8076,32'd5820,32'd-3876,32'd-3669,32'd-1420,32'd-6342,32'd3269,32'd-737,32'd517,32'd3483,32'd2595,32'd3510,32'd2164,32'd-6391,32'd-1878,32'd255,32'd-5532,32'd3015,32'd3637,32'd-3913,32'd-4428,32'd-3525,32'd-1054,32'd-386,32'd-3718,32'd4677,32'd392,32'd760,32'd2032,32'd2998,32'd-5585,32'd-7636,32'd-1973,32'd-3261,32'd713,32'd2626,32'd-5166,32'd-5537,32'd5791,32'd5864,32'd12470,32'd4631,32'd7558,32'd-3425,32'd-2712,32'd6440,32'd-1408,32'd1613,32'd-2956,32'd7924,32'd3874,32'd645,32'd2321,32'd2531,32'd-10429,32'd487,32'd6958,32'd1711,32'd-5913,32'd-88,32'd1588,32'd-1314,32'd-4790,32'd-3999,32'd5917,32'd-5410,32'd-5590,32'd473,32'd7651,32'd-1652,32'd2491,32'd-1522,32'd7739,32'd2570,32'd135,32'd1522,32'd-3957,32'd-2226,32'd3747,32'd1738,32'd8774,32'd-1752,32'd3500,32'd489,32'd2153,32'd1474,32'd-1479,32'd-2016,32'd2413,32'd-339,32'd621,32'd11191,32'd-2631,32'd-11328,32'd-1295,32'd-6933,32'd-1114};
    Wx[13]='{32'd-690,32'd7216,32'd2331,32'd-437,32'd683,32'd-2758,32'd2795,32'd1540,32'd503,32'd960,32'd5849,32'd-396,32'd2420,32'd3854,32'd-3522,32'd1235,32'd1663,32'd3103,32'd2910,32'd1090,32'd-1198,32'd3093,32'd-2536,32'd2313,32'd3063,32'd1972,32'd3100,32'd3942,32'd2320,32'd-7060,32'd-1040,32'd-167,32'd5185,32'd2235,32'd5478,32'd3779,32'd-12,32'd825,32'd-7563,32'd2442,32'd4606,32'd4272,32'd-2846,32'd398,32'd-2563,32'd-648,32'd-1239,32'd3481,32'd3183,32'd-4550,32'd3308,32'd6181,32'd-704,32'd-2407,32'd-3808,32'd5234,32'd1737,32'd5917,32'd5283,32'd3217,32'd-254,32'd2827,32'd-745,32'd4111,32'd-1469,32'd-1989,32'd4614,32'd11699,32'd4211,32'd-1942,32'd-4680,32'd5175,32'd-4501,32'd38,32'd-1762,32'd2626,32'd1180,32'd3889,32'd1801,32'd6059,32'd3479,32'd1518,32'd9072,32'd-3203,32'd331,32'd2707,32'd-2315,32'd1497,32'd1215,32'd1378,32'd1574,32'd5683,32'd1513,32'd-3620,32'd3476,32'd7119,32'd1994,32'd1184,32'd5830,32'd8305,32'd-5156,32'd18837,32'd1055,32'd-2349,32'd-6772,32'd258,32'd13603,32'd-5122,32'd7900,32'd960,32'd-3454,32'd-4091,32'd7412,32'd17998,32'd4851,32'd2565,32'd7700,32'd-8461,32'd1202,32'd-1127,32'd-1148,32'd8159,32'd-2939,32'd9746,32'd7993,32'd5405,32'd6474,32'd-278,32'd-5390,32'd1324,32'd-6547,32'd4453,32'd-29218,32'd3254,32'd7060,32'd-1856,32'd12070,32'd2897,32'd11855,32'd-3999,32'd7832,32'd-13291,32'd-12744,32'd2492,32'd-13847,32'd5639,32'd-9536,32'd9555,32'd-6865,32'd746,32'd14892,32'd-11914,32'd-1834,32'd-25,32'd6196,32'd-582,32'd6650,32'd-1564,32'd2871,32'd5190,32'd3471,32'd6210,32'd9633,32'd348,32'd2490,32'd1564,32'd-2890,32'd-1934,32'd-1470,32'd-2249,32'd-3698,32'd-4645,32'd-5805,32'd2846,32'd-10927,32'd2083,32'd5971,32'd-2583,32'd11591,32'd-4104,32'd7636,32'd13369,32'd-4116,32'd8427,32'd-4938,32'd19501,32'd4770,32'd-3552,32'd1372,32'd1412,32'd6254,32'd-3217,32'd-6806,32'd-1783,32'd8588,32'd-555,32'd13134,32'd4970,32'd4814,32'd15566,32'd2687,32'd3676,32'd1882,32'd6186,32'd-850,32'd-794,32'd3562,32'd5913,32'd451,32'd-916,32'd2941,32'd120,32'd-1640,32'd-2338,32'd4038,32'd-5434,32'd-1657,32'd4641,32'd3090,32'd2288,32'd-994,32'd925,32'd-2360,32'd6650,32'd486,32'd-4204,32'd-1588,32'd1616,32'd-2133,32'd2517,32'd3376,32'd-4624,32'd-5410,32'd-119,32'd-9462,32'd-3928,32'd-4628,32'd-702,32'd-931,32'd-4873,32'd648,32'd-16396,32'd-2583,32'd4226,32'd3796,32'd-2739,32'd-16113,32'd-4272,32'd-2105,32'd3083,32'd-2315,32'd2614,32'd1343,32'd-2897,32'd-685,32'd-3469,32'd-3715,32'd2980,32'd10087,32'd-2023,32'd3359,32'd-5512,32'd-5209,32'd3586,32'd-4746,32'd-635,32'd3088,32'd-5991,32'd4919,32'd-2770,32'd-512,32'd-7192,32'd1290,32'd-566,32'd-1799,32'd-5292,32'd-1110,32'd96,32'd4055,32'd-4125,32'd1530,32'd4589,32'd-49,32'd1634,32'd-4592,32'd-1616,32'd-827,32'd131,32'd330,32'd246,32'd8930,32'd-9228,32'd5849,32'd-2480,32'd-3083,32'd1791,32'd8598,32'd-6889,32'd5810,32'd-689,32'd3457,32'd7470,32'd6367,32'd1785,32'd-3955,32'd4877,32'd9848,32'd1529,32'd8876,32'd-9052,32'd-1914,32'd3095,32'd5502,32'd2050,32'd-6411,32'd-2178,32'd9023,32'd-1899,32'd7958,32'd9111,32'd-1391,32'd-817,32'd384,32'd5751,32'd-5673,32'd3244,32'd852,32'd844,32'd12197,32'd7998,32'd4523,32'd3073,32'd-6840,32'd3754,32'd2626,32'd-7612,32'd1015,32'd3583,32'd296,32'd-1903,32'd4892,32'd3144,32'd2414,32'd-1865,32'd676,32'd-270,32'd7700,32'd-3730,32'd4716,32'd-84,32'd7797,32'd2539,32'd3564,32'd-1370,32'd-2355,32'd4316,32'd3200,32'd11718,32'd8183,32'd10654,32'd-407,32'd2492,32'd-2631,32'd5107,32'd-7016,32'd-5390,32'd10322,32'd-5405,32'd13164,32'd14628,32'd-2517,32'd4680,32'd3142,32'd-944,32'd-9472,32'd5615,32'd5908,32'd5249,32'd-4291,32'd5463,32'd8017,32'd7246,32'd6621,32'd-363,32'd2454,32'd-1061,32'd-3952,32'd366,32'd3054,32'd8281,32'd1717,32'd-15234,32'd493,32'd-710,32'd-10058,32'd3623,32'd7250,32'd2890,32'd3977,32'd8891};
    Wx[14]='{32'd3645,32'd8798,32'd1480,32'd-1552,32'd2460,32'd914,32'd5844,32'd614,32'd1738,32'd-974,32'd5673,32'd301,32'd-6533,32'd-2303,32'd-7783,32'd486,32'd-7075,32'd2722,32'd-467,32'd2580,32'd-4311,32'd-3745,32'd-364,32'd1625,32'd1246,32'd-1855,32'd1431,32'd-3063,32'd5791,32'd-2092,32'd-946,32'd-1861,32'd-3847,32'd-594,32'd2458,32'd-2866,32'd403,32'd-2099,32'd3930,32'd-2070,32'd-2269,32'd5312,32'd-2156,32'd-3120,32'd6977,32'd-2619,32'd-5107,32'd-4394,32'd-1708,32'd-566,32'd-4682,32'd1485,32'd-963,32'd-2442,32'd945,32'd88,32'd1041,32'd4145,32'd-1473,32'd-762,32'd2500,32'd-5268,32'd-6459,32'd-1491,32'd-853,32'd864,32'd-821,32'd657,32'd459,32'd303,32'd3518,32'd-4558,32'd1056,32'd-1677,32'd-1104,32'd-3527,32'd-5551,32'd-2398,32'd-5654,32'd4660,32'd-1566,32'd-481,32'd-1508,32'd1091,32'd726,32'd-862,32'd-2196,32'd2597,32'd-5214,32'd-2099,32'd-2597,32'd5068,32'd-3757,32'd2719,32'd2626,32'd-5078,32'd-2548,32'd1293,32'd971,32'd-1164,32'd1439,32'd1871,32'd-1008,32'd-4897,32'd-2077,32'd-1182,32'd7968,32'd4963,32'd-1240,32'd-4396,32'd4519,32'd7670,32'd-2961,32'd391,32'd9550,32'd423,32'd6782,32'd-3203,32'd-3024,32'd5473,32'd28,32'd-1296,32'd-693,32'd2421,32'd1347,32'd-3017,32'd389,32'd2890,32'd9086,32'd6401,32'd6503,32'd2404,32'd5175,32'd-891,32'd-3666,32'd-3388,32'd516,32'd-4440,32'd10966,32'd671,32'd-11416,32'd4555,32'd7958,32'd-5996,32'd-1289,32'd-4716,32'd1778,32'd3786,32'd6015,32'd-194,32'd-4333,32'd-2415,32'd1820,32'd-6142,32'd-3518,32'd-5688,32'd8994,32'd293,32'd-2851,32'd-502,32'd-3874,32'd-3549,32'd6733,32'd-3762,32'd6791,32'd62,32'd313,32'd4594,32'd-1629,32'd501,32'd881,32'd-1507,32'd-578,32'd6503,32'd-933,32'd-2486,32'd-3937,32'd-6303,32'd-3615,32'd-2388,32'd2998,32'd-8378,32'd2165,32'd640,32'd5566,32'd-9243,32'd188,32'd3989,32'd895,32'd-2666,32'd5937,32'd7216,32'd2963,32'd1694,32'd305,32'd1826,32'd1357,32'd-5415,32'd3105,32'd6059,32'd2445,32'd761,32'd2047,32'd993,32'd211,32'd-1844,32'd-1848,32'd-1693,32'd-2929,32'd-2322,32'd-2220,32'd97,32'd2966,32'd5449,32'd-5791,32'd4243,32'd11337,32'd3305,32'd-1300,32'd2054,32'd-2429,32'd-3903,32'd2810,32'd-2011,32'd-564,32'd-1207,32'd315,32'd-3872,32'd1111,32'd-2216,32'd-3825,32'd9189,32'd2858,32'd-352,32'd1627,32'd1644,32'd697,32'd-4125,32'd2280,32'd4877,32'd-1182,32'd-1884,32'd9091,32'd-4494,32'd1998,32'd1490,32'd4157,32'd1945,32'd5463,32'd5468,32'd11201,32'd1112,32'd-1040,32'd6674,32'd-3703,32'd5444,32'd5981,32'd4152,32'd-2187,32'd-16,32'd-3247,32'd7958,32'd-1411,32'd-1491,32'd-1605,32'd-4240,32'd-314,32'd11142,32'd870,32'd2023,32'd963,32'd-133,32'd6977,32'd5698,32'd1046,32'd1690,32'd-25,32'd154,32'd-5971,32'd1883,32'd-542,32'd3557,32'd5249,32'd-3225,32'd2563,32'd-962,32'd1943,32'd-956,32'd646,32'd2392,32'd-9379,32'd4638,32'd2998,32'd6411,32'd3996,32'd168,32'd-1442,32'd-4499,32'd-1999,32'd6557,32'd1185,32'd-198,32'd1115,32'd-505,32'd-1091,32'd4753,32'd-703,32'd9326,32'd-3996,32'd-6533,32'd3081,32'd-691,32'd204,32'd846,32'd-3308,32'd49,32'd1719,32'd2200,32'd-9677,32'd731,32'd-3354,32'd-3862,32'd-596,32'd-107,32'd1116,32'd2514,32'd-690,32'd-6523,32'd4213,32'd-4287,32'd-6601,32'd-856,32'd320,32'd-4489,32'd6083,32'd-4094,32'd-509,32'd-7705,32'd2320,32'd-2648,32'd-1407,32'd2788,32'd3603,32'd-7749,32'd-4116,32'd-4592,32'd1728,32'd-6376,32'd936,32'd2167,32'd-1381,32'd-434,32'd-1475,32'd138,32'd-6601,32'd6376,32'd3095,32'd-1341,32'd-1081,32'd-523,32'd-3974,32'd-733,32'd-6796,32'd-8764,32'd1839,32'd4614,32'd-2758,32'd13681,32'd7573,32'd-4577,32'd5786,32'd2316,32'd-1726,32'd871,32'd-8520,32'd-7939,32'd-4514,32'd-6274,32'd-5581,32'd5410,32'd-925,32'd-5727,32'd6938,32'd-1391,32'd4040,32'd533,32'd4453,32'd6225,32'd-2260,32'd-1500,32'd-8627,32'd-9008,32'd4733,32'd4274,32'd2186,32'd-5776,32'd-4172,32'd-756,32'd250,32'd1243};
    Wx[15]='{32'd-397,32'd-9116,32'd685,32'd-3522,32'd-3063,32'd-651,32'd-5478,32'd-880,32'd3334,32'd653,32'd-3054,32'd-3203,32'd191,32'd543,32'd-1318,32'd-3745,32'd-1540,32'd-4470,32'd1523,32'd974,32'd1870,32'd-4096,32'd-3876,32'd-547,32'd-2189,32'd-2849,32'd1014,32'd-1437,32'd-1870,32'd-4362,32'd2294,32'd3676,32'd-6621,32'd-5698,32'd273,32'd-2305,32'd1039,32'd-5229,32'd2399,32'd-2714,32'd-2437,32'd-1379,32'd2060,32'd-3066,32'd-4196,32'd676,32'd1319,32'd-2316,32'd1480,32'd625,32'd-2054,32'd-6440,32'd802,32'd6279,32'd-1162,32'd-11103,32'd1309,32'd1301,32'd-423,32'd-6440,32'd-737,32'd-346,32'd-6733,32'd674,32'd-1113,32'd1434,32'd-303,32'd6,32'd-4062,32'd-4460,32'd1799,32'd-3559,32'd1434,32'd-1390,32'd1235,32'd610,32'd-2685,32'd119,32'd-2104,32'd-4284,32'd1829,32'd254,32'd-2819,32'd-4140,32'd-5483,32'd-3420,32'd1906,32'd-2355,32'd484,32'd250,32'd1787,32'd-3444,32'd825,32'd-2099,32'd1265,32'd-874,32'd-5556,32'd-2438,32'd-3879,32'd-1881,32'd3562,32'd-11904,32'd-2397,32'd7539,32'd4450,32'd-1699,32'd567,32'd1633,32'd-7465,32'd884,32'd14228,32'd1779,32'd6333,32'd-516,32'd2452,32'd-1778,32'd1961,32'd-6474,32'd-2734,32'd-487,32'd-1203,32'd-1317,32'd8339,32'd-5781,32'd-2912,32'd-2276,32'd-2196,32'd1297,32'd-8447,32'd-1235,32'd3103,32'd-7006,32'd-5493,32'd-5405,32'd-6811,32'd1533,32'd-548,32'd-2995,32'd11757,32'd697,32'd2717,32'd-2384,32'd2526,32'd14833,32'd1160,32'd-10742,32'd-7055,32'd-5649,32'd-1672,32'd4548,32'd-14863,32'd127,32'd-571,32'd-14677,32'd-737,32'd7641,32'd2954,32'd-782,32'd4465,32'd-1743,32'd-120,32'd16162,32'd2145,32'd-395,32'd-5981,32'd-92,32'd1884,32'd-7387,32'd2490,32'd1115,32'd9208,32'd471,32'd3427,32'd4565,32'd3708,32'd12363,32'd7744,32'd-3129,32'd-16718,32'd-3237,32'd2839,32'd9199,32'd-6352,32'd656,32'd4331,32'd-8881,32'd2434,32'd-4692,32'd2753,32'd83,32'd-5361,32'd15117,32'd4121,32'd1929,32'd-7861,32'd-7089,32'd-2116,32'd9228,32'd-3991,32'd-3532,32'd-1701,32'd-4689,32'd-2148,32'd629,32'd2780,32'd1140,32'd7246,32'd420,32'd-4797,32'd503,32'd-3823,32'd-1312,32'd-2714,32'd-1146,32'd4863,32'd5024,32'd1842,32'd-1774,32'd2408,32'd-510,32'd2832,32'd-277,32'd-2514,32'd1875,32'd3874,32'd-2052,32'd-667,32'd494,32'd319,32'd5776,32'd-1206,32'd2561,32'd5766,32'd-974,32'd-3676,32'd-3642,32'd60,32'd-2866,32'd-5302,32'd-4670,32'd-597,32'd3459,32'd-3583,32'd-953,32'd-1802,32'd-4113,32'd833,32'd-2832,32'd4743,32'd-1358,32'd-4169,32'd-4416,32'd1022,32'd-7465,32'd-1674,32'd5888,32'd3537,32'd-3886,32'd-6069,32'd1997,32'd-3017,32'd-856,32'd-3342,32'd-1057,32'd-8701,32'd-1650,32'd-3083,32'd10156,32'd-2768,32'd-2995,32'd-3574,32'd5312,32'd4135,32'd-1809,32'd2805,32'd2490,32'd-7055,32'd-3151,32'd1120,32'd-1270,32'd3491,32'd-10195,32'd5468,32'd10146,32'd620,32'd1848,32'd-1358,32'd-3813,32'd-320,32'd130,32'd-2144,32'd4604,32'd-4807,32'd212,32'd1680,32'd3063,32'd922,32'd4453,32'd-3056,32'd-1306,32'd3918,32'd-6694,32'd-7895,32'd-5058,32'd-197,32'd-6113,32'd717,32'd637,32'd-4189,32'd5678,32'd207,32'd-1638,32'd-5620,32'd-3964,32'd-4118,32'd850,32'd-2766,32'd1127,32'd4658,32'd-1400,32'd-12363,32'd2432,32'd993,32'd-1242,32'd6240,32'd-705,32'd-971,32'd-6806,32'd-5625,32'd997,32'd-3869,32'd704,32'd-369,32'd-10263,32'd-3181,32'd-455,32'd1590,32'd-2995,32'd-6933,32'd-3276,32'd-2498,32'd-119,32'd705,32'd2568,32'd-2612,32'd-6044,32'd4160,32'd7441,32'd52,32'd1390,32'd-7558,32'd-4897,32'd2154,32'd4870,32'd-8935,32'd-12333,32'd-1538,32'd3813,32'd1888,32'd-5214,32'd1502,32'd-2073,32'd2462,32'd-10507,32'd-665,32'd2717,32'd-1629,32'd-1307,32'd-5009,32'd-4184,32'd3537,32'd2470,32'd374,32'd-4875,32'd1801,32'd-1998,32'd-7192,32'd2199,32'd-3068,32'd-5541,32'd8569,32'd-4514,32'd-942,32'd6552,32'd-14521,32'd-4482,32'd-1289,32'd-3046,32'd-3032,32'd2291,32'd2963,32'd6611,32'd-4885,32'd-2961,32'd-1746,32'd548,32'd2863,32'd-1231,32'd5034,32'd-3935};
    Wx[16]='{32'd736,32'd2915,32'd-1203,32'd137,32'd-946,32'd-639,32'd1292,32'd-2744,32'd-1357,32'd-106,32'd1485,32'd1206,32'd2800,32'd-462,32'd7426,32'd-301,32'd-4072,32'd1011,32'd-2357,32'd-1416,32'd2871,32'd-1794,32'd3891,32'd3063,32'd-1062,32'd-144,32'd3774,32'd1219,32'd1078,32'd3715,32'd-1789,32'd-2495,32'd2614,32'd2797,32'd936,32'd-5913,32'd-1336,32'd950,32'd3085,32'd2985,32'd1621,32'd509,32'd-957,32'd3237,32'd10039,32'd-869,32'd14951,32'd3117,32'd-1122,32'd-72,32'd4470,32'd2553,32'd2946,32'd2949,32'd-4155,32'd310,32'd3168,32'd3769,32'd-81,32'd-663,32'd-371,32'd-1016,32'd3923,32'd-603,32'd5615,32'd2181,32'd-320,32'd1524,32'd-2998,32'd3710,32'd1431,32'd4907,32'd-3754,32'd1335,32'd-627,32'd-173,32'd4765,32'd3884,32'd2690,32'd-6,32'd706,32'd-188,32'd3967,32'd4538,32'd4458,32'd4645,32'd-1578,32'd2561,32'd-993,32'd-210,32'd1350,32'd-1181,32'd1518,32'd1910,32'd1918,32'd-2514,32'd488,32'd1705,32'd-1156,32'd2416,32'd-1998,32'd-6684,32'd-2639,32'd-1411,32'd-262,32'd194,32'd-4121,32'd9492,32'd638,32'd-5957,32'd-548,32'd3239,32'd2995,32'd2770,32'd-154,32'd4453,32'd-9458,32'd90,32'd9091,32'd-3730,32'd4768,32'd-5297,32'd1750,32'd-7128,32'd-933,32'd3090,32'd-2218,32'd-9550,32'd-756,32'd7534,32'd-4309,32'd11962,32'd3588,32'd216,32'd5117,32'd-594,32'd-464,32'd-3120,32'd21328,32'd-10468,32'd-3723,32'd5917,32'd3830,32'd-2380,32'd5541,32'd16757,32'd-4367,32'd3327,32'd3022,32'd-3452,32'd-4016,32'd10976,32'd2331,32'd622,32'd2338,32'd-155,32'd-1408,32'd803,32'd-516,32'd-368,32'd971,32'd11562,32'd544,32'd-7568,32'd-2244,32'd-1988,32'd440,32'd-5083,32'd1917,32'd-1571,32'd-6826,32'd-5126,32'd3803,32'd-2197,32'd-1052,32'd-17187,32'd-3911,32'd15839,32'd1450,32'd342,32'd-5434,32'd-1922,32'd-1120,32'd7700,32'd5273,32'd-6997,32'd4189,32'd-7172,32'd2658,32'd725,32'd4724,32'd-9023,32'd-9555,32'd1187,32'd5527,32'd3740,32'd-12177,32'd11474,32'd-1348,32'd4130,32'd1909,32'd-218,32'd-2027,32'd-2521,32'd-116,32'd58,32'd-5776,32'd1364,32'd-17,32'd-1201,32'd-31,32'd-3063,32'd3913,32'd1972,32'd-10078,32'd-1726,32'd-1827,32'd637,32'd-4931,32'd809,32'd-823,32'd1744,32'd-1339,32'd2387,32'd2790,32'd3522,32'd2709,32'd-1484,32'd-1453,32'd-3591,32'd283,32'd-3247,32'd-3303,32'd2103,32'd714,32'd-9,32'd-1287,32'd3554,32'd405,32'd-4648,32'd3605,32'd362,32'd-4919,32'd4201,32'd-2198,32'd-1690,32'd1409,32'd-1748,32'd-930,32'd-1757,32'd-2973,32'd-2246,32'd36,32'd-7,32'd-5253,32'd-2529,32'd-6997,32'd2714,32'd-3713,32'd-1865,32'd-4023,32'd-8793,32'd-4436,32'd2578,32'd-3083,32'd1569,32'd-3894,32'd-12500,32'd-3039,32'd-1282,32'd-4384,32'd-1243,32'd3930,32'd-4545,32'd-2524,32'd-13701,32'd-3986,32'd228,32'd6210,32'd-1898,32'd-1018,32'd-5776,32'd2187,32'd-4770,32'd1141,32'd-8432,32'd-1925,32'd151,32'd991,32'd921,32'd-960,32'd-1470,32'd1995,32'd955,32'd2095,32'd-421,32'd-2275,32'd-4521,32'd-751,32'd-233,32'd5800,32'd-882,32'd-6020,32'd681,32'd726,32'd46,32'd538,32'd-1308,32'd-1237,32'd1490,32'd2832,32'd-3669,32'd-196,32'd2075,32'd-5502,32'd-6728,32'd-2529,32'd6875,32'd-4243,32'd2668,32'd5405,32'd3635,32'd-2,32'd2556,32'd6704,32'd125,32'd7055,32'd1475,32'd6171,32'd-3486,32'd1048,32'd-2320,32'd-3032,32'd6601,32'd3686,32'd-3144,32'd-592,32'd-1818,32'd1806,32'd25,32'd3430,32'd4211,32'd-955,32'd-839,32'd-4284,32'd-2663,32'd2626,32'd900,32'd-160,32'd612,32'd3312,32'd-5776,32'd3327,32'd1188,32'd1623,32'd5654,32'd2839,32'd-6240,32'd1981,32'd-1209,32'd-3383,32'd-5434,32'd-4370,32'd6318,32'd1970,32'd7934,32'd-1466,32'd-10927,32'd2114,32'd3181,32'd-289,32'd2714,32'd5507,32'd-2385,32'd-2861,32'd-9140,32'd5170,32'd-1398,32'd1462,32'd-7226,32'd-958,32'd-12636,32'd1832,32'd-5478,32'd4753,32'd-1409,32'd-6489,32'd2866,32'd-1400,32'd-3044,32'd1960,32'd2241,32'd3613,32'd-2138,32'd5126,32'd486,32'd4777,32'd-7597,32'd1490,32'd-1084};
    Wx[17]='{32'd-1833,32'd-3581,32'd869,32'd519,32'd-225,32'd2176,32'd-750,32'd-6733,32'd-1621,32'd2897,32'd-8520,32'd2563,32'd-3054,32'd-2622,32'd-3361,32'd-653,32'd-6054,32'd1139,32'd-1221,32'd2044,32'd603,32'd-4741,32'd-2888,32'd-483,32'd223,32'd-4167,32'd-3928,32'd-1605,32'd-2958,32'd-3645,32'd-2105,32'd-3696,32'd-4995,32'd-5317,32'd-6933,32'd2242,32'd-1524,32'd573,32'd-6489,32'd-472,32'd-1341,32'd-2578,32'd91,32'd1184,32'd1062,32'd-3244,32'd-12451,32'd3952,32'd-2103,32'd2280,32'd-5458,32'd-15693,32'd-4421,32'd-6152,32'd-5073,32'd-8662,32'd-1843,32'd-515,32'd-2980,32'd-5146,32'd-4958,32'd3220,32'd-627,32'd-3012,32'd-7685,32'd512,32'd-1353,32'd2705,32'd3920,32'd-1877,32'd-3708,32'd-416,32'd796,32'd-1015,32'd-847,32'd-538,32'd1127,32'd-3439,32'd-3854,32'd-454,32'd3281,32'd157,32'd-775,32'd-4194,32'd-274,32'd-3293,32'd628,32'd1380,32'd-2924,32'd-3559,32'd339,32'd-6992,32'd-2995,32'd464,32'd-6127,32'd-8818,32'd275,32'd-5468,32'd-527,32'd-7104,32'd839,32'd-2277,32'd-801,32'd932,32'd-1480,32'd-1580,32'd-2337,32'd225,32'd4277,32'd-7719,32'd-4541,32'd4501,32'd-4204,32'd5112,32'd794,32'd1420,32'd-2644,32'd5864,32'd-2714,32'd157,32'd-1286,32'd-3696,32'd2387,32'd713,32'd-4782,32'd-4382,32'd7758,32'd5795,32'd-6464,32'd-4916,32'd2673,32'd3498,32'd2427,32'd7646,32'd-2802,32'd3352,32'd-1129,32'd4680,32'd-9760,32'd-6132,32'd-5463,32'd-5209,32'd6357,32'd3972,32'd-1224,32'd-15537,32'd769,32'd450,32'd-44,32'd6699,32'd2697,32'd-12509,32'd-267,32'd9194,32'd-1296,32'd-2729,32'd1352,32'd-285,32'd-3305,32'd-445,32'd-6459,32'd-2795,32'd-6259,32'd-1645,32'd-9257,32'd-3264,32'd-1380,32'd-6,32'd-990,32'd-2990,32'd-7934,32'd-2736,32'd729,32'd-10966,32'd-564,32'd-1550,32'd15166,32'd3110,32'd-5151,32'd-3100,32'd2509,32'd-7001,32'd-486,32'd-720,32'd410,32'd4311,32'd-6845,32'd11572,32'd2479,32'd-6152,32'd-9599,32'd8862,32'd-480,32'd115,32'd-4296,32'd-7861,32'd3366,32'd-409,32'd1242,32'd-2238,32'd-413,32'd12402,32'd611,32'd1182,32'd758,32'd2827,32'd2775,32'd-4697,32'd4716,32'd2277,32'd-732,32'd63,32'd-353,32'd-2885,32'd12910,32'd6865,32'd-1911,32'd35,32'd3715,32'd1730,32'd687,32'd-629,32'd-3845,32'd-3779,32'd-447,32'd2462,32'd-1813,32'd-1419,32'd3315,32'd7050,32'd-893,32'd8608,32'd-365,32'd5512,32'd-1027,32'd-1665,32'd3466,32'd204,32'd353,32'd7407,32'd5839,32'd15371,32'd-10644,32'd1553,32'd-5874,32'd10761,32'd812,32'd-4665,32'd-609,32'd3686,32'd2905,32'd7324,32'd1912,32'd3332,32'd-1188,32'd7177,32'd5913,32'd833,32'd2858,32'd-3391,32'd-4089,32'd4382,32'd5131,32'd-5034,32'd4748,32'd3281,32'd3952,32'd-5024,32'd1927,32'd549,32'd1574,32'd6069,32'd-2412,32'd3259,32'd3410,32'd1674,32'd6259,32'd3823,32'd3154,32'd3388,32'd1239,32'd-4667,32'd4863,32'd-1541,32'd3513,32'd-3774,32'd492,32'd5092,32'd-686,32'd1281,32'd-54,32'd7954,32'd-6918,32'd-2302,32'd7426,32'd-3630,32'd5556,32'd-382,32'd-2272,32'd2626,32'd-507,32'd11650,32'd4370,32'd-343,32'd-1872,32'd2479,32'd4099,32'd-8613,32'd-3378,32'd1306,32'd-2452,32'd-641,32'd-4255,32'd-3603,32'd7099,32'd2015,32'd-550,32'd-932,32'd5244,32'd1629,32'd-2121,32'd-3051,32'd-4733,32'd1116,32'd115,32'd-1597,32'd-3232,32'd-34,32'd-3085,32'd1569,32'd-3176,32'd778,32'd3535,32'd3405,32'd-7670,32'd3601,32'd-3962,32'd-1593,32'd-1097,32'd1505,32'd5039,32'd4924,32'd-3967,32'd2148,32'd-2287,32'd1486,32'd-4165,32'd884,32'd-4963,32'd144,32'd-572,32'd-5175,32'd-9462,32'd-4897,32'd4951,32'd-2154,32'd3569,32'd-3061,32'd-101,32'd-1981,32'd-762,32'd3256,32'd1262,32'd-4243,32'd1763,32'd3198,32'd5512,32'd807,32'd4335,32'd-3840,32'd-1511,32'd9477,32'd-861,32'd5126,32'd4050,32'd5126,32'd4470,32'd-1146,32'd-6958,32'd32,32'd875,32'd-488,32'd1846,32'd9257,32'd5966,32'd994,32'd-2983,32'd8876,32'd-3957,32'd2429,32'd-5625,32'd3027,32'd-4926,32'd2673,32'd11816,32'd-5302,32'd7456,32'd-1334,32'd-972,32'd2670};
    Wx[18]='{32'd783,32'd1519,32'd-754,32'd873,32'd133,32'd1511,32'd3508,32'd-1226,32'd-687,32'd296,32'd-3156,32'd-753,32'd7260,32'd1734,32'd1590,32'd6166,32'd-1072,32'd-2519,32'd-504,32'd1973,32'd-3637,32'd-271,32'd-981,32'd143,32'd1170,32'd2026,32'd136,32'd639,32'd-3837,32'd3623,32'd-2749,32'd-9008,32'd-4487,32'd-563,32'd1164,32'd2475,32'd-1555,32'd243,32'd2402,32'd-1978,32'd1076,32'd-3154,32'd-297,32'd-292,32'd-5463,32'd2954,32'd-617,32'd-1159,32'd-1903,32'd-251,32'd2030,32'd-6103,32'd333,32'd-1086,32'd1701,32'd1993,32'd47,32'd-3083,32'd1785,32'd4992,32'd-272,32'd-3547,32'd-931,32'd3503,32'd-316,32'd1262,32'd-283,32'd1059,32'd1285,32'd265,32'd-1992,32'd2392,32'd-5629,32'd-3681,32'd2352,32'd-234,32'd1318,32'd3308,32'd1926,32'd-3615,32'd1604,32'd-1505,32'd1697,32'd6928,32'd-1977,32'd-1639,32'd19,32'd1224,32'd-1501,32'd1945,32'd514,32'd4162,32'd-341,32'd3410,32'd-4172,32'd3020,32'd13,32'd-2425,32'd-1926,32'd-2551,32'd-4121,32'd1857,32'd783,32'd-5727,32'd2917,32'd2795,32'd3249,32'd-3508,32'd-727,32'd-135,32'd7465,32'd-5180,32'd-366,32'd-2741,32'd-605,32'd-3615,32'd-82,32'd-3127,32'd-6298,32'd5283,32'd1053,32'd-1436,32'd-4394,32'd2502,32'd-3044,32'd5312,32'd1501,32'd-3442,32'd632,32'd-3781,32'd864,32'd6689,32'd-4567,32'd-7998,32'd83,32'd-895,32'd2352,32'd4018,32'd1216,32'd-4772,32'd2590,32'd-2504,32'd6547,32'd-9682,32'd-2546,32'd-4006,32'd12617,32'd5004,32'd-73,32'd2486,32'd8740,32'd334,32'd1414,32'd10419,32'd-4848,32'd169,32'd-1513,32'd1473,32'd-1824,32'd-1497,32'd-3974,32'd9028,32'd-8081,32'd6953,32'd-8203,32'd-1798,32'd-7578,32'd-3786,32'd-2810,32'd-1215,32'd-3125,32'd6005,32'd-2442,32'd-1037,32'd3505,32'd-6450,32'd10625,32'd-598,32'd6469,32'd-36,32'd-2021,32'd-2863,32'd-5976,32'd10117,32'd2534,32'd-5864,32'd1289,32'd3374,32'd3034,32'd-3103,32'd-2258,32'd-10341,32'd205,32'd2980,32'd-69,32'd-896,32'd-1816,32'd-9711,32'd-1347,32'd-806,32'd-4143,32'd-7285,32'd1436,32'd3193,32'd2478,32'd1480,32'd-3029,32'd3903,32'd3024,32'd-112,32'd8608,32'd-1883,32'd2900,32'd-2150,32'd-1422,32'd-1929,32'd-2534,32'd-470,32'd-1075,32'd3415,32'd-628,32'd-531,32'd3728,32'd989,32'd471,32'd1115,32'd3347,32'd-2116,32'd-1567,32'd-133,32'd-111,32'd9462,32'd3447,32'd4182,32'd3454,32'd-1448,32'd-1889,32'd1211,32'd-902,32'd915,32'd-2452,32'd-710,32'd8071,32'd3798,32'd-2888,32'd-3208,32'd-4741,32'd-1054,32'd455,32'd-2470,32'd-3906,32'd3508,32'd-337,32'd-4687,32'd-2039,32'd-2208,32'd-2048,32'd3684,32'd-1380,32'd-9394,32'd-1885,32'd-1223,32'd701,32'd-3356,32'd8173,32'd860,32'd-1323,32'd-9370,32'd467,32'd2352,32'd-4553,32'd-1063,32'd1469,32'd241,32'd2385,32'd4455,32'd-1550,32'd5625,32'd3935,32'd-3063,32'd1142,32'd6635,32'd1926,32'd2127,32'd4831,32'd2037,32'd2360,32'd-1948,32'd-1939,32'd4343,32'd-3159,32'd5410,32'd5400,32'd679,32'd-2651,32'd-3461,32'd-6015,32'd897,32'd-2313,32'd3103,32'd-894,32'd-1716,32'd-3674,32'd1823,32'd3867,32'd-2170,32'd-348,32'd-4609,32'd-851,32'd4848,32'd3427,32'd-1345,32'd5712,32'd2687,32'd1173,32'd622,32'd-2254,32'd1317,32'd6513,32'd-3420,32'd-2910,32'd-1549,32'd299,32'd749,32'd-2512,32'd2021,32'd1452,32'd-602,32'd-5678,32'd-650,32'd-5830,32'd2780,32'd-2722,32'd-341,32'd208,32'd-2590,32'd2131,32'd-2297,32'd4548,32'd4050,32'd-2043,32'd-1088,32'd568,32'd-3618,32'd-2147,32'd-3928,32'd-6958,32'd-3835,32'd3601,32'd-1829,32'd-6757,32'd596,32'd7241,32'd-7573,32'd-2100,32'd-466,32'd-3269,32'd-692,32'd-2739,32'd-6025,32'd-3537,32'd-2263,32'd-5156,32'd5180,32'd1654,32'd8813,32'd6049,32'd-6269,32'd-14736,32'd4252,32'd3391,32'd-1751,32'd3903,32'd281,32'd905,32'd-3579,32'd-2695,32'd2486,32'd1222,32'd-141,32'd-1807,32'd673,32'd2521,32'd-551,32'd7104,32'd3476,32'd1604,32'd165,32'd225,32'd-6313,32'd-1926,32'd-2304,32'd2463,32'd3857,32'd-5029,32'd-3286,32'd-326,32'd-4770,32'd-181,32'd-2401};
    Wx[19]='{32'd200,32'd-3798,32'd1516,32'd458,32'd-2873,32'd-1663,32'd4665,32'd1318,32'd-353,32'd-3630,32'd-1562,32'd306,32'd-3505,32'd-4011,32'd-861,32'd2868,32'd1516,32'd211,32'd-791,32'd292,32'd957,32'd127,32'd1074,32'd-582,32'd1395,32'd2592,32'd2327,32'd3029,32'd1273,32'd733,32'd1130,32'd-3430,32'd5561,32'd2595,32'd-4111,32'd1278,32'd177,32'd-1202,32'd1036,32'd1152,32'd-1170,32'd1582,32'd833,32'd-3571,32'd-1673,32'd-2236,32'd-1837,32'd880,32'd-1021,32'd-2314,32'd-1490,32'd5263,32'd1934,32'd7968,32'd4194,32'd739,32'd21,32'd2973,32'd265,32'd2097,32'd2680,32'd2239,32'd-5092,32'd-2110,32'd887,32'd-1889,32'd389,32'd1933,32'd-1860,32'd-1392,32'd-4387,32'd-488,32'd-3557,32'd-1155,32'd-869,32'd1029,32'd3061,32'd-1757,32'd-2590,32'd-858,32'd-2023,32'd-8154,32'd-1837,32'd-1550,32'd-3085,32'd-3088,32'd133,32'd107,32'd388,32'd-2272,32'd-6552,32'd6000,32'd-1408,32'd-1553,32'd540,32'd-458,32'd-3173,32'd-40,32'd5566,32'd-4370,32'd2176,32'd-1356,32'd-57,32'd12978,32'd-2939,32'd1397,32'd3845,32'd473,32'd153,32'd-220,32'd9199,32'd1795,32'd6459,32'd10869,32'd-5595,32'd5751,32'd-4460,32'd-2070,32'd467,32'd2573,32'd1285,32'd6206,32'd-6489,32'd13437,32'd1651,32'd-9995,32'd-2167,32'd808,32'd2320,32'd-8081,32'd6093,32'd592,32'd-994,32'd-4033,32'd-2486,32'd-275,32'd-1019,32'd-9301,32'd-5932,32'd13740,32'd4975,32'd-7412,32'd-1414,32'd15234,32'd11152,32'd-632,32'd-4924,32'd5224,32'd-22968,32'd716,32'd10419,32'd8139,32'd9150,32'd-9438,32'd-1094,32'd-4006,32'd5048,32'd-2463,32'd-356,32'd1342,32'd8017,32'd-161,32'd-6132,32'd8666,32'd15380,32'd1173,32'd-811,32'd-2697,32'd2580,32'd-3232,32'd-3395,32'd-3854,32'd-4482,32'd-12880,32'd1124,32'd-3508,32'd-3652,32'd-2900,32'd-13662,32'd-7500,32'd5375,32'd11962,32'd3635,32'd-1845,32'd3168,32'd-6508,32'd957,32'd3840,32'd-2963,32'd-1468,32'd3662,32'd-7192,32'd-4758,32'd-355,32'd-1925,32'd9140,32'd4736,32'd3571,32'd10654,32'd-24199,32'd-2568,32'd16152,32'd-2465,32'd3818,32'd-1467,32'd-23,32'd2229,32'd4128,32'd-460,32'd143,32'd-1798,32'd-642,32'd-3295,32'd2695,32'd-2631,32'd4145,32'd9165,32'd-3762,32'd160,32'd2338,32'd1472,32'd-1050,32'd-1557,32'd-5327,32'd-3847,32'd-1232,32'd-3598,32'd-2680,32'd-8725,32'd5771,32'd-1311,32'd-6298,32'd-850,32'd-1523,32'd1721,32'd-1508,32'd-1343,32'd-3259,32'd-1109,32'd3542,32'd-545,32'd2768,32'd12197,32'd-3784,32'd-5522,32'd-1035,32'd4943,32'd894,32'd3002,32'd-513,32'd-375,32'd-947,32'd8022,32'd6835,32'd3583,32'd8500,32'd3063,32'd-2490,32'd250,32'd162,32'd185,32'd-5400,32'd-3930,32'd-5190,32'd-1127,32'd52,32'd2312,32'd6289,32'd878,32'd-1395,32'd1855,32'd-5517,32'd-4140,32'd5473,32'd-3139,32'd-5224,32'd7075,32'd-1403,32'd5263,32'd725,32'd1102,32'd-1881,32'd-676,32'd-936,32'd769,32'd3969,32'd528,32'd-1877,32'd6318,32'd2490,32'd-6347,32'd-2763,32'd-3674,32'd1887,32'd-2653,32'd-2600,32'd-5629,32'd-13925,32'd591,32'd-1490,32'd-1590,32'd9047,32'd-6665,32'd-3854,32'd-6582,32'd-18505,32'd-4914,32'd8422,32'd5947,32'd8173,32'd-439,32'd1439,32'd6005,32'd-1794,32'd-1733,32'd3610,32'd8798,32'd-1977,32'd-4379,32'd1687,32'd-12392,32'd-5493,32'd-3039,32'd872,32'd-2358,32'd3432,32'd4260,32'd-5004,32'd7124,32'd8715,32'd4460,32'd2276,32'd-1810,32'd-4477,32'd4418,32'd278,32'd172,32'd-3100,32'd-1651,32'd-4162,32'd2812,32'd2238,32'd1049,32'd4772,32'd3059,32'd1585,32'd-5668,32'd-891,32'd-9121,32'd-567,32'd9077,32'd-2100,32'd1856,32'd-994,32'd-5961,32'd188,32'd3144,32'd-5097,32'd3061,32'd6230,32'd2435,32'd7421,32'd97,32'd-2502,32'd-1152,32'd-14062,32'd-2634,32'd-1921,32'd2130,32'd-6640,32'd1674,32'd-1607,32'd-7832,32'd2670,32'd-3825,32'd-1222,32'd5126,32'd-1353,32'd5087,32'd7631,32'd5380,32'd-2150,32'd483,32'd1968,32'd477,32'd3583,32'd-92,32'd-3315,32'd2167,32'd585,32'd-8017,32'd1682,32'd-1915,32'd10234,32'd1628,32'd4785,32'd-1846,32'd3388,32'd7836,32'd-2670};
    Wx[20]='{32'd531,32'd-6928,32'd-305,32'd-2481,32'd3520,32'd1820,32'd-526,32'd7148,32'd1315,32'd35,32'd1309,32'd-2758,32'd-1826,32'd-2456,32'd1812,32'd0,32'd-1599,32'd2858,32'd3134,32'd-218,32'd2490,32'd4448,32'd-2082,32'd57,32'd-1734,32'd-1541,32'd1307,32'd2015,32'd4130,32'd-3859,32'd256,32'd5698,32'd928,32'd-2441,32'd2368,32'd2196,32'd3369,32'd1624,32'd932,32'd-1270,32'd1142,32'd-1367,32'd1036,32'd-1439,32'd-2448,32'd3557,32'd-8564,32'd-4560,32'd4934,32'd145,32'd4577,32'd1804,32'd597,32'd-2155,32'd-3247,32'd-5351,32'd-1887,32'd-2133,32'd-686,32'd1378,32'd3,32'd5649,32'd-5698,32'd498,32'd8813,32'd-3395,32'd1348,32'd2437,32'd3208,32'd1414,32'd6572,32'd-4372,32'd-3437,32'd-4909,32'd1904,32'd-40,32'd-1020,32'd409,32'd5288,32'd3225,32'd-371,32'd-5571,32'd1782,32'd-4570,32'd-1403,32'd-3295,32'd122,32'd-761,32'd1577,32'd-1529,32'd797,32'd-6025,32'd-395,32'd2086,32'd936,32'd3903,32'd-4453,32'd2514,32'd-458,32'd-211,32'd-155,32'd2602,32'd1326,32'd-3613,32'd13564,32'd-1744,32'd-3610,32'd3793,32'd-2805,32'd8120,32'd-9833,32'd-3774,32'd1821,32'd1352,32'd-8974,32'd-5625,32'd-2034,32'd546,32'd5170,32'd-433,32'd5327,32'd303,32'd3259,32'd2902,32'd7412,32'd-10439,32'd2333,32'd-1383,32'd-3542,32'd4526,32'd-533,32'd9589,32'd-5585,32'd-3964,32'd3093,32'd2690,32'd2401,32'd400,32'd7529,32'd-4475,32'd-1113,32'd-15957,32'd9379,32'd9731,32'd9257,32'd2493,32'd6333,32'd-10341,32'd1190,32'd5742,32'd-1285,32'd-12617,32'd8041,32'd-8403,32'd8447,32'd1453,32'd4326,32'd5239,32'd3300,32'd-1256,32'd6577,32'd7226,32'd306,32'd3840,32'd-3071,32'd-3234,32'd-2604,32'd8588,32'd1063,32'd-2318,32'd2551,32'd-3425,32'd-2139,32'd22343,32'd155,32'd-1911,32'd-15146,32'd7026,32'd-6088,32'd4489,32'd-3190,32'd5976,32'd-872,32'd10175,32'd-10253,32'd4790,32'd1129,32'd4548,32'd7,32'd322,32'd8686,32'd637,32'd1362,32'd903,32'd-2893,32'd2575,32'd-5966,32'd4404,32'd5419,32'd-15468,32'd-1547,32'd-6479,32'd2287,32'd4204,32'd7866,32'd2082,32'd6181,32'd-7695,32'd-4260,32'd591,32'd-2041,32'd1918,32'd2435,32'd-1398,32'd11582,32'd-4738,32'd-736,32'd511,32'd1335,32'd-5278,32'd472,32'd-997,32'd6708,32'd2060,32'd1004,32'd2607,32'd-3322,32'd4323,32'd4416,32'd5922,32'd-1246,32'd-243,32'd-2863,32'd-1257,32'd-545,32'd1923,32'd-4658,32'd-1552,32'd-2495,32'd678,32'd6064,32'd-6650,32'd-8994,32'd3183,32'd26738,32'd-2524,32'd-9418,32'd4848,32'd-1141,32'd3554,32'd1291,32'd4255,32'd3076,32'd-6318,32'd1788,32'd3142,32'd4819,32'd-217,32'd-807,32'd3398,32'd-1270,32'd7060,32'd4597,32'd-5810,32'd-6821,32'd-2304,32'd1291,32'd-1903,32'd-1636,32'd-2888,32'd4509,32'd4738,32'd3300,32'd-1674,32'd3715,32'd-1364,32'd-2315,32'd-2995,32'd210,32'd5708,32'd836,32'd-9956,32'd2478,32'd2939,32'd-5439,32'd7128,32'd1517,32'd-3281,32'd5087,32'd-1148,32'd1271,32'd306,32'd-255,32'd1097,32'd-2382,32'd1179,32'd1530,32'd-4968,32'd2279,32'd-3381,32'd-3000,32'd3825,32'd181,32'd4040,32'd6010,32'd5229,32'd9316,32'd-1965,32'd-2778,32'd1021,32'd-1270,32'd5200,32'd-1136,32'd5742,32'd2014,32'd-2580,32'd-4982,32'd2556,32'd133,32'd1624,32'd-302,32'd384,32'd4428,32'd1881,32'd1180,32'd-2429,32'd-2666,32'd3793,32'd7836,32'd3540,32'd-3261,32'd2030,32'd-3176,32'd-2059,32'd-1679,32'd1768,32'd-3522,32'd-29,32'd-8168,32'd22,32'd4548,32'd-5014,32'd1740,32'd7363,32'd13085,32'd-622,32'd-2792,32'd2336,32'd8945,32'd-913,32'd5952,32'd-1121,32'd3395,32'd-4072,32'd5141,32'd-1486,32'd3559,32'd1182,32'd-1861,32'd-2773,32'd2308,32'd9404,32'd2648,32'd4790,32'd3020,32'd-789,32'd2424,32'd4855,32'd14248,32'd11826,32'd1864,32'd6176,32'd3757,32'd-780,32'd1754,32'd4450,32'd4624,32'd4,32'd-1115,32'd7470,32'd6650,32'd-3122,32'd2443,32'd9160,32'd-8583,32'd5449,32'd2822,32'd1683,32'd-1815,32'd12880,32'd58,32'd2003,32'd-1575,32'd16083,32'd5288,32'd3322,32'd-3317,32'd6640,32'd1873,32'd3105};
    Wx[21]='{32'd467,32'd-5493,32'd486,32'd-1389,32'd25,32'd536,32'd-3127,32'd-2384,32'd397,32'd-3715,32'd3564,32'd1763,32'd667,32'd993,32'd-7963,32'd-4865,32'd6816,32'd3107,32'd3027,32'd1428,32'd3298,32'd-3933,32'd-2717,32'd-1317,32'd1790,32'd-1167,32'd3439,32'd1943,32'd-4160,32'd-2731,32'd649,32'd-2344,32'd3178,32'd1243,32'd-2243,32'd-1193,32'd-308,32'd-443,32'd2426,32'd5092,32'd-546,32'd-654,32'd-3269,32'd-4099,32'd-7504,32'd1162,32'd2050,32'd6772,32'd827,32'd2685,32'd-1096,32'd-1541,32'd3977,32'd415,32'd2744,32'd4357,32'd-1851,32'd4399,32'd341,32'd2919,32'd-541,32'd4223,32'd-4624,32'd4460,32'd-8305,32'd460,32'd3059,32'd1268,32'd280,32'd2954,32'd2025,32'd-1034,32'd729,32'd1551,32'd-224,32'd-656,32'd3000,32'd292,32'd2346,32'd-1966,32'd50,32'd-23,32'd-4672,32'd-7485,32'd142,32'd1881,32'd3269,32'd-3225,32'd-1588,32'd98,32'd2795,32'd2226,32'd-2402,32'd-1024,32'd89,32'd-170,32'd-670,32'd3471,32'd299,32'd1325,32'd2802,32'd7260,32'd3261,32'd4821,32'd9946,32'd-2010,32'd-2854,32'd11582,32'd-1385,32'd3376,32'd-7690,32'd-309,32'd2653,32'd-8037,32'd6533,32'd819,32'd-3635,32'd-5375,32'd-987,32'd-3364,32'd2766,32'd-8056,32'd-207,32'd-3784,32'd-985,32'd54,32'd337,32'd-2452,32'd-15419,32'd-3115,32'd2968,32'd15312,32'd20781,32'd-6406,32'd-3566,32'd2854,32'd402,32'd3159,32'd-810,32'd-2175,32'd-4760,32'd15703,32'd-6313,32'd-14589,32'd-10742,32'd-6181,32'd-14648,32'd11318,32'd-398,32'd3215,32'd2807,32'd10917,32'd2193,32'd-5732,32'd2939,32'd-9194,32'd-3212,32'd1824,32'd6464,32'd-2912,32'd4372,32'd35,32'd1467,32'd-4436,32'd4521,32'd256,32'd-5429,32'd-7607,32'd450,32'd-791,32'd9204,32'd-11816,32'd-3078,32'd2257,32'd-2785,32'd6000,32'd-7841,32'd12695,32'd1733,32'd-7177,32'd2250,32'd3508,32'd-6796,32'd-164,32'd-8168,32'd12958,32'd362,32'd-5507,32'd3593,32'd7788,32'd6611,32'd3159,32'd-7622,32'd-3498,32'd-180,32'd-2403,32'd8295,32'd-1013,32'd10703,32'd-14033,32'd-1184,32'd13222,32'd647,32'd2308,32'd100,32'd772,32'd66,32'd9326,32'd-4819,32'd2136,32'd1580,32'd4338,32'd930,32'd-11464,32'd4116,32'd2565,32'd10371,32'd7031,32'd2193,32'd-2158,32'd4445,32'd1624,32'd5244,32'd-4472,32'd5478,32'd1183,32'd-6948,32'd1499,32'd5566,32'd5488,32'd-6479,32'd4873,32'd-4423,32'd5839,32'd-3701,32'd-4516,32'd203,32'd-2827,32'd5268,32'd3300,32'd-2702,32'd6425,32'd6821,32'd-12744,32'd9287,32'd4477,32'd-4260,32'd-2912,32'd-1929,32'd3969,32'd3811,32'd3725,32'd-2209,32'd8593,32'd8671,32'd-941,32'd6054,32'd-96,32'd3002,32'd4838,32'd-3242,32'd-6113,32'd5410,32'd2961,32'd6284,32'd-848,32'd6069,32'd16826,32'd-163,32'd1623,32'd492,32'd7324,32'd-10,32'd8930,32'd108,32'd1468,32'd6464,32'd-345,32'd-3464,32'd304,32'd3259,32'd2335,32'd2252,32'd-869,32'd474,32'd-254,32'd-556,32'd2341,32'd3178,32'd1567,32'd-3483,32'd3767,32'd3732,32'd567,32'd-449,32'd1054,32'd3952,32'd2341,32'd3808,32'd2966,32'd-1906,32'd8842,32'd35,32'd-2797,32'd-3083,32'd9560,32'd-3239,32'd9873,32'd1956,32'd-253,32'd1201,32'd2944,32'd-6000,32'd-1320,32'd-4367,32'd-1026,32'd3034,32'd-2565,32'd3876,32'd-7343,32'd7753,32'd1485,32'd-1848,32'd-1665,32'd-4494,32'd4946,32'd245,32'd323,32'd7880,32'd-1586,32'd5981,32'd4807,32'd-3884,32'd475,32'd-336,32'd4345,32'd6821,32'd-1508,32'd-1778,32'd3447,32'd-214,32'd4284,32'd388,32'd-7885,32'd-948,32'd5107,32'd5263,32'd4753,32'd-4238,32'd3229,32'd9433,32'd7138,32'd-6787,32'd433,32'd1157,32'd-7441,32'd7075,32'd1373,32'd-4116,32'd1250,32'd3393,32'd6689,32'd435,32'd-4108,32'd-2023,32'd-872,32'd6372,32'd8261,32'd-15546,32'd-4985,32'd-955,32'd12431,32'd2866,32'd7495,32'd5693,32'd2298,32'd-7197,32'd-3251,32'd1395,32'd-4187,32'd-2493,32'd-3845,32'd2010,32'd17861,32'd-1257,32'd7265,32'd-3747,32'd6586,32'd4086,32'd3759,32'd-635,32'd1605,32'd-1172,32'd-1002,32'd-4477,32'd7763,32'd7255,32'd9233,32'd-122,32'd1674};
    Wx[22]='{32'd-3217,32'd-5507,32'd670,32'd83,32'd-6831,32'd-2100,32'd2285,32'd845,32'd-1473,32'd-1005,32'd-1380,32'd304,32'd1271,32'd-467,32'd751,32'd-1950,32'd6542,32'd-549,32'd1717,32'd589,32'd215,32'd1189,32'd920,32'd3764,32'd-2543,32'd2858,32'd-2386,32'd2103,32'd8237,32'd-3842,32'd1379,32'd4741,32'd6674,32'd5151,32'd-3327,32'd-3178,32'd-117,32'd-1644,32'd1359,32'd-1094,32'd1026,32'd-8330,32'd3962,32'd-1383,32'd415,32'd-3461,32'd407,32'd-4367,32'd1258,32'd1640,32'd-7749,32'd-3557,32'd5585,32'd-3750,32'd498,32'd-4238,32'd241,32'd3459,32'd-2041,32'd-164,32'd1017,32'd6445,32'd-1545,32'd-826,32'd-4770,32'd295,32'd1607,32'd-1036,32'd-2534,32'd-1009,32'd-2298,32'd-1307,32'd4409,32'd-3139,32'd1945,32'd1745,32'd4831,32'd5415,32'd1282,32'd-2614,32'd3701,32'd4907,32'd-1666,32'd-1533,32'd-1971,32'd3598,32'd343,32'd-1207,32'd-3005,32'd5000,32'd1871,32'd-3098,32'd1859,32'd-445,32'd-842,32'd-853,32'd-3891,32'd1348,32'd5253,32'd841,32'd-4211,32'd-11201,32'd-3044,32'd-2756,32'd977,32'd-436,32'd8510,32'd-2797,32'd18,32'd3239,32'd-5327,32'd4624,32'd7602,32'd629,32'd16689,32'd-1229,32'd-437,32'd-11132,32'd8491,32'd1259,32'd691,32'd6811,32'd1627,32'd-1795,32'd-164,32'd973,32'd-11,32'd-997,32'd4260,32'd10898,32'd797,32'd2386,32'd8291,32'd3398,32'd4191,32'd300,32'd-1821,32'd-2802,32'd8510,32'd-9301,32'd-1608,32'd-6782,32'd-409,32'd10107,32'd1839,32'd2998,32'd299,32'd11357,32'd449,32'd-1414,32'd-3996,32'd4863,32'd10273,32'd-2285,32'd526,32'd5332,32'd12109,32'd-6342,32'd11181,32'd2279,32'd-3745,32'd10419,32'd4169,32'd-3852,32'd5825,32'd-1082,32'd360,32'd-19550,32'd1911,32'd-2098,32'd10048,32'd-2266,32'd3889,32'd2880,32'd-3410,32'd874,32'd11826,32'd3857,32'd-9179,32'd-9526,32'd-4638,32'd-6933,32'd4291,32'd8945,32'd3864,32'd-367,32'd6157,32'd2366,32'd-2407,32'd-523,32'd10605,32'd-2155,32'd-7211,32'd-3100,32'd4045,32'd-525,32'd-11513,32'd9531,32'd-2116,32'd-4699,32'd971,32'd5771,32'd-1893,32'd2073,32'd-7285,32'd-1501,32'd-3486,32'd1143,32'd843,32'd-1778,32'd-2430,32'd3073,32'd-2099,32'd-3056,32'd4211,32'd-4260,32'd-10742,32'd3103,32'd-3254,32'd4326,32'd2172,32'd-1164,32'd-6210,32'd2580,32'd4450,32'd-2687,32'd4812,32'd-3376,32'd-1492,32'd2026,32'd328,32'd-17207,32'd4372,32'd-6772,32'd4104,32'd4929,32'd-2296,32'd-3435,32'd-2475,32'd-3796,32'd5327,32'd-7050,32'd4711,32'd-3269,32'd10810,32'd-4948,32'd2303,32'd707,32'd-1766,32'd4025,32'd-11132,32'd-121,32'd1765,32'd-4086,32'd4643,32'd2326,32'd-487,32'd245,32'd1436,32'd-892,32'd1936,32'd-2509,32'd-6411,32'd5322,32'd-7421,32'd683,32'd806,32'd-16689,32'd-392,32'd-3137,32'd6308,32'd-3527,32'd1721,32'd5107,32'd-681,32'd-1696,32'd-4277,32'd-10693,32'd1597,32'd-5068,32'd-82,32'd-6630,32'd9282,32'd-4787,32'd1649,32'd-3349,32'd-310,32'd105,32'd5874,32'd-2020,32'd2983,32'd-2993,32'd5981,32'd-690,32'd8964,32'd1435,32'd-3623,32'd-6474,32'd-805,32'd2000,32'd-808,32'd-4113,32'd3261,32'd-9350,32'd-6943,32'd-6147,32'd2015,32'd3959,32'd3073,32'd-4377,32'd2136,32'd-1055,32'd1394,32'd-9814,32'd-7539,32'd-4299,32'd-2039,32'd5512,32'd4160,32'd8564,32'd-10302,32'd-1154,32'd-571,32'd3537,32'd3007,32'd3479,32'd2927,32'd-6694,32'd7500,32'd11728,32'd1751,32'd-6596,32'd3576,32'd-5458,32'd-1489,32'd1715,32'd-2022,32'd-10820,32'd-6484,32'd-1596,32'd2770,32'd-7504,32'd1948,32'd-4340,32'd7846,32'd-8193,32'd-1285,32'd2244,32'd-10302,32'd7153,32'd657,32'd-4379,32'd2519,32'd-7475,32'd3381,32'd1652,32'd4260,32'd10234,32'd1241,32'd2661,32'd1483,32'd1956,32'd790,32'd4233,32'd-6083,32'd-2619,32'd-7490,32'd-10810,32'd-11894,32'd-6005,32'd5874,32'd-4274,32'd-7221,32'd1906,32'd-4257,32'd-100,32'd-1596,32'd-453,32'd4228,32'd-5014,32'd2600,32'd-9833,32'd9506,32'd-4538,32'd-8354,32'd-6718,32'd-751,32'd-1618,32'd-5351,32'd7856,32'd8422,32'd76,32'd2819,32'd-7592,32'd301,32'd5239,32'd-1936,32'd-2846,32'd-4775,32'd-4108};
    Wx[23]='{32'd-684,32'd5375,32'd-1573,32'd-1748,32'd3486,32'd-496,32'd1864,32'd12,32'd-39,32'd-205,32'd5102,32'd-779,32'd1285,32'd-3767,32'd749,32'd6015,32'd2125,32'd552,32'd1271,32'd161,32'd-5444,32'd983,32'd-1196,32'd-1170,32'd-708,32'd1341,32'd-142,32'd-2673,32'd53,32'd8056,32'd-1313,32'd8178,32'd64,32'd-910,32'd-3671,32'd-447,32'd1704,32'd405,32'd1802,32'd3786,32'd-318,32'd4001,32'd202,32'd-844,32'd5688,32'd2604,32'd6875,32'd5483,32'd4169,32'd3166,32'd2778,32'd6811,32'd-1141,32'd132,32'd2296,32'd4531,32'd-7685,32'd-4902,32'd3027,32'd5727,32'd-5200,32'd-284,32'd3251,32'd-333,32'd8930,32'd74,32'd-1004,32'd4228,32'd646,32'd-1375,32'd-1068,32'd5439,32'd3630,32'd-812,32'd3054,32'd-229,32'd966,32'd-599,32'd3703,32'd-444,32'd1882,32'd4458,32'd-5566,32'd13701,32'd760,32'd897,32'd2856,32'd-3508,32'd1110,32'd-927,32'd6430,32'd-755,32'd-152,32'd2575,32'd2476,32'd2008,32'd3005,32'd379,32'd259,32'd5502,32'd5058,32'd-5224,32'd1511,32'd-8969,32'd-1469,32'd657,32'd5009,32'd-10507,32'd-2827,32'd134,32'd-9672,32'd-6284,32'd-8081,32'd-5415,32'd-7021,32'd-7148,32'd18671,32'd1918,32'd254,32'd636,32'd-2912,32'd1051,32'd-975,32'd-5541,32'd2695,32'd-3107,32'd1542,32'd1585,32'd4636,32'd2531,32'd4060,32'd-1324,32'd-2543,32'd-10117,32'd-463,32'd2409,32'd-774,32'd-172,32'd9526,32'd-4140,32'd-6484,32'd18623,32'd655,32'd-2734,32'd-3540,32'd12939,32'd-4689,32'd-7402,32'd3671,32'd3054,32'd-11630,32'd-13027,32'd3242,32'd13496,32'd-2052,32'd-3850,32'd-12880,32'd765,32'd-2076,32'd-4367,32'd-4487,32'd-12333,32'd-11738,32'd-4741,32'd-6464,32'd-1032,32'd1964,32'd-12988,32'd1633,32'd-2355,32'd12187,32'd-7968,32'd4545,32'd-16767,32'd1141,32'd3498,32'd-5688,32'd9560,32'd-6762,32'd4948,32'd6186,32'd1413,32'd-2023,32'd-729,32'd-671,32'd-4455,32'd-2126,32'd-6333,32'd4089,32'd-4702,32'd-3112,32'd-8320,32'd-2220,32'd2978,32'd-9809,32'd7500,32'd-2565,32'd-2186,32'd-5571,32'd15498,32'd-1151,32'd1907,32'd-553,32'd-3479,32'd-1271,32'd828,32'd-5649,32'd-1263,32'd6635,32'd-3405,32'd3898,32'd596,32'd-549,32'd-8950,32'd-4379,32'd-5449,32'd-5185,32'd-232,32'd-1782,32'd6269,32'd-3566,32'd-3493,32'd1252,32'd3725,32'd-370,32'd-5195,32'd-3645,32'd-2819,32'd2678,32'd-4846,32'd-1046,32'd217,32'd-7666,32'd-10605,32'd10878,32'd2305,32'd-67,32'd465,32'd-10087,32'd-559,32'd17,32'd-3125,32'd1501,32'd-1816,32'd-2260,32'd-3769,32'd9501,32'd-1962,32'd-1196,32'd2397,32'd6074,32'd-8979,32'd-2454,32'd861,32'd29,32'd-4667,32'd-1622,32'd1419,32'd-9199,32'd-3427,32'd-758,32'd9702,32'd3000,32'd-3330,32'd-16142,32'd421,32'd-2995,32'd11542,32'd873,32'd-1673,32'd-7036,32'd292,32'd-276,32'd484,32'd-1466,32'd4367,32'd-653,32'd3110,32'd-1541,32'd-2264,32'd3647,32'd6928,32'd5571,32'd4121,32'd-6918,32'd8354,32'd5551,32'd5620,32'd-832,32'd3376,32'd-3083,32'd1055,32'd2519,32'd2452,32'd4279,32'd844,32'd-6821,32'd-10029,32'd-1704,32'd2216,32'd2629,32'd-1450,32'd-3857,32'd1238,32'd-470,32'd1939,32'd-5024,32'd3872,32'd4992,32'd-4172,32'd-2709,32'd1840,32'd1932,32'd-12011,32'd2512,32'd-358,32'd-4475,32'd-5874,32'd-2841,32'd-2224,32'd-721,32'd-716,32'd-1624,32'd788,32'd3356,32'd-4672,32'd-6845,32'd-3417,32'd12304,32'd-4445,32'd-3193,32'd-1483,32'd-838,32'd-5390,32'd4357,32'd770,32'd-1723,32'd2106,32'd7861,32'd-1751,32'd-3337,32'd12568,32'd310,32'd-1733,32'd-1187,32'd106,32'd5019,32'd-4333,32'd2019,32'd-2165,32'd4343,32'd-4594,32'd4033,32'd-3601,32'd823,32'd-6333,32'd-585,32'd-11386,32'd478,32'd-751,32'd487,32'd2091,32'd9838,32'd4077,32'd406,32'd8774,32'd4621,32'd2489,32'd1014,32'd-9477,32'd-1677,32'd1654,32'd1968,32'd9990,32'd-3684,32'd3937,32'd6298,32'd-1480,32'd-786,32'd-3757,32'd528,32'd1529,32'd-2915,32'd7963,32'd-13701,32'd1998,32'd7055,32'd-2119,32'd2541,32'd692,32'd2612,32'd6240,32'd5688,32'd7597,32'd2758,32'd6669,32'd-343,32'd-2457,32'd-4211,32'd786};
    Wx[24]='{32'd-1484,32'd7475,32'd-4870,32'd-2083,32'd-2121,32'd445,32'd8271,32'd-3049,32'd-1505,32'd2729,32'd-5273,32'd-198,32'd-3674,32'd-223,32'd2736,32'd-5830,32'd-8168,32'd4262,32'd3903,32'd-591,32'd2142,32'd2929,32'd1445,32'd1431,32'd-552,32'd-933,32'd2580,32'd1934,32'd9687,32'd710,32'd1676,32'd3193,32'd683,32'd-1655,32'd-1196,32'd-864,32'd-4255,32'd-629,32'd-468,32'd1047,32'd2481,32'd5322,32'd1721,32'd370,32'd1923,32'd2966,32'd3493,32'd-2597,32'd-3049,32'd2181,32'd5546,32'd-1796,32'd864,32'd2335,32'd-1501,32'd3149,32'd-3508,32'd-2131,32'd2304,32'd378,32'd5180,32'd2949,32'd-235,32'd-1140,32'd-3937,32'd3071,32'd961,32'd-4982,32'd259,32'd2468,32'd1427,32'd4265,32'd-2841,32'd-1992,32'd-362,32'd-2103,32'd942,32'd-674,32'd941,32'd4060,32'd-3769,32'd1744,32'd-1043,32'd-4436,32'd-4846,32'd2541,32'd-3500,32'd-33,32'd-476,32'd-1801,32'd-5717,32'd-52,32'd736,32'd640,32'd2150,32'd-1444,32'd-303,32'd-906,32'd-1068,32'd-1550,32'd316,32'd17460,32'd8593,32'd12558,32'd8017,32'd-2883,32'd-10302,32'd17070,32'd-2247,32'd-89,32'd-13310,32'd-1503,32'd1287,32'd-8315,32'd-6025,32'd-9985,32'd122,32'd7626,32'd165,32'd-256,32'd235,32'd-6503,32'd-4216,32'd247,32'd5424,32'd-2426,32'd-2622,32'd-13144,32'd2934,32'd788,32'd-3344,32'd-2302,32'd9360,32'd1600,32'd-4650,32'd662,32'd3823,32'd-5068,32'd-2900,32'd-1834,32'd-3579,32'd7148,32'd4865,32'd2885,32'd3491,32'd-2214,32'd-2087,32'd-7993,32'd-1702,32'd806,32'd-2949,32'd11875,32'd-4445,32'd-12294,32'd6191,32'd-19179,32'd3916,32'd4611,32'd2491,32'd-127,32'd6298,32'd-3825,32'd8227,32'd-7363,32'd-5097,32'd314,32'd811,32'd-34335,32'd-1535,32'd4599,32'd12578,32'd-10556,32'd-69,32'd6333,32'd8315,32'd-24589,32'd13144,32'd-832,32'd-5332,32'd6250,32'd9887,32'd-2980,32'd-2462,32'd-9565,32'd-12578,32'd8115,32'd6166,32'd2229,32'd-4523,32'd-6181,32'd-1173,32'd-3750,32'd13437,32'd212,32'd13076,32'd-4565,32'd3256,32'd-7646,32'd1749,32'd-11240,32'd1699,32'd-10957,32'd-5009,32'd3112,32'd-461,32'd635,32'd6040,32'd-1503,32'd-5087,32'd2604,32'd-424,32'd-3632,32'd1719,32'd-2624,32'd-2008,32'd4584,32'd-2636,32'd-3615,32'd4975,32'd-511,32'd558,32'd2496,32'd102,32'd1311,32'd1816,32'd-4572,32'd1511,32'd254,32'd927,32'd-8251,32'd1989,32'd-2268,32'd-266,32'd3564,32'd-1346,32'd1400,32'd1030,32'd-488,32'd4912,32'd1396,32'd1932,32'd437,32'd-3046,32'd-5610,32'd-3774,32'd293,32'd-8569,32'd1506,32'd-1417,32'd1853,32'd2861,32'd-6918,32'd6000,32'd4904,32'd464,32'd-3139,32'd-4467,32'd1862,32'd-2077,32'd2854,32'd3117,32'd8012,32'd-1289,32'd9155,32'd955,32'd-3068,32'd4196,32'd-1810,32'd1577,32'd-1038,32'd-3740,32'd-571,32'd1203,32'd158,32'd1223,32'd4709,32'd11132,32'd-1575,32'd2263,32'd-2705,32'd-1015,32'd-6083,32'd-2209,32'd-102,32'd-5454,32'd-6,32'd-966,32'd-467,32'd3098,32'd-3696,32'd2301,32'd-4504,32'd-1917,32'd96,32'd4812,32'd3205,32'd-440,32'd2795,32'd4482,32'd-1308,32'd3156,32'd-6435,32'd-5922,32'd4831,32'd2492,32'd10761,32'd7055,32'd770,32'd-1640,32'd6093,32'd-11250,32'd-5024,32'd-869,32'd3803,32'd186,32'd-4521,32'd5288,32'd-721,32'd6235,32'd-4858,32'd6406,32'd5092,32'd-136,32'd-1730,32'd4138,32'd-8129,32'd8291,32'd472,32'd7915,32'd-5893,32'd-1630,32'd-3159,32'd-2147,32'd3271,32'd1795,32'd-1049,32'd-1558,32'd2790,32'd3999,32'd-3366,32'd3166,32'd133,32'd-4379,32'd-4399,32'd-47,32'd3193,32'd2900,32'd-5742,32'd-3354,32'd-398,32'd7802,32'd7866,32'd4418,32'd6127,32'd7939,32'd8364,32'd-4997,32'd-3771,32'd411,32'd8349,32'd-2800,32'd5112,32'd-6191,32'd2656,32'd3591,32'd635,32'd-1462,32'd-1634,32'd13955,32'd8149,32'd3234,32'd-2110,32'd3891,32'd-3771,32'd5458,32'd997,32'd3947,32'd-1041,32'd2237,32'd-20,32'd-697,32'd-7915,32'd-2995,32'd-10087,32'd-9174,32'd-825,32'd-3679,32'd-890,32'd-2475,32'd-2254,32'd2072,32'd3515,32'd-3366,32'd-7573,32'd-2897,32'd286,32'd245,32'd14199,32'd8759,32'd3850};
    Wx[25]='{32'd-964,32'd3039,32'd68,32'd4521,32'd-159,32'd-1945,32'd-216,32'd2147,32'd1508,32'd-5639,32'd-681,32'd618,32'd-541,32'd1530,32'd2521,32'd3051,32'd6782,32'd857,32'd1843,32'd-1031,32'd-1511,32'd647,32'd701,32'd-112,32'd1480,32'd-3037,32'd1525,32'd-1480,32'd3061,32'd-1334,32'd5263,32'd-8872,32'd-463,32'd-3754,32'd-2242,32'd-428,32'd566,32'd1580,32'd2127,32'd-3300,32'd1141,32'd939,32'd4035,32'd-4353,32'd2443,32'd-869,32'd2521,32'd5151,32'd3540,32'd4003,32'd4570,32'd326,32'd116,32'd667,32'd-307,32'd4575,32'd2895,32'd-3227,32'd3613,32'd-581,32'd-1348,32'd3657,32'd5771,32'd-1335,32'd581,32'd-1236,32'd-1065,32'd-7929,32'd-1195,32'd392,32'd-1535,32'd-3408,32'd2741,32'd2719,32'd-676,32'd548,32'd1346,32'd379,32'd4548,32'd-2088,32'd1660,32'd-5820,32'd121,32'd-4079,32'd1584,32'd-662,32'd2448,32'd-2025,32'd1497,32'd5761,32'd1857,32'd-5302,32'd7260,32'd-2305,32'd2524,32'd3632,32'd5874,32'd3664,32'd982,32'd-1921,32'd1724,32'd-8774,32'd-2199,32'd2078,32'd-9316,32'd-1832,32'd2988,32'd6079,32'd-1064,32'd7778,32'd4836,32'd-4802,32'd12011,32'd12412,32'd-6362,32'd7568,32'd3471,32'd531,32'd-2165,32'd-808,32'd1076,32'd4768,32'd473,32'd-3171,32'd2844,32'd4106,32'd168,32'd2148,32'd3994,32'd6791,32'd-550,32'd1602,32'd10439,32'd-3330,32'd-850,32'd-8012,32'd-8300,32'd-1962,32'd3000,32'd-6679,32'd4907,32'd8955,32'd4877,32'd1109,32'd-20253,32'd-378,32'd-3605,32'd-9609,32'd-2509,32'd2795,32'd-19365,32'd-4011,32'd-4787,32'd10595,32'd-1654,32'd3134,32'd3635,32'd412,32'd-901,32'd6679,32'd3471,32'd8408,32'd5058,32'd3679,32'd1844,32'd-3937,32'd4348,32'd18818,32'd-778,32'd1234,32'd1850,32'd9648,32'd3850,32'd-5493,32'd338,32'd5288,32'd12109,32'd-7607,32'd7026,32'd-11308,32'd-1444,32'd-10097,32'd1092,32'd4909,32'd-723,32'd59,32'd-488,32'd-8261,32'd-2612,32'd2326,32'd-4016,32'd-10898,32'd-1881,32'd969,32'd-2370,32'd7016,32'd4892,32'd-6191,32'd-623,32'd-7387,32'd-1860,32'd1776,32'd605,32'd-1435,32'd-3261,32'd57,32'd-1826,32'd-5292,32'd-4653,32'd-1342,32'd8349,32'd-2429,32'd-3608,32'd6723,32'd-6254,32'd1777,32'd7377,32'd467,32'd5507,32'd-735,32'd-587,32'd-106,32'd-1201,32'd-4531,32'd367,32'd-4028,32'd1472,32'd-912,32'd-6308,32'd2990,32'd4814,32'd-10839,32'd-13613,32'd-8676,32'd-4650,32'd-574,32'd-9091,32'd-3522,32'd-8784,32'd-888,32'd-4309,32'd-798,32'd-7949,32'd5424,32'd-2644,32'd-5102,32'd-9365,32'd-3166,32'd-219,32'd3193,32'd145,32'd-404,32'd273,32'd-1494,32'd-480,32'd-10468,32'd2180,32'd-6010,32'd-948,32'd2856,32'd195,32'd-3435,32'd-9663,32'd8188,32'd-11660,32'd-3706,32'd-5244,32'd-2102,32'd859,32'd-1314,32'd-6621,32'd2442,32'd4335,32'd3032,32'd-2912,32'd-8217,32'd-8642,32'd-6860,32'd-1112,32'd-769,32'd67,32'd505,32'd-2619,32'd3891,32'd1282,32'd-1064,32'd-1234,32'd-2032,32'd-792,32'd1881,32'd4201,32'd2519,32'd-4338,32'd-2071,32'd-5361,32'd-834,32'd-1822,32'd-621,32'd-8061,32'd-8793,32'd1256,32'd5878,32'd6455,32'd-1872,32'd1424,32'd-6245,32'd3251,32'd-10039,32'd-2973,32'd-6562,32'd11445,32'd5927,32'd5405,32'd-2546,32'd-8300,32'd-2983,32'd957,32'd16005,32'd713,32'd5996,32'd-5112,32'd4926,32'd2961,32'd-407,32'd3242,32'd4714,32'd1400,32'd-6748,32'd785,32'd5117,32'd6811,32'd-3730,32'd-11640,32'd-9799,32'd2418,32'd819,32'd-1044,32'd-4033,32'd-1024,32'd-141,32'd1395,32'd-2283,32'd3784,32'd1021,32'd2081,32'd-2332,32'd-8227,32'd466,32'd-2014,32'd7221,32'd-1308,32'd-3527,32'd6191,32'd4829,32'd4721,32'd-4587,32'd9926,32'd8437,32'd5776,32'd83,32'd-1489,32'd3071,32'd-1028,32'd1293,32'd-4477,32'd-11650,32'd-3493,32'd-5156,32'd-2731,32'd-1260,32'd4282,32'd-4072,32'd-397,32'd5917,32'd-132,32'd5112,32'd-3486,32'd7436,32'd5737,32'd-3881,32'd-94,32'd3305,32'd1214,32'd-8720,32'd-4128,32'd-506,32'd-3098,32'd-413,32'd3696,32'd4755,32'd6894,32'd16757,32'd1012,32'd-2476,32'd-1416,32'd-819,32'd5561,32'd-10273,32'd-6611,32'd1579};
    Wx[26]='{32'd-447,32'd-125,32'd1287,32'd2673,32'd-460,32'd-1406,32'd-3466,32'd-1964,32'd-1406,32'd-3203,32'd599,32'd881,32'd2563,32'd-1958,32'd2448,32'd4489,32'd-2915,32'd-5893,32'd2070,32'd3464,32'd3327,32'd1652,32'd-181,32'd1114,32'd-130,32'd3066,32'd12,32'd-1879,32'd-6059,32'd614,32'd-1425,32'd-1214,32'd4108,32'd-4165,32'd2683,32'd-1052,32'd-1212,32'd1614,32'd1379,32'd-4187,32'd758,32'd-3503,32'd-7836,32'd-2768,32'd5117,32'd-928,32'd7456,32'd1270,32'd-1084,32'd3713,32'd-5068,32'd-2047,32'd-123,32'd3500,32'd2021,32'd4438,32'd-2778,32'd2454,32'd-852,32'd-1763,32'd-2683,32'd-2060,32'd2817,32'd-3281,32'd2465,32'd-1016,32'd-393,32'd3127,32'd-1989,32'd1824,32'd4953,32'd3579,32'd4155,32'd-5185,32'd2360,32'd4924,32'd-2644,32'd593,32'd217,32'd-4831,32'd-1466,32'd2463,32'd438,32'd-5336,32'd2014,32'd-3635,32'd884,32'd-2768,32'd-1431,32'd2656,32'd-1010,32'd5112,32'd-313,32'd-1871,32'd25,32'd-1304,32'd-515,32'd-3012,32'd-6298,32'd989,32'd2946,32'd-10986,32'd2539,32'd-5527,32'd734,32'd-1929,32'd9995,32'd-7612,32'd-4709,32'd-2805,32'd2139,32'd4890,32'd-4333,32'd-5541,32'd2403,32'd-5307,32'd-2690,32'd6889,32'd-2751,32'd2897,32'd1510,32'd2427,32'd3449,32'd2176,32'd-2249,32'd-11953,32'd-11367,32'd3366,32'd-6738,32'd-7363,32'd362,32'd-1425,32'd-7885,32'd-1257,32'd1250,32'd4086,32'd-17,32'd2580,32'd-1271,32'd6933,32'd-5219,32'd-9272,32'd-11074,32'd-1510,32'd-1045,32'd940,32'd-14267,32'd-3701,32'd-1264,32'd-8525,32'd2469,32'd-23593,32'd-15,32'd3498,32'd3488,32'd-2980,32'd-3017,32'd-866,32'd10595,32'd3540,32'd-4946,32'd-7739,32'd-1416,32'd5151,32'd-5961,32'd-329,32'd-5986,32'd-4089,32'd-651,32'd3886,32'd2841,32'd13798,32'd357,32'd11787,32'd-988,32'd3098,32'd9350,32'd-10488,32'd3503,32'd-10107,32'd-8129,32'd-1887,32'd3205,32'd-22617,32'd919,32'd7280,32'd-1367,32'd-5468,32'd-3684,32'd-871,32'd-2570,32'd-4626,32'd1997,32'd-1815,32'd-2070,32'd-2504,32'd-4785,32'd2639,32'd-738,32'd-7060,32'd1040,32'd-1030,32'd-4001,32'd-1501,32'd189,32'd-478,32'd1586,32'd402,32'd-133,32'd-1899,32'd-1215,32'd1201,32'd1539,32'd-1089,32'd3508,32'd480,32'd3923,32'd5083,32'd7265,32'd219,32'd2288,32'd-16,32'd1365,32'd-2254,32'd-4648,32'd-8955,32'd-1323,32'd-2517,32'd4135,32'd-4729,32'd1188,32'd7104,32'd-256,32'd-10097,32'd4233,32'd3215,32'd-3876,32'd1614,32'd-5732,32'd4782,32'd1240,32'd4582,32'd-2349,32'd3852,32'd-3303,32'd796,32'd5234,32'd-1042,32'd1419,32'd-4641,32'd8330,32'd7641,32'd-831,32'd-3518,32'd-1470,32'd8505,32'd-1159,32'd-5048,32'd1917,32'd3894,32'd-2012,32'd-1654,32'd-7226,32'd-654,32'd-5571,32'd817,32'd-318,32'd-12333,32'd177,32'd4665,32'd-2375,32'd-3283,32'd-881,32'd4824,32'd146,32'd4194,32'd1140,32'd3891,32'd-2597,32'd-2719,32'd-1568,32'd3876,32'd-85,32'd874,32'd-1112,32'd2678,32'd2027,32'd3166,32'd2387,32'd-6079,32'd107,32'd-2968,32'd-1130,32'd-773,32'd-3984,32'd-3457,32'd1945,32'd6743,32'd-4941,32'd-265,32'd-1994,32'd3178,32'd277,32'd-56,32'd3549,32'd-4262,32'd7065,32'd-5395,32'd-4677,32'd-2658,32'd-3959,32'd-1099,32'd944,32'd2817,32'd-2496,32'd-3540,32'd-3715,32'd-3159,32'd6757,32'd244,32'd-677,32'd-1992,32'd-3061,32'd-3288,32'd2376,32'd1446,32'd-6748,32'd-8286,32'd5234,32'd2269,32'd424,32'd4785,32'd2293,32'd-5966,32'd-1140,32'd533,32'd-1451,32'd-427,32'd1855,32'd-640,32'd54,32'd2702,32'd-1617,32'd-2169,32'd-936,32'd-1192,32'd5747,32'd6547,32'd70,32'd835,32'd8652,32'd-1844,32'd-1374,32'd-2763,32'd-12226,32'd4011,32'd1845,32'd7695,32'd1754,32'd-5971,32'd1356,32'd-1661,32'd11435,32'd-6030,32'd-9521,32'd6538,32'd-6992,32'd126,32'd-10927,32'd-1033,32'd1273,32'd-6870,32'd-2391,32'd325,32'd1169,32'd1068,32'd8432,32'd1124,32'd752,32'd-8076,32'd-5131,32'd-863,32'd6435,32'd3400,32'd-1951,32'd5009,32'd1379,32'd3957,32'd4545,32'd11308,32'd-3251,32'd-16318,32'd-1971,32'd-6635,32'd-970,32'd-1040,32'd-2966,32'd1154,32'd-3164,32'd4870};
    Wx[27]='{32'd2622,32'd-3686,32'd-2746,32'd-317,32'd2895,32'd974,32'd-4682,32'd-2670,32'd5268,32'd5766,32'd-3461,32'd35,32'd516,32'd-5703,32'd4182,32'd-3767,32'd2188,32'd1459,32'd1358,32'd-172,32'd3620,32'd-1263,32'd-3537,32'd16,32'd-2406,32'd2410,32'd-2039,32'd2275,32'd-2526,32'd3942,32'd4479,32'd-4101,32'd-7177,32'd-5234,32'd4775,32'd-2188,32'd7543,32'd690,32'd-2397,32'd-4812,32'd-212,32'd-2727,32'd-421,32'd-3254,32'd-10224,32'd1916,32'd-6220,32'd589,32'd-2490,32'd-1794,32'd5620,32'd-3767,32'd-3806,32'd2902,32'd-2719,32'd-3115,32'd-1907,32'd2668,32'd-259,32'd312,32'd-490,32'd-500,32'd-6713,32'd-620,32'd-249,32'd-3454,32'd2103,32'd-11992,32'd746,32'd-3481,32'd-3320,32'd-328,32'd-383,32'd1002,32'd2092,32'd-2907,32'd-4609,32'd8105,32'd-5693,32'd-4709,32'd176,32'd-12548,32'd-5161,32'd-9589,32'd2097,32'd5810,32'd5107,32'd776,32'd366,32'd-2878,32'd1010,32'd-9262,32'd-1878,32'd-2039,32'd-7851,32'd1520,32'd206,32'd-5024,32'd32,32'd-1530,32'd1844,32'd-12734,32'd282,32'd6513,32'd4899,32'd207,32'd6240,32'd-7631,32'd1496,32'd-98,32'd2310,32'd-5268,32'd-9277,32'd7739,32'd6704,32'd-2692,32'd6225,32'd8881,32'd-2958,32'd1591,32'd2539,32'd5200,32'd14833,32'd778,32'd-3750,32'd381,32'd1938,32'd-6040,32'd3913,32'd-234,32'd1181,32'd-6416,32'd-125,32'd-1285,32'd3986,32'd-820,32'd4211,32'd-3229,32'd-1179,32'd-9179,32'd4941,32'd-23671,32'd-11972,32'd6787,32'd10664,32'd-4758,32'd-5043,32'd8027,32'd-1267,32'd9472,32'd4079,32'd-12705,32'd1447,32'd-1520,32'd6391,32'd5947,32'd6494,32'd-5078,32'd5986,32'd2536,32'd-2517,32'd9140,32'd-123,32'd3000,32'd12851,32'd1436,32'd2182,32'd-4772,32'd2268,32'd-3386,32'd-8085,32'd-5854,32'd-2890,32'd15117,32'd-1522,32'd-3686,32'd-7705,32'd-12558,32'd-6899,32'd6113,32'd1039,32'd14560,32'd4167,32'd7158,32'd3159,32'd-12626,32'd-463,32'd-3979,32'd3991,32'd-5834,32'd-4675,32'd6650,32'd-1727,32'd1155,32'd-1149,32'd-10693,32'd1650,32'd12089,32'd-8154,32'd5683,32'd226,32'd1103,32'd3149,32'd-2856,32'd3234,32'd1922,32'd10771,32'd-111,32'd334,32'd1213,32'd-8515,32'd3620,32'd-141,32'd-1958,32'd8461,32'd3718,32'd140,32'd-495,32'd-1227,32'd512,32'd4516,32'd333,32'd-2883,32'd-982,32'd-1896,32'd2824,32'd-5429,32'd3010,32'd399,32'd186,32'd-2832,32'd4929,32'd3913,32'd1036,32'd-1474,32'd1925,32'd-2802,32'd-2971,32'd-2565,32'd-2497,32'd1888,32'd-7207,32'd5229,32'd-1756,32'd3918,32'd-4719,32'd-1254,32'd2890,32'd-1556,32'd5727,32'd-3188,32'd184,32'd1170,32'd361,32'd-3283,32'd-15585,32'd5410,32'd2587,32'd-4340,32'd-9287,32'd-2661,32'd-5268,32'd-1795,32'd738,32'd-2152,32'd-780,32'd2641,32'd-2283,32'd-1597,32'd1165,32'd-1131,32'd-5585,32'd-1114,32'd-106,32'd2834,32'd-5507,32'd-4523,32'd408,32'd4482,32'd4365,32'd-2766,32'd-241,32'd838,32'd2371,32'd-3469,32'd-2856,32'd-2517,32'd-8798,32'd-5747,32'd-959,32'd1958,32'd5410,32'd1761,32'd-92,32'd-1032,32'd9794,32'd4965,32'd7221,32'd2543,32'd-1000,32'd-1356,32'd-6708,32'd-3813,32'd-2377,32'd-1061,32'd-3378,32'd6987,32'd-1228,32'd3193,32'd14218,32'd-7514,32'd2166,32'd-2175,32'd-4133,32'd9428,32'd-528,32'd-2709,32'd-2871,32'd2020,32'd5053,32'd-6689,32'd2152,32'd-386,32'd-1350,32'd6333,32'd603,32'd-5107,32'd7299,32'd-3149,32'd2282,32'd4780,32'd-8081,32'd2088,32'd-7519,32'd2435,32'd1522,32'd1102,32'd5424,32'd-4104,32'd-5683,32'd4030,32'd-2561,32'd9921,32'd-4597,32'd-1384,32'd-10039,32'd-1594,32'd7055,32'd-1494,32'd1997,32'd5693,32'd-3039,32'd-4667,32'd2922,32'd-3352,32'd4396,32'd2624,32'd-232,32'd2260,32'd4721,32'd2163,32'd-2685,32'd-680,32'd6816,32'd2812,32'd-1704,32'd-3769,32'd-2266,32'd14843,32'd-5893,32'd1989,32'd-9931,32'd-3090,32'd3391,32'd-3562,32'd-12246,32'd3203,32'd-3029,32'd6860,32'd-254,32'd-85,32'd-3908,32'd-4802,32'd-7832,32'd189,32'd-6000,32'd4914,32'd-6206,32'd1885,32'd-6865,32'd4960,32'd-1055,32'd-2963,32'd-7875,32'd-1337,32'd12832,32'd2558,32'd2866,32'd2812,32'd-3601};
    Wx[28]='{32'd2086,32'd1036,32'd-2094,32'd-2707,32'd987,32'd3969,32'd1832,32'd1342,32'd-116,32'd-928,32'd1945,32'd-1751,32'd2402,32'd6352,32'd-2712,32'd-734,32'd-286,32'd-184,32'd2054,32'd1049,32'd-158,32'd-3305,32'd259,32'd2220,32'd105,32'd238,32'd4360,32'd-842,32'd1280,32'd-1126,32'd2391,32'd7133,32'd-2486,32'd-3186,32'd-1207,32'd-4096,32'd4057,32'd-179,32'd-1663,32'd-1981,32'd2391,32'd-5200,32'd2600,32'd1273,32'd-103,32'd225,32'd-9462,32'd-1888,32'd-597,32'd784,32'd-5429,32'd-5585,32'd-2812,32'd549,32'd1748,32'd4375,32'd682,32'd-1973,32'd-6069,32'd-1870,32'd4653,32'd1379,32'd1166,32'd-7299,32'd-2980,32'd877,32'd-3830,32'd-7880,32'd2161,32'd3432,32'd1195,32'd-2254,32'd3737,32'd2780,32'd-3117,32'd2810,32'd-1831,32'd-1040,32'd-2396,32'd8081,32'd949,32'd-9184,32'd1610,32'd-4987,32'd2485,32'd-2963,32'd-2178,32'd-1468,32'd2507,32'd1004,32'd-3432,32'd-4111,32'd79,32'd-931,32'd3725,32'd-3078,32'd-457,32'd1568,32'd4743,32'd-1685,32'd-1496,32'd8974,32'd-2347,32'd-11748,32'd1395,32'd-1547,32'd6967,32'd6118,32'd-3669,32'd4287,32'd-8632,32'd-6899,32'd-1624,32'd-8100,32'd-8486,32'd-9990,32'd2607,32'd2929,32'd-780,32'd2705,32'd1531,32'd-2697,32'd-5727,32'd1788,32'd1418,32'd-7031,32'd-5366,32'd4243,32'd-808,32'd17402,32'd858,32'd12304,32'd12343,32'd-18066,32'd-4614,32'd-8051,32'd-4750,32'd3171,32'd5410,32'd2132,32'd-8188,32'd5380,32'd5556,32'd-8876,32'd206,32'd-2243,32'd1015,32'd-11718,32'd5380,32'd-11962,32'd1374,32'd-2949,32'd-8002,32'd12500,32'd-3115,32'd-10439,32'd-13505,32'd1789,32'd1636,32'd3618,32'd56,32'd6855,32'd3669,32'd1534,32'd-9174,32'd-2641,32'd7919,32'd10566,32'd-3166,32'd-1821,32'd9965,32'd762,32'd1545,32'd-14208,32'd-1921,32'd7456,32'd13437,32'd10996,32'd-8774,32'd-3942,32'd160,32'd7993,32'd12529,32'd-13964,32'd-2067,32'd5249,32'd2290,32'd1107,32'd-1412,32'd4313,32'd-494,32'd4057,32'd4890,32'd256,32'd-535,32'd1607,32'd-12880,32'd13222,32'd12460,32'd2432,32'd-2783,32'd-3544,32'd-1021,32'd5605,32'd-3273,32'd-285,32'd-865,32'd938,32'd-1909,32'd-5683,32'd-1722,32'd-1214,32'd-3127,32'd1351,32'd-3791,32'd1750,32'd1647,32'd5668,32'd4309,32'd-1090,32'd1530,32'd-2670,32'd-3166,32'd-304,32'd14,32'd-891,32'd-974,32'd-1166,32'd-8916,32'd2653,32'd3237,32'd-403,32'd-1973,32'd-729,32'd-6220,32'd3847,32'd-6635,32'd-4536,32'd4621,32'd3588,32'd-1267,32'd-7998,32'd126,32'd-2058,32'd4184,32'd-665,32'd-10166,32'd1190,32'd1168,32'd2707,32'd4572,32'd-7436,32'd-1965,32'd-1669,32'd702,32'd-1943,32'd1689,32'd-487,32'd-11210,32'd679,32'd-2387,32'd-5234,32'd4077,32'd-3432,32'd-6074,32'd1953,32'd-6362,32'd-8261,32'd3674,32'd-1130,32'd950,32'd221,32'd1560,32'd2619,32'd-2590,32'd-6474,32'd14980,32'd8623,32'd3781,32'd5581,32'd-7377,32'd2137,32'd2053,32'd-2136,32'd-5302,32'd380,32'd-1811,32'd1990,32'd5927,32'd-4379,32'd-1234,32'd-5126,32'd6865,32'd1129,32'd4704,32'd1774,32'd-1544,32'd2597,32'd-5239,32'd409,32'd1405,32'd-1668,32'd-4653,32'd8193,32'd209,32'd-9038,32'd-5854,32'd1304,32'd12001,32'd-12148,32'd9414,32'd1938,32'd1271,32'd5156,32'd-11367,32'd772,32'd-2526,32'd6923,32'd-2753,32'd1285,32'd-7583,32'd-1850,32'd-181,32'd2797,32'd-4038,32'd-2570,32'd-2492,32'd-1510,32'd13017,32'd728,32'd6347,32'd2416,32'd-252,32'd930,32'd-1387,32'd-4958,32'd2529,32'd-8500,32'd-2364,32'd1956,32'd788,32'd8359,32'd-3364,32'd2150,32'd3884,32'd5229,32'd-9003,32'd-4760,32'd-2919,32'd-4758,32'd2851,32'd-1400,32'd-1975,32'd5092,32'd6347,32'd1901,32'd7524,32'd-5439,32'd-8544,32'd3007,32'd-995,32'd1925,32'd-1788,32'd-4826,32'd-4479,32'd-2988,32'd-12236,32'd-3317,32'd-975,32'd-1008,32'd-6000,32'd-29,32'd374,32'd4311,32'd-2644,32'd-4677,32'd9902,32'd10449,32'd797,32'd2897,32'd-11425,32'd1226,32'd4077,32'd-140,32'd6943,32'd6962,32'd-211,32'd-281,32'd7998,32'd17275,32'd-6113,32'd-1662,32'd2829,32'd1409,32'd121,32'd-4548,32'd-3977,32'd1708,32'd1178,32'd4597};
    Wx[29]='{32'd863,32'd-5468,32'd-3239,32'd-3564,32'd1238,32'd60,32'd-1130,32'd-3410,32'd-447,32'd1319,32'd2951,32'd-497,32'd-2934,32'd-7202,32'd-5175,32'd-12304,32'd-6708,32'd-343,32'd-195,32'd-2558,32'd-192,32'd-2963,32'd-4753,32'd-3334,32'd-664,32'd-2250,32'd-1973,32'd602,32'd-1166,32'd889,32'd1912,32'd-8427,32'd-626,32'd-7050,32'd-1331,32'd-1414,32'd-694,32'd-919,32'd-2724,32'd-3820,32'd-3847,32'd-2041,32'd-5234,32'd-4907,32'd-3000,32'd-2327,32'd-9541,32'd-6923,32'd-2827,32'd-2324,32'd-5322,32'd-4636,32'd6230,32'd-4628,32'd-3886,32'd-150,32'd-1049,32'd-2675,32'd-2188,32'd5444,32'd-2529,32'd-143,32'd-2727,32'd-7783,32'd-7026,32'd78,32'd950,32'd-6376,32'd-820,32'd597,32'd-4924,32'd-4909,32'd-2470,32'd651,32'd2072,32'd-5332,32'd-1174,32'd-723,32'd-4812,32'd4145,32'd1144,32'd-5556,32'd-1932,32'd-4445,32'd-231,32'd-831,32'd-2254,32'd-210,32'd-159,32'd-1127,32'd-741,32'd-5190,32'd-946,32'd-2502,32'd-3679,32'd-1429,32'd-2734,32'd1691,32'd-2583,32'd-8720,32'd446,32'd24902,32'd1676,32'd929,32'd2252,32'd1398,32'd-5805,32'd-123,32'd-1793,32'd-7182,32'd-1989,32'd476,32'd-1391,32'd4357,32'd-7075,32'd-10585,32'd5034,32'd2636,32'd-4536,32'd-3850,32'd-1056,32'd-55,32'd5429,32'd-10029,32'd3505,32'd2893,32'd8505,32'd-948,32'd4064,32'd-3439,32'd596,32'd8911,32'd-5742,32'd12070,32'd-608,32'd7241,32'd-202,32'd2008,32'd-119,32'd-9545,32'd3635,32'd3835,32'd1287,32'd9467,32'd721,32'd-1621,32'd-1260,32'd7158,32'd-1757,32'd4836,32'd5776,32'd-15498,32'd-52,32'd-2464,32'd3671,32'd10205,32'd2685,32'd-261,32'd-3942,32'd1451,32'd-2139,32'd-6362,32'd-6440,32'd-8598,32'd3762,32'd-834,32'd-3107,32'd293,32'd3728,32'd3540,32'd3005,32'd-4897,32'd3581,32'd-8720,32'd-977,32'd3195,32'd-10351,32'd17587,32'd2541,32'd-3027,32'd5805,32'd4655,32'd-1097,32'd12363,32'd-1139,32'd-8339,32'd441,32'd1262,32'd-1508,32'd309,32'd-2805,32'd26445,32'd-51,32'd-2493,32'd-9340,32'd-4953,32'd8496,32'd9321,32'd2917,32'd13457,32'd2241,32'd-5351,32'd-1557,32'd-847,32'd3886,32'd2083,32'd438,32'd-2683,32'd273,32'd-1392,32'd893,32'd-1854,32'd764,32'd-3898,32'd3833,32'd2841,32'd-4685,32'd-3642,32'd5649,32'd3342,32'd207,32'd-4096,32'd-491,32'd3137,32'd1666,32'd-3659,32'd2978,32'd2017,32'd-1541,32'd-1578,32'd1534,32'd-1001,32'd-3688,32'd-1785,32'd4548,32'd-28,32'd8515,32'd2534,32'd-10839,32'd2330,32'd3452,32'd5234,32'd2083,32'd-3610,32'd4018,32'd-4904,32'd8505,32'd339,32'd-3625,32'd2666,32'd-5097,32'd-1922,32'd5668,32'd6875,32'd-4140,32'd-4399,32'd-3801,32'd1663,32'd-7666,32'd-6044,32'd-4042,32'd-1682,32'd6430,32'd-1061,32'd-2320,32'd-2237,32'd-670,32'd3254,32'd-3081,32'd908,32'd-3007,32'd-6708,32'd-4335,32'd-8833,32'd788,32'd1141,32'd1477,32'd1552,32'd1254,32'd-1759,32'd-942,32'd-7045,32'd4687,32'd861,32'd945,32'd-7104,32'd-853,32'd3046,32'd7177,32'd1838,32'd2807,32'd-513,32'd-667,32'd-3510,32'd-68,32'd-5024,32'd-5903,32'd-2224,32'd4404,32'd-2861,32'd3671,32'd-69,32'd4084,32'd164,32'd-783,32'd16650,32'd-348,32'd-1827,32'd-4089,32'd-4721,32'd-1535,32'd-263,32'd-5058,32'd-4575,32'd-1591,32'd-4062,32'd-5292,32'd-3867,32'd11953,32'd-523,32'd283,32'd-2030,32'd-1802,32'd653,32'd3127,32'd-7314,32'd2094,32'd3911,32'd-6181,32'd-6093,32'd-708,32'd-5273,32'd1986,32'd-574,32'd-4130,32'd1799,32'd-3889,32'd7294,32'd-10585,32'd-5541,32'd891,32'd-6152,32'd-4113,32'd-1302,32'd-5478,32'd-11259,32'd-507,32'd-9106,32'd-2243,32'd1983,32'd-2463,32'd-5556,32'd6132,32'd-795,32'd-2204,32'd1506,32'd-2705,32'd-6997,32'd-855,32'd-6660,32'd-180,32'd-428,32'd378,32'd242,32'd-817,32'd5200,32'd5761,32'd1044,32'd3176,32'd5493,32'd3576,32'd-13369,32'd-130,32'd-4567,32'd1528,32'd-2165,32'd-2028,32'd-3088,32'd-1307,32'd2342,32'd-3208,32'd-2114,32'd-7495,32'd-2551,32'd-3945,32'd-10166,32'd-563,32'd-3022,32'd-7563,32'd-5576,32'd7055,32'd-1975,32'd-94,32'd-12675,32'd-11962,32'd-2678,32'd9428,32'd-1040,32'd5253,32'd-6601};
    Wx[30]='{32'd2231,32'd-14150,32'd-1365,32'd2551,32'd-953,32'd320,32'd5644,32'd-5390,32'd1663,32'd433,32'd276,32'd-659,32'd454,32'd-2783,32'd-4028,32'd-7587,32'd2351,32'd3859,32'd292,32'd356,32'd1733,32'd531,32'd-1813,32'd-3845,32'd-175,32'd-466,32'd1402,32'd398,32'd3369,32'd-1240,32'd-816,32'd-572,32'd-946,32'd-4482,32'd2114,32'd1503,32'd1212,32'd-197,32'd-318,32'd1303,32'd1251,32'd-2399,32'd-7221,32'd-4746,32'd3173,32'd3640,32'd-5937,32'd1196,32'd2034,32'd-62,32'd-3601,32'd469,32'd-3342,32'd-1951,32'd-3527,32'd-3806,32'd-1790,32'd2464,32'd-1335,32'd824,32'd-1772,32'd6977,32'd1231,32'd2539,32'd-1074,32'd-2449,32'd2369,32'd664,32'd1047,32'd2734,32'd184,32'd-2016,32'd-5424,32'd-584,32'd1877,32'd309,32'd-1146,32'd-2370,32'd-2548,32'd-1203,32'd2088,32'd-3388,32'd2172,32'd-166,32'd3027,32'd823,32'd-1441,32'd-3818,32'd1572,32'd-3112,32'd-348,32'd-3618,32'd77,32'd730,32'd-6313,32'd2719,32'd-2100,32'd3620,32'd-6635,32'd-1765,32'd-1513,32'd-137,32'd2315,32'd-4682,32'd2224,32'd-1311,32'd256,32'd-11464,32'd8750,32'd959,32'd-4265,32'd1846,32'd-2604,32'd4785,32'd-728,32'd3266,32'd20019,32'd-7114,32'd-1779,32'd-2766,32'd1745,32'd1271,32'd-533,32'd-1600,32'd-3947,32'd-8144,32'd6484,32'd3833,32'd-460,32'd-6123,32'd3659,32'd-5336,32'd-3549,32'd-748,32'd4882,32'd1546,32'd3779,32'd-3171,32'd-3154,32'd5268,32'd598,32'd-10849,32'd-518,32'd-1258,32'd4113,32'd-5166,32'd928,32'd-2283,32'd3623,32'd-1831,32'd-3759,32'd-2644,32'd5722,32'd-2597,32'd2858,32'd8466,32'd-1016,32'd-39,32'd4670,32'd545,32'd1608,32'd-4528,32'd-3259,32'd1109,32'd9365,32'd-139,32'd-1470,32'd6196,32'd-3095,32'd-68,32'd-13974,32'd-5253,32'd-3486,32'd3698,32'd-618,32'd-7299,32'd-6704,32'd217,32'd-2841,32'd-7543,32'd652,32'd-6977,32'd-186,32'd7832,32'd6235,32'd2303,32'd-1923,32'd-267,32'd-725,32'd-3488,32'd2739,32'd-1901,32'd1994,32'd573,32'd1374,32'd2457,32'd2683,32'd531,32'd-3759,32'd2958,32'd1781,32'd15468,32'd-1172,32'd27,32'd3842,32'd579,32'd1958,32'd-4499,32'd-1144,32'd2961,32'd182,32'd483,32'd383,32'd3583,32'd-1251,32'd-2624,32'd6987,32'd-179,32'd1176,32'd-1539,32'd-1445,32'd-1234,32'd882,32'd-2006,32'd1494,32'd1640,32'd-582,32'd-381,32'd10029,32'd-5610,32'd-6176,32'd2403,32'd737,32'd6284,32'd-3586,32'd-6870,32'd-4914,32'd2106,32'd850,32'd2246,32'd7041,32'd4814,32'd4650,32'd2429,32'd182,32'd7441,32'd1749,32'd-200,32'd573,32'd-629,32'd4384,32'd8618,32'd1439,32'd3696,32'd-3994,32'd-1988,32'd-1199,32'd158,32'd4711,32'd-5805,32'd173,32'd4035,32'd-729,32'd2919,32'd3813,32'd-2371,32'd5937,32'd4589,32'd-1870,32'd823,32'd1071,32'd-1791,32'd805,32'd3291,32'd2161,32'd1206,32'd640,32'd6040,32'd-1464,32'd-3452,32'd2932,32'd1678,32'd-1860,32'd-4077,32'd-2298,32'd-1636,32'd1152,32'd2592,32'd-902,32'd-697,32'd8,32'd6250,32'd-4697,32'd921,32'd3049,32'd5834,32'd6523,32'd40,32'd3237,32'd431,32'd2919,32'd13164,32'd6206,32'd-466,32'd1781,32'd5175,32'd6914,32'd-5170,32'd-5932,32'd-2670,32'd-8315,32'd322,32'd124,32'd5371,32'd-7797,32'd-7685,32'd8500,32'd4140,32'd-4338,32'd839,32'd3508,32'd668,32'd-5537,32'd526,32'd520,32'd916,32'd-136,32'd1342,32'd13398,32'd-290,32'd-2841,32'd2009,32'd-4042,32'd4460,32'd-10898,32'd-3188,32'd107,32'd-219,32'd4345,32'd3481,32'd3742,32'd9765,32'd3510,32'd-658,32'd1004,32'd-2022,32'd2543,32'd6342,32'd-3872,32'd3015,32'd886,32'd-5029,32'd5078,32'd1518,32'd-4201,32'd-3203,32'd-5200,32'd14023,32'd1718,32'd-3525,32'd3588,32'd4003,32'd-656,32'd4189,32'd190,32'd1872,32'd6396,32'd2907,32'd3913,32'd8876,32'd2558,32'd5385,32'd-249,32'd-2592,32'd-1881,32'd5122,32'd4221,32'd2807,32'd-4536,32'd-3559,32'd8803,32'd2250,32'd-653,32'd5839,32'd-5141,32'd8286,32'd209,32'd-2436,32'd3164,32'd4926,32'd-4,32'd-523,32'd-3645,32'd9594,32'd1058,32'd7548,32'd10166,32'd-299,32'd230,32'd5102};
    Wx[31]='{32'd2614,32'd3015,32'd-81,32'd456,32'd-994,32'd-2834,32'd232,32'd5268,32'd469,32'd2296,32'd3713,32'd738,32'd1759,32'd6352,32'd-1688,32'd3247,32'd4172,32'd2902,32'd3249,32'd511,32'd-1168,32'd343,32'd-1514,32'd-1536,32'd3403,32'd-148,32'd38,32'd2298,32'd2888,32'd-3828,32'd3078,32'd2376,32'd4829,32'd1922,32'd3923,32'd-403,32'd-1198,32'd-2841,32'd-1346,32'd-192,32'd509,32'd-2207,32'd-815,32'd526,32'd-7729,32'd6333,32'd5961,32'd-504,32'd-1165,32'd656,32'd-4487,32'd3730,32'd-7353,32'd-53,32'd-8281,32'd-5766,32'd245,32'd-5517,32'd-2437,32'd836,32'd4045,32'd3007,32'd-36,32'd-263,32'd7968,32'd2491,32'd2215,32'd2281,32'd-2841,32'd-74,32'd-3833,32'd312,32'd2597,32'd-4599,32'd886,32'd-1232,32'd-344,32'd2484,32'd-3205,32'd-607,32'd2705,32'd-523,32'd1446,32'd-1047,32'd-889,32'd952,32'd-4318,32'd-5161,32'd-983,32'd-265,32'd3676,32'd-6987,32'd1156,32'd-2636,32'd7412,32'd7495,32'd-991,32'd-4265,32'd4433,32'd2949,32'd-988,32'd-7597,32'd-3601,32'd-7167,32'd712,32'd3486,32'd4440,32'd704,32'd-1608,32'd1630,32'd-14179,32'd6391,32'd11328,32'd3151,32'd2487,32'd3962,32'd141,32'd3466,32'd-1545,32'd-4550,32'd-4953,32'd-3452,32'd2792,32'd2700,32'd2604,32'd1430,32'd-7138,32'd-3054,32'd2440,32'd7583,32'd-7695,32'd-13115,32'd4174,32'd10605,32'd6787,32'd5483,32'd4909,32'd-1549,32'd-9355,32'd3874,32'd2257,32'd-1584,32'd-1717,32'd6997,32'd2653,32'd7363,32'd958,32'd-1311,32'd-2159,32'd1330,32'd12597,32'd13730,32'd-19257,32'd7617,32'd6416,32'd9331,32'd4467,32'd2648,32'd-3129,32'd53,32'd3359,32'd-3388,32'd-5815,32'd3686,32'd-1572,32'd3034,32'd-4655,32'd-5507,32'd4814,32'd3513,32'd2497,32'd-10429,32'd-8823,32'd-7192,32'd4252,32'd360,32'd11464,32'd-17402,32'd15224,32'd-60,32'd6835,32'd5444,32'd5341,32'd11005,32'd-632,32'd3498,32'd2194,32'd-19785,32'd-220,32'd-9038,32'd-8061,32'd6157,32'd8374,32'd1502,32'd1834,32'd7182,32'd4042,32'd-3750,32'd2597,32'd1959,32'd1997,32'd-6318,32'd5278,32'd6440,32'd1915,32'd-1102,32'd3430,32'd8715,32'd734,32'd3610,32'd4680,32'd1782,32'd2478,32'd-4897,32'd-991,32'd2001,32'd-2211,32'd-78,32'd3420,32'd1300,32'd-124,32'd2274,32'd-2145,32'd4968,32'd3398,32'd-3840,32'd1827,32'd593,32'd1181,32'd7973,32'd-3681,32'd-8110,32'd-3808,32'd1888,32'd-3376,32'd7949,32'd993,32'd-2241,32'd1059,32'd1206,32'd-362,32'd-1168,32'd-2023,32'd6293,32'd4150,32'd2176,32'd-7661,32'd916,32'd-1654,32'd5917,32'd12460,32'd-3112,32'd-416,32'd3845,32'd-562,32'd221,32'd-1079,32'd-5380,32'd11376,32'd-3530,32'd2653,32'd9384,32'd1150,32'd-1420,32'd-4541,32'd2019,32'd8725,32'd-7661,32'd-2365,32'd-1888,32'd-1378,32'd-1032,32'd401,32'd9077,32'd1052,32'd4382,32'd8164,32'd11542,32'd1641,32'd-6074,32'd2147,32'd-16396,32'd-1657,32'd-4157,32'd-4104,32'd-1613,32'd-77,32'd1276,32'd97,32'd-3459,32'd7910,32'd2386,32'd1245,32'd-2910,32'd-11357,32'd3442,32'd5366,32'd4692,32'd838,32'd-453,32'd1766,32'd-11943,32'd4719,32'd-106,32'd3078,32'd-4299,32'd-5439,32'd3862,32'd3454,32'd11650,32'd-2467,32'd895,32'd1112,32'd134,32'd-2597,32'd488,32'd745,32'd-2897,32'd4221,32'd7265,32'd2741,32'd1674,32'd-3281,32'd1236,32'd3085,32'd-555,32'd4819,32'd994,32'd-1800,32'd-550,32'd-4750,32'd-5556,32'd-229,32'd6450,32'd-20,32'd3601,32'd-2722,32'd1390,32'd-960,32'd3774,32'd2998,32'd-2592,32'd-9702,32'd-1314,32'd-7358,32'd8535,32'd7631,32'd-68,32'd-4919,32'd509,32'd9106,32'd1496,32'd-8676,32'd-6411,32'd119,32'd-717,32'd1271,32'd3833,32'd3547,32'd-6010,32'd2088,32'd3959,32'd7617,32'd-4816,32'd205,32'd693,32'd10976,32'd-3925,32'd2624,32'd773,32'd-1240,32'd5000,32'd-2208,32'd556,32'd14140,32'd11855,32'd-7250,32'd770,32'd-7685,32'd-1243,32'd4663,32'd-7412,32'd5244,32'd-3732,32'd5849,32'd2788,32'd-386,32'd-8457,32'd623,32'd-4948,32'd11074,32'd-5151,32'd-1376,32'd-1892,32'd-5366,32'd1143,32'd-273,32'd3645,32'd3776,32'd4074};
    Wx[32]='{32'd968,32'd1072,32'd-785,32'd4270,32'd-2056,32'd997,32'd-444,32'd1931,32'd-1044,32'd1503,32'd-11259,32'd-1184,32'd-1012,32'd-2600,32'd701,32'd-1490,32'd2780,32'd-6284,32'd-289,32'd1439,32'd2452,32'd2761,32'd3476,32'd805,32'd2790,32'd-4467,32'd1064,32'd-476,32'd-123,32'd-430,32'd-737,32'd629,32'd879,32'd-1854,32'd378,32'd-841,32'd-1423,32'd916,32'd717,32'd2385,32'd-186,32'd-17,32'd-7778,32'd4003,32'd-6118,32'd-27,32'd10947,32'd-4370,32'd-3212,32'd-4584,32'd1590,32'd3276,32'd1623,32'd-1867,32'd3149,32'd-365,32'd-1564,32'd784,32'd-1846,32'd1652,32'd4870,32'd781,32'd6166,32'd4223,32'd-4619,32'd440,32'd-72,32'd-3835,32'd1348,32'd-1944,32'd-1428,32'd2265,32'd-115,32'd-2871,32'd2457,32'd-1752,32'd-3208,32'd-1081,32'd1418,32'd1534,32'd134,32'd4599,32'd1949,32'd-2145,32'd1702,32'd3193,32'd433,32'd5922,32'd-3491,32'd-261,32'd2836,32'd-1643,32'd-753,32'd-572,32'd5107,32'd2663,32'd-495,32'd-9223,32'd795,32'd267,32'd-791,32'd-10429,32'd-1134,32'd20,32'd2135,32'd-2467,32'd-4875,32'd5058,32'd-1018,32'd-1359,32'd979,32'd4890,32'd-946,32'd-3808,32'd5087,32'd-3300,32'd-22773,32'd6201,32'd357,32'd4707,32'd3037,32'd1109,32'd-58,32'd-791,32'd1955,32'd-3493,32'd-6298,32'd-4108,32'd12070,32'd7592,32'd1306,32'd10283,32'd-186,32'd-5014,32'd895,32'd-1616,32'd-3359,32'd600,32'd-2539,32'd-1271,32'd5869,32'd3862,32'd3620,32'd1765,32'd11376,32'd-4047,32'd-14179,32'd-305,32'd5717,32'd5249,32'd866,32'd4497,32'd7119,32'd2770,32'd1091,32'd3984,32'd2766,32'd2476,32'd-4079,32'd445,32'd5424,32'd-151,32'd7504,32'd-986,32'd-11464,32'd-4802,32'd717,32'd-8344,32'd-437,32'd-1130,32'd4909,32'd7636,32'd1246,32'd2944,32'd6474,32'd-5590,32'd3830,32'd6166,32'd-12636,32'd-1296,32'd-731,32'd9960,32'd8842,32'd-1188,32'd6538,32'd-3803,32'd-1387,32'd8256,32'd3134,32'd-3854,32'd488,32'd-2827,32'd2088,32'd-4194,32'd6083,32'd991,32'd-656,32'd-11250,32'd-7158,32'd-9052,32'd-2529,32'd-7617,32'd-1068,32'd-824,32'd-3139,32'd1586,32'd9501,32'd-4677,32'd2814,32'd-1229,32'd5981,32'd-1322,32'd3095,32'd-6123,32'd4189,32'd-3544,32'd6040,32'd-1951,32'd1291,32'd-727,32'd-321,32'd-2403,32'd2296,32'd-1336,32'd6474,32'd1193,32'd-4155,32'd-1614,32'd-7250,32'd7514,32'd661,32'd-1071,32'd-1453,32'd4255,32'd-541,32'd3349,32'd0,32'd2592,32'd1457,32'd-1210,32'd-3891,32'd1575,32'd6855,32'd5581,32'd4799,32'd-676,32'd-6127,32'd-3723,32'd5058,32'd740,32'd-611,32'd1403,32'd5786,32'd7758,32'd-1693,32'd-4750,32'd6811,32'd-1158,32'd-934,32'd-3217,32'd5087,32'd852,32'd7978,32'd3276,32'd3786,32'd4526,32'd1761,32'd7255,32'd-1122,32'd-922,32'd4895,32'd2039,32'd-1986,32'd6440,32'd1430,32'd-3657,32'd2049,32'd820,32'd-709,32'd13,32'd2277,32'd0,32'd1328,32'd6367,32'd93,32'd-1789,32'd2766,32'd-3850,32'd5590,32'd-904,32'd3898,32'd2248,32'd-1411,32'd3288,32'd5429,32'd-201,32'd5703,32'd-3747,32'd333,32'd176,32'd-2863,32'd-8222,32'd-7578,32'd-5727,32'd2702,32'd289,32'd5317,32'd-174,32'd-805,32'd7988,32'd417,32'd-4936,32'd5180,32'd-1567,32'd-2695,32'd1079,32'd716,32'd-7524,32'd291,32'd2160,32'd1633,32'd2282,32'd-1436,32'd-396,32'd3115,32'd-6406,32'd6162,32'd-2766,32'd-5375,32'd757,32'd-3581,32'd439,32'd-1870,32'd-1291,32'd-1386,32'd4882,32'd2232,32'd6606,32'd-4519,32'd-4899,32'd-3908,32'd-1223,32'd1134,32'd-3208,32'd-5009,32'd773,32'd6098,32'd885,32'd-2802,32'd-2832,32'd-4460,32'd4064,32'd5869,32'd839,32'd6333,32'd2498,32'd-1574,32'd3205,32'd288,32'd1520,32'd-3459,32'd2539,32'd90,32'd-5468,32'd-3251,32'd3854,32'd4868,32'd2983,32'd7172,32'd-10185,32'd6303,32'd-1649,32'd-4057,32'd1409,32'd5214,32'd-3195,32'd-1502,32'd-264,32'd-524,32'd472,32'd7104,32'd-2595,32'd9311,32'd5683,32'd4355,32'd2709,32'd2080,32'd-1394,32'd2988,32'd2668,32'd6694,32'd-10117,32'd-1763,32'd-7553,32'd4926,32'd4819,32'd6542,32'd1191,32'd301,32'd-1662};
    Wx[33]='{32'd687,32'd-2313,32'd653,32'd-1684,32'd-538,32'd908,32'd7,32'd-1911,32'd-5532,32'd-2407,32'd-908,32'd-2949,32'd1148,32'd-2402,32'd-8837,32'd9653,32'd3964,32'd-6635,32'd-376,32'd2349,32'd-1147,32'd-1293,32'd-1322,32'd-1771,32'd1184,32'd994,32'd-1931,32'd2220,32'd3164,32'd586,32'd632,32'd1448,32'd-1627,32'd3269,32'd-2519,32'd536,32'd2900,32'd-1213,32'd-2897,32'd-5517,32'd1589,32'd5439,32'd7749,32'd499,32'd2059,32'd5771,32'd1408,32'd190,32'd-3798,32'd1621,32'd9975,32'd2592,32'd3383,32'd4099,32'd4897,32'd7231,32'd-2382,32'd2042,32'd-4023,32'd5014,32'd3513,32'd5283,32'd-1903,32'd885,32'd2427,32'd1341,32'd-3730,32'd5449,32'd-2924,32'd-3728,32'd-28,32'd1275,32'd996,32'd-1101,32'd2309,32'd-7656,32'd-3852,32'd-3691,32'd2160,32'd-3928,32'd-2393,32'd76,32'd3181,32'd-10009,32'd-2144,32'd8789,32'd-406,32'd1104,32'd5048,32'd-73,32'd-5468,32'd-1428,32'd850,32'd1898,32'd-2038,32'd-377,32'd5859,32'd-8349,32'd1666,32'd-270,32'd-5473,32'd-2373,32'd-523,32'd-6777,32'd3811,32'd-1177,32'd-7050,32'd-4592,32'd-2805,32'd6542,32'd3562,32'd-5620,32'd10869,32'd-10351,32'd2475,32'd-1993,32'd-2265,32'd10048,32'd4104,32'd1337,32'd567,32'd9902,32'd-11435,32'd1573,32'd225,32'd382,32'd-2514,32'd-6787,32'd-3750,32'd-107,32'd3024,32'd-17832,32'd-6494,32'd2069,32'd-7841,32'd-2470,32'd-1848,32'd-5585,32'd-4084,32'd-9926,32'd3884,32'd-5380,32'd7138,32'd-673,32'd-19169,32'd-17617,32'd-3493,32'd10195,32'd-11337,32'd4196,32'd9755,32'd-11113,32'd-5771,32'd1365,32'd1209,32'd-11103,32'd-442,32'd310,32'd-1843,32'd-5395,32'd-737,32'd8115,32'd-2082,32'd4216,32'd3366,32'd-1931,32'd-2790,32'd-1859,32'd1412,32'd-164,32'd8588,32'd1489,32'd-1735,32'd5385,32'd-430,32'd-8305,32'd-12910,32'd12929,32'd6953,32'd-863,32'd-2958,32'd16220,32'd1517,32'd-12666,32'd-1688,32'd20878,32'd-96,32'd8686,32'd44,32'd-2305,32'd892,32'd5932,32'd-7324,32'd-448,32'd-4826,32'd-2941,32'd5834,32'd-12236,32'd8076,32'd-9121,32'd-4418,32'd-5214,32'd-1420,32'd2222,32'd3798,32'd751,32'd1254,32'd-122,32'd-353,32'd-2075,32'd-2666,32'd-888,32'd-1387,32'd-4162,32'd-14638,32'd-6079,32'd-5332,32'd-4418,32'd-3571,32'd570,32'd-1635,32'd-833,32'd3540,32'd-499,32'd-6264,32'd-6025,32'd-11953,32'd1011,32'd-2292,32'd4558,32'd4362,32'd-5751,32'd-267,32'd-10292,32'd-4243,32'd612,32'd-7680,32'd-4040,32'd591,32'd-991,32'd-3481,32'd2592,32'd2595,32'd-2717,32'd-1184,32'd-4721,32'd5625,32'd5190,32'd4414,32'd70,32'd-6074,32'd-2736,32'd-304,32'd-1187,32'd5913,32'd-5522,32'd2668,32'd-5117,32'd5742,32'd-1211,32'd8007,32'd-3222,32'd-2183,32'd-198,32'd-2445,32'd-7587,32'd-5395,32'd-4794,32'd2249,32'd-2883,32'd-601,32'd-1466,32'd-2142,32'd2927,32'd1206,32'd3703,32'd98,32'd-6708,32'd382,32'd-1400,32'd-4946,32'd4851,32'd-4870,32'd1674,32'd-3515,32'd-5253,32'd-5312,32'd-2990,32'd5249,32'd-567,32'd8413,32'd-1018,32'd3537,32'd-1781,32'd-397,32'd-4382,32'd2509,32'd-238,32'd-2678,32'd-3110,32'd-4011,32'd-941,32'd-8261,32'd-4787,32'd2294,32'd241,32'd2442,32'd6181,32'd-7441,32'd-1650,32'd-449,32'd1571,32'd699,32'd-4895,32'd-15625,32'd56,32'd-4353,32'd-13398,32'd3354,32'd-2222,32'd-3337,32'd-702,32'd3603,32'd-3271,32'd-6181,32'd-2976,32'd-6875,32'd-133,32'd-4074,32'd6430,32'd4001,32'd-184,32'd3625,32'd-8007,32'd-1300,32'd-1557,32'd-5253,32'd4975,32'd-4697,32'd-4270,32'd-3552,32'd3325,32'd4086,32'd2758,32'd-129,32'd-537,32'd2595,32'd9218,32'd-5029,32'd1624,32'd-3244,32'd-1915,32'd-1186,32'd908,32'd-87,32'd-6113,32'd-1033,32'd5224,32'd-6069,32'd-3608,32'd3315,32'd1740,32'd-3518,32'd421,32'd-2531,32'd-16083,32'd-3471,32'd-6948,32'd834,32'd-4152,32'd1118,32'd1920,32'd-2086,32'd-12753,32'd-2731,32'd2467,32'd-5976,32'd-6884,32'd436,32'd-2609,32'd-7788,32'd-368,32'd-4299,32'd3981,32'd-22539,32'd-4743,32'd-7705,32'd-7539,32'd-524,32'd-1538,32'd-2587,32'd-3527,32'd-56,32'd-1650,32'd-1630,32'd-2578,32'd-1704,32'd-7265,32'd-7729,32'd-22};
    Wx[34]='{32'd-390,32'd-1538,32'd-456,32'd573,32'd124,32'd967,32'd555,32'd-8867,32'd-2900,32'd2125,32'd183,32'd100,32'd-1728,32'd1827,32'd-1517,32'd-3212,32'd-2066,32'd2980,32'd854,32'd-1718,32'd-1474,32'd1063,32'd-1401,32'd-1264,32'd474,32'd837,32'd1022,32'd-1088,32'd-3063,32'd2114,32'd-5209,32'd4997,32'd2868,32'd4628,32'd453,32'd1270,32'd-3537,32'd-1387,32'd5039,32'd5605,32'd-371,32'd2196,32'd-1821,32'd4433,32'd1179,32'd-223,32'd154,32'd-1405,32'd-491,32'd-1270,32'd2568,32'd2797,32'd1424,32'd2661,32'd5219,32'd-100,32'd3491,32'd-913,32'd1958,32'd-809,32'd1820,32'd2500,32'd83,32'd-391,32'd-3559,32'd1385,32'd2117,32'd5590,32'd-386,32'd2092,32'd2724,32'd-1221,32'd-1655,32'd-1151,32'd-5927,32'd-323,32'd10537,32'd2252,32'd1400,32'd-2207,32'd1617,32'd4001,32'd3339,32'd5058,32'd-2067,32'd5156,32'd1387,32'd2309,32'd-2844,32'd-4108,32'd846,32'd6513,32'd697,32'd-2115,32'd1434,32'd-2888,32'd2551,32'd-6547,32'd-1571,32'd2349,32'd-5014,32'd12773,32'd-3798,32'd14765,32'd-1206,32'd1927,32'd-1258,32'd9096,32'd2126,32'd3,32'd1197,32'd-7348,32'd-1462,32'd6577,32'd563,32'd9907,32'd1469,32'd-3510,32'd3720,32'd-3,32'd580,32'd-6157,32'd-179,32'd5419,32'd1407,32'd7060,32'd5932,32'd-1563,32'd10761,32'd6752,32'd1809,32'd4462,32'd4406,32'd-10546,32'd-2614,32'd1950,32'd908,32'd-651,32'd-5014,32'd-3271,32'd6582,32'd4423,32'd11572,32'd3298,32'd2917,32'd-11904,32'd12216,32'd2746,32'd-7866,32'd-4299,32'd-11259,32'd10351,32'd-5708,32'd-3215,32'd-1772,32'd-16210,32'd5859,32'd2487,32'd8603,32'd957,32'd5717,32'd12597,32'd7675,32'd689,32'd-8051,32'd-546,32'd9487,32'd-20273,32'd1557,32'd-3544,32'd-14287,32'd-12861,32'd-6420,32'd-5458,32'd5576,32'd-8925,32'd-7368,32'd6181,32'd-9301,32'd993,32'd5878,32'd3933,32'd3569,32'd3566,32'd-3415,32'd2565,32'd2294,32'd-87,32'd1148,32'd-5727,32'd-4489,32'd-14091,32'd-405,32'd-1508,32'd4494,32'd-4169,32'd6313,32'd7553,32'd223,32'd-4653,32'd1312,32'd4804,32'd333,32'd-164,32'd-1223,32'd-939,32'd-2119,32'd-3227,32'd682,32'd4235,32'd274,32'd-1303,32'd479,32'd-5424,32'd-176,32'd-391,32'd5629,32'd-2604,32'd2283,32'd2958,32'd-2883,32'd2636,32'd164,32'd196,32'd7285,32'd574,32'd-1068,32'd2014,32'd2534,32'd-9804,32'd1209,32'd155,32'd-3383,32'd1223,32'd7568,32'd-1656,32'd-3627,32'd2026,32'd-3957,32'd-825,32'd-2727,32'd-4370,32'd-3671,32'd613,32'd-4104,32'd-1986,32'd7451,32'd-6796,32'd-4560,32'd1074,32'd-1990,32'd-8125,32'd-2137,32'd-1406,32'd2043,32'd6904,32'd264,32'd99,32'd-5883,32'd7231,32'd-3229,32'd-10673,32'd1381,32'd5029,32'd7543,32'd1063,32'd-4104,32'd-7915,32'd1549,32'd-685,32'd4504,32'd-1715,32'd-1416,32'd-3898,32'd1284,32'd-1608,32'd-5688,32'd-6840,32'd2163,32'd2469,32'd-2030,32'd3566,32'd1982,32'd1864,32'd-5942,32'd-4123,32'd-3071,32'd3645,32'd3041,32'd-4060,32'd-4851,32'd-571,32'd-4345,32'd-1838,32'd-13320,32'd-2254,32'd-755,32'd-9433,32'd5468,32'd214,32'd2366,32'd2,32'd8691,32'd1594,32'd2578,32'd-503,32'd-3496,32'd-2756,32'd-1401,32'd-186,32'd-2551,32'd-4379,32'd3271,32'd513,32'd3476,32'd1794,32'd7885,32'd-4228,32'd-1060,32'd4409,32'd2467,32'd657,32'd-4138,32'd1094,32'd515,32'd-3085,32'd6577,32'd5800,32'd3759,32'd-4890,32'd-1906,32'd-5888,32'd-8408,32'd4008,32'd422,32'd-1221,32'd4575,32'd-2663,32'd-8779,32'd-610,32'd4968,32'd54,32'd-5654,32'd3869,32'd50,32'd3596,32'd12236,32'd-3735,32'd3029,32'd-948,32'd-3864,32'd2783,32'd-3959,32'd-926,32'd17753,32'd11357,32'd-3159,32'd-665,32'd4211,32'd11367,32'd392,32'd-3864,32'd-15283,32'd6215,32'd-3784,32'd12382,32'd-2578,32'd1121,32'd9604,32'd5903,32'd4680,32'd-1195,32'd-4533,32'd-689,32'd1033,32'd2690,32'd-4892,32'd-7241,32'd2467,32'd3356,32'd-513,32'd8403,32'd411,32'd-3066,32'd12617,32'd-5434,32'd3320,32'd4907,32'd4912,32'd-4257,32'd1010,32'd-8149,32'd773,32'd8984,32'd-10908,32'd-5336,32'd917,32'd3586,32'd7182,32'd-3806};
    Wx[35]='{32'd-198,32'd-4685,32'd-1555,32'd-895,32'd2097,32'd-40,32'd4731,32'd-3317,32'd-421,32'd1031,32'd-408,32'd-1434,32'd305,32'd2521,32'd-889,32'd3999,32'd-1082,32'd166,32'd598,32'd2127,32'd-470,32'd-2956,32'd-1912,32'd4494,32'd-2384,32'd1372,32'd-1427,32'd-74,32'd-14,32'd3842,32'd-817,32'd9672,32'd-1904,32'd2939,32'd245,32'd6381,32'd-2121,32'd958,32'd-2493,32'd2060,32'd866,32'd1728,32'd-1267,32'd-684,32'd3366,32'd5068,32'd-4719,32'd331,32'd3046,32'd141,32'd-2502,32'd7480,32'd-1751,32'd1356,32'd-2452,32'd-5898,32'd679,32'd3796,32'd-879,32'd-944,32'd-2493,32'd-230,32'd-1293,32'd-706,32'd2753,32'd3361,32'd-2602,32'd8642,32'd3220,32'd-3303,32'd-621,32'd3325,32'd289,32'd3208,32'd-1400,32'd722,32'd4658,32'd1012,32'd-2573,32'd-2297,32'd4833,32'd2221,32'd-1621,32'd5507,32'd-2741,32'd3474,32'd2199,32'd4584,32'd-3293,32'd1352,32'd3076,32'd2744,32'd-3076,32'd463,32'd-5034,32'd3366,32'd2194,32'd-2995,32'd-2095,32'd-1560,32'd-2086,32'd-1296,32'd-1063,32'd-276,32'd-1511,32'd914,32'd-3671,32'd3557,32'd6206,32'd-4965,32'd3947,32'd-3652,32'd523,32'd-3435,32'd11064,32'd-3767,32'd-8901,32'd2583,32'd-1243,32'd3540,32'd-1881,32'd131,32'd5014,32'd-2054,32'd-1975,32'd-21,32'd208,32'd6997,32'd7846,32'd-11523,32'd6040,32'd8066,32'd8916,32'd-3066,32'd7343,32'd8823,32'd-251,32'd3041,32'd-8452,32'd-8247,32'd4362,32'd8330,32'd10898,32'd-9829,32'd-7241,32'd-12314,32'd18164,32'd-1243,32'd-6450,32'd9863,32'd386,32'd1402,32'd7792,32'd6528,32'd-1968,32'd7421,32'd-3315,32'd-1596,32'd4616,32'd3388,32'd2354,32'd-2800,32'd-11835,32'd-694,32'd-4511,32'd95,32'd7368,32'd3771,32'd2558,32'd-4584,32'd-2519,32'd2065,32'd-969,32'd-11933,32'd3071,32'd-21835,32'd-976,32'd25019,32'd-3896,32'd4313,32'd-2216,32'd22539,32'd828,32'd-7431,32'd3395,32'd1735,32'd-558,32'd10654,32'd870,32'd-759,32'd-9741,32'd5434,32'd5742,32'd-1968,32'd362,32'd2888,32'd-60,32'd-8334,32'd1345,32'd-2736,32'd-4252,32'd6425,32'd-941,32'd4833,32'd-1275,32'd1909,32'd-4973,32'd1044,32'd1859,32'd1085,32'd2824,32'd-1285,32'd4213,32'd-4663,32'd-4411,32'd1691,32'd-250,32'd347,32'd-1195,32'd3876,32'd-2055,32'd-539,32'd3496,32'd1183,32'd3791,32'd3417,32'd-522,32'd-2678,32'd971,32'd4748,32'd1889,32'd975,32'd-671,32'd-1062,32'd-327,32'd-3354,32'd-2797,32'd3942,32'd1064,32'd1467,32'd-727,32'd12,32'd-648,32'd5942,32'd2788,32'd1971,32'd-1242,32'd-3676,32'd-3112,32'd3500,32'd5346,32'd-5039,32'd1494,32'd639,32'd-50,32'd-4565,32'd-2656,32'd2177,32'd641,32'd-6899,32'd-2919,32'd3195,32'd5712,32'd-3276,32'd143,32'd3955,32'd-3491,32'd-12197,32'd716,32'd-6914,32'd-1859,32'd4277,32'd-130,32'd2763,32'd-2127,32'd-12939,32'd-1530,32'd-1972,32'd-4797,32'd5244,32'd-1966,32'd-31,32'd1099,32'd-2983,32'd-1016,32'd-6118,32'd1367,32'd-855,32'd4370,32'd3962,32'd-2746,32'd-6035,32'd-4082,32'd-2290,32'd906,32'd-1168,32'd4731,32'd-94,32'd-2309,32'd-1461,32'd-6093,32'd8691,32'd-4338,32'd2059,32'd-567,32'd-10039,32'd-1816,32'd2084,32'd3688,32'd-4064,32'd3300,32'd411,32'd3793,32'd4462,32'd2556,32'd3371,32'd6821,32'd-5458,32'd1089,32'd-4858,32'd-3747,32'd-3583,32'd2734,32'd6552,32'd-3339,32'd3554,32'd-1988,32'd-6367,32'd4328,32'd2388,32'd1480,32'd8701,32'd-8251,32'd-3620,32'd6508,32'd1749,32'd918,32'd1833,32'd-1673,32'd4599,32'd-1447,32'd6367,32'd947,32'd-83,32'd-3569,32'd551,32'd414,32'd-5371,32'd-2105,32'd84,32'd4233,32'd-4777,32'd1555,32'd-3393,32'd-6113,32'd-8486,32'd-5278,32'd3142,32'd-5961,32'd-10673,32'd-1308,32'd-3212,32'd691,32'd-1549,32'd-167,32'd6694,32'd-8032,32'd-715,32'd-4914,32'd-12871,32'd760,32'd1153,32'd-913,32'd-84,32'd162,32'd-5683,32'd-3854,32'd13,32'd-425,32'd1810,32'd-2463,32'd5273,32'd-106,32'd6381,32'd299,32'd-814,32'd4067,32'd830,32'd603,32'd6865,32'd-513,32'd-6323,32'd-4558,32'd14511,32'd-405,32'd7802,32'd2374,32'd5249,32'd-3249,32'd2534};
    Wx[36]='{32'd459,32'd1117,32'd-1539,32'd148,32'd-646,32'd-4135,32'd3310,32'd-2366,32'd1102,32'd1804,32'd536,32'd-695,32'd2403,32'd-469,32'd-5214,32'd2128,32'd-5688,32'd-353,32'd-607,32'd892,32'd-4111,32'd-257,32'd4572,32'd355,32'd513,32'd-296,32'd-177,32'd-340,32'd268,32'd2178,32'd328,32'd-7084,32'd-2871,32'd638,32'd-450,32'd-7,32'd4174,32'd-1171,32'd-2377,32'd-4257,32'd3593,32'd2305,32'd-1492,32'd-7656,32'd6547,32'd-6352,32'd8520,32'd2358,32'd1984,32'd-1385,32'd1473,32'd-562,32'd2404,32'd2352,32'd1418,32'd-4550,32'd-167,32'd-1161,32'd-19,32'd-314,32'd237,32'd-1459,32'd250,32'd-752,32'd-1624,32'd-2158,32'd-815,32'd-4133,32'd-1049,32'd933,32'd642,32'd-3322,32'd-1958,32'd2976,32'd-1003,32'd-3518,32'd-565,32'd1616,32'd-1112,32'd-5698,32'd-433,32'd-4291,32'd2519,32'd-4965,32'd107,32'd-3679,32'd4135,32'd-1848,32'd1319,32'd371,32'd-1317,32'd-957,32'd5307,32'd-2514,32'd4418,32'd-676,32'd-347,32'd254,32'd-31,32'd-885,32'd-1085,32'd-15097,32'd-1585,32'd2258,32'd-3002,32'd3842,32'd-8286,32'd-12666,32'd-5429,32'd4453,32'd7153,32'd537,32'd-5502,32'd-3410,32'd1339,32'd12939,32'd19550,32'd3105,32'd6401,32'd-457,32'd-589,32'd-1414,32'd-3317,32'd-4858,32'd3950,32'd-3237,32'd-4887,32'd915,32'd-4157,32'd-2156,32'd1306,32'd6489,32'd1507,32'd-534,32'd5708,32'd-6733,32'd5405,32'd2858,32'd1416,32'd16191,32'd-2683,32'd1204,32'd-5449,32'd3869,32'd-7104,32'd11484,32'd10097,32'd-7875,32'd8276,32'd-8852,32'd-8383,32'd1389,32'd-4589,32'd-2102,32'd6435,32'd3854,32'd-5795,32'd-407,32'd6367,32'd-664,32'd4431,32'd-1961,32'd3017,32'd3317,32'd2117,32'd-679,32'd3693,32'd-10976,32'd-218,32'd-1539,32'd1795,32'd-5820,32'd2932,32'd1766,32'd-1662,32'd-12304,32'd-16914,32'd6181,32'd-7382,32'd4538,32'd-4555,32'd-7573,32'd-2841,32'd-2954,32'd546,32'd11845,32'd1496,32'd-70,32'd1477,32'd-1669,32'd114,32'd4895,32'd-4077,32'd102,32'd682,32'd-7578,32'd-2353,32'd7041,32'd-505,32'd-8559,32'd-691,32'd2812,32'd-964,32'd-473,32'd-416,32'd-876,32'd2961,32'd-2290,32'd-1921,32'd-2058,32'd2009,32'd1862,32'd4411,32'd5185,32'd-2646,32'd9140,32'd-1591,32'd-2396,32'd-1608,32'd-599,32'd-439,32'd2653,32'd396,32'd1089,32'd5019,32'd7661,32'd4255,32'd895,32'd-6928,32'd-456,32'd1580,32'd3962,32'd147,32'd4707,32'd-8442,32'd5708,32'd815,32'd-1568,32'd-3579,32'd-3847,32'd-7470,32'd-210,32'd-12333,32'd6000,32'd8710,32'd-7666,32'd3920,32'd1826,32'd-352,32'd-4262,32'd-1106,32'd-8452,32'd93,32'd1638,32'd-221,32'd-871,32'd-92,32'd-4943,32'd-2922,32'd-886,32'd1442,32'd5063,32'd-8876,32'd3076,32'd-1047,32'd2156,32'd-896,32'd7963,32'd2238,32'd24,32'd12089,32'd-1832,32'd4924,32'd16,32'd-4323,32'd896,32'd-474,32'd1756,32'd-2117,32'd1552,32'd-4858,32'd-2232,32'd4040,32'd5385,32'd-315,32'd587,32'd551,32'd-1717,32'd-2578,32'd-1705,32'd-1427,32'd-2398,32'd487,32'd-601,32'd-5874,32'd4357,32'd1562,32'd-2379,32'd1601,32'd-3676,32'd-2539,32'd-2922,32'd-5922,32'd657,32'd-3178,32'd-12148,32'd5292,32'd-4555,32'd1733,32'd-935,32'd-366,32'd-671,32'd2224,32'd-2176,32'd-1962,32'd920,32'd-1833,32'd2514,32'd-9741,32'd-5839,32'd-9472,32'd3271,32'd3073,32'd-1258,32'd5649,32'd-3337,32'd3041,32'd-5874,32'd447,32'd-5141,32'd-4677,32'd5166,32'd1719,32'd-1790,32'd2980,32'd2260,32'd1269,32'd-4809,32'd8662,32'd1979,32'd-3686,32'd783,32'd6000,32'd5683,32'd4191,32'd-9008,32'd1768,32'd-1389,32'd5292,32'd-1213,32'd3554,32'd-5341,32'd3476,32'd4912,32'd-8334,32'd-1728,32'd-2700,32'd-2539,32'd-4406,32'd5800,32'd776,32'd200,32'd-6074,32'd-108,32'd3449,32'd-290,32'd-5585,32'd1752,32'd4602,32'd-5019,32'd3364,32'd4465,32'd1743,32'd-406,32'd-5307,32'd-1909,32'd3093,32'd-1578,32'd-1434,32'd-9008,32'd-1656,32'd-3601,32'd-704,32'd-4694,32'd-9770,32'd3005,32'd5537,32'd-1652,32'd4282,32'd-4682,32'd-1043,32'd785,32'd3061,32'd2829,32'd-498,32'd5200,32'd-8164,32'd-3979,32'd-610,32'd-825};
    Wx[37]='{32'd-784,32'd-660,32'd1374,32'd35,32'd1210,32'd-2098,32'd-618,32'd1026,32'd-1065,32'd2812,32'd5117,32'd-299,32'd210,32'd5268,32'd397,32'd-1741,32'd8852,32'd2060,32'd-1492,32'd-78,32'd-1707,32'd1971,32'd-252,32'd-527,32'd-2193,32'd443,32'd527,32'd2521,32'd-1915,32'd1352,32'd-1673,32'd-1163,32'd-2399,32'd-1478,32'd-2846,32'd-1467,32'd1865,32'd1734,32'd3857,32'd4938,32'd-1141,32'd1552,32'd1601,32'd291,32'd7529,32'd515,32'd1988,32'd1430,32'd3691,32'd1340,32'd-4714,32'd4904,32'd-687,32'd-480,32'd-2209,32'd-3337,32'd-3403,32'd-4367,32'd1932,32'd-4169,32'd-8266,32'd-1384,32'd-1198,32'd-962,32'd5161,32'd-65,32'd838,32'd6313,32'd-2053,32'd1767,32'd0,32'd7622,32'd-140,32'd-2387,32'd4826,32'd-179,32'd2966,32'd640,32'd2187,32'd5097,32'd745,32'd6679,32'd-1023,32'd-3190,32'd-861,32'd721,32'd-809,32'd-3818,32'd-94,32'd-2229,32'd-2083,32'd1030,32'd-1862,32'd431,32'd2810,32'd-1017,32'd3862,32'd8637,32'd-1955,32'd2119,32'd-5751,32'd-14814,32'd1333,32'd-1140,32'd3728,32'd1100,32'd-2333,32'd-6967,32'd-245,32'd-1931,32'd-21113,32'd-1911,32'd-2509,32'd-10244,32'd-10009,32'd3603,32'd11621,32'd-2467,32'd4465,32'd-4067,32'd-660,32'd4682,32'd9892,32'd-3337,32'd-1682,32'd-12158,32'd124,32'd1983,32'd-7714,32'd-7475,32'd2011,32'd-3703,32'd6669,32'd-2,32'd2039,32'd4477,32'd1046,32'd3178,32'd-2022,32'd-7236,32'd4338,32'd-6796,32'd-4418,32'd-5859,32'd5810,32'd14609,32'd-6440,32'd-8779,32'd1196,32'd-485,32'd16,32'd4589,32'd-7724,32'd7910,32'd-2246,32'd-4880,32'd866,32'd1713,32'd9770,32'd-2646,32'd1622,32'd7299,32'd-4499,32'd8525,32'd-393,32'd-3342,32'd-1473,32'd19892,32'd4855,32'd-1279,32'd9941,32'd-9184,32'd-1052,32'd-1240,32'd3464,32'd-5776,32'd-2893,32'd3576,32'd8642,32'd-5244,32'd-1713,32'd-5898,32'd-2277,32'd-15888,32'd-6704,32'd-11738,32'd-838,32'd-1381,32'd2392,32'd-4150,32'd-4116,32'd-2880,32'd1652,32'd1160,32'd7275,32'd1693,32'd-1065,32'd7016,32'd1679,32'd-9438,32'd871,32'd4912,32'd-887,32'd1687,32'd2137,32'd-1552,32'd6674,32'd1972,32'd-4274,32'd841,32'd1401,32'd3774,32'd1624,32'd891,32'd1694,32'd-6591,32'd2814,32'd787,32'd-3781,32'd-817,32'd-2375,32'd-3027,32'd-2281,32'd3918,32'd-2807,32'd6782,32'd827,32'd1376,32'd13876,32'd-491,32'd-828,32'd3417,32'd247,32'd6591,32'd-7094,32'd-408,32'd-8120,32'd534,32'd358,32'd-527,32'd-1406,32'd-1677,32'd-1370,32'd10898,32'd-7651,32'd1619,32'd2171,32'd2207,32'd-2626,32'd3698,32'd6157,32'd-6655,32'd-897,32'd-7368,32'd748,32'd-2292,32'd-3532,32'd-6000,32'd535,32'd4401,32'd-3215,32'd2565,32'd6254,32'd143,32'd2086,32'd3295,32'd4013,32'd-4914,32'd-4384,32'd1867,32'd4384,32'd5019,32'd-1600,32'd-3933,32'd1060,32'd-4597,32'd-1381,32'd-844,32'd6674,32'd1710,32'd-2614,32'd-2531,32'd4189,32'd-4665,32'd-828,32'd-9799,32'd-1040,32'd2929,32'd1557,32'd-1889,32'd-881,32'd-2153,32'd-4377,32'd2344,32'd-192,32'd2170,32'd184,32'd6884,32'd-3115,32'd4396,32'd765,32'd13574,32'd7412,32'd8330,32'd-1190,32'd-4023,32'd4609,32'd757,32'd-490,32'd-8530,32'd4262,32'd5883,32'd1928,32'd5952,32'd-845,32'd-899,32'd6801,32'd5585,32'd-2121,32'd4003,32'd734,32'd-651,32'd-3225,32'd971,32'd-3264,32'd3288,32'd-869,32'd1120,32'd10751,32'd3891,32'd566,32'd6152,32'd-2524,32'd8881,32'd-11435,32'd-2861,32'd-6879,32'd-5405,32'd-3356,32'd8491,32'd3271,32'd2382,32'd3850,32'd19335,32'd829,32'd5317,32'd5834,32'd-1708,32'd-3635,32'd-54,32'd8081,32'd-8974,32'd-275,32'd1962,32'd-1687,32'd4172,32'd4033,32'd3813,32'd2324,32'd-23,32'd4152,32'd5444,32'd10458,32'd7949,32'd3857,32'd1157,32'd5874,32'd5351,32'd-6425,32'd8452,32'd2110,32'd16279,32'd-1766,32'd10185,32'd-1857,32'd-960,32'd7900,32'd3654,32'd7490,32'd1932,32'd-1807,32'd1876,32'd6645,32'd1535,32'd-6875,32'd9584,32'd2829,32'd-3767,32'd2561,32'd5605,32'd-2324,32'd9521,32'd-3269,32'd6035,32'd2200,32'd-290,32'd-2666,32'd2049,32'd-1030,32'd6596};
    Wx[38]='{32'd-501,32'd-4880,32'd-1663,32'd1889,32'd-192,32'd-349,32'd-1437,32'd2294,32'd3481,32'd2944,32'd-1040,32'd5151,32'd-2651,32'd-981,32'd-3181,32'd-1503,32'd328,32'd2661,32'd-530,32'd794,32'd678,32'd2910,32'd-649,32'd-1629,32'd2512,32'd-993,32'd3735,32'd-1978,32'd-5410,32'd1196,32'd-2181,32'd-7153,32'd3579,32'd-6586,32'd357,32'd-975,32'd806,32'd-54,32'd466,32'd2199,32'd-4707,32'd-6367,32'd-4550,32'd848,32'd-4716,32'd2612,32'd-3527,32'd-1605,32'd3251,32'd-3583,32'd205,32'd-1116,32'd-3041,32'd-2775,32'd-1665,32'd-591,32'd-2005,32'd-3601,32'd6030,32'd693,32'd-5766,32'd-6210,32'd-901,32'd304,32'd599,32'd2722,32'd3237,32'd-7963,32'd946,32'd1701,32'd-3308,32'd-974,32'd-1790,32'd1348,32'd173,32'd-5913,32'd2873,32'd-2045,32'd-5566,32'd-1694,32'd641,32'd-14794,32'd-2973,32'd408,32'd-29,32'd-3176,32'd1781,32'd-323,32'd811,32'd1121,32'd-780,32'd-6596,32'd-2653,32'd-872,32'd3708,32'd1926,32'd2819,32'd-3078,32'd-2393,32'd5200,32'd-1638,32'd13691,32'd-798,32'd5429,32'd-3171,32'd-2978,32'd-2177,32'd3464,32'd1822,32'd-3605,32'd-11210,32'd-4204,32'd341,32'd1549,32'd2355,32'd12695,32'd1679,32'd-6694,32'd2470,32'd-1552,32'd637,32'd1455,32'd-236,32'd-70,32'd-93,32'd-240,32'd3920,32'd5039,32'd1925,32'd-1259,32'd-939,32'd-4077,32'd5390,32'd183,32'd2149,32'd-3862,32'd-2622,32'd1596,32'd4553,32'd-2736,32'd11142,32'd-12011,32'd8867,32'd5307,32'd-8242,32'd-11416,32'd14345,32'd-1837,32'd-384,32'd13291,32'd-1538,32'd-8857,32'd7973,32'd3044,32'd-5644,32'd-600,32'd4909,32'd2666,32'd-5952,32'd453,32'd6196,32'd-9687,32'd4875,32'd-2770,32'd96,32'd-4296,32'd-213,32'd5083,32'd1906,32'd133,32'd-4069,32'd-9873,32'd2832,32'd9072,32'd2381,32'd-11132,32'd-5932,32'd-2553,32'd7216,32'd10195,32'd2137,32'd6430,32'd-2832,32'd-2115,32'd-2749,32'd-20078,32'd-7807,32'd-150,32'd2032,32'd645,32'd-197,32'd-6669,32'd-4726,32'd2393,32'd9399,32'd2102,32'd8208,32'd-3435,32'd-2167,32'd-1210,32'd1350,32'd12578,32'd40,32'd-2436,32'd-1003,32'd400,32'd3173,32'd5830,32'd-1384,32'd574,32'd5961,32'd-6977,32'd3996,32'd5180,32'd961,32'd10566,32'd475,32'd3959,32'd-3168,32'd-2868,32'd-1057,32'd-2487,32'd375,32'd3518,32'd2094,32'd6503,32'd-1420,32'd-150,32'd2768,32'd3308,32'd-1939,32'd7646,32'd2802,32'd4907,32'd3547,32'd602,32'd-2927,32'd-4116,32'd8139,32'd4184,32'd5019,32'd6923,32'd3732,32'd224,32'd-14316,32'd2398,32'd-9575,32'd-3251,32'd482,32'd4997,32'd-3027,32'd-4191,32'd-1245,32'd-3381,32'd1650,32'd-4853,32'd5156,32'd2479,32'd434,32'd-3549,32'd629,32'd-1240,32'd13134,32'd8159,32'd-1988,32'd-2221,32'd1076,32'd4353,32'd1872,32'd-819,32'd4958,32'd-3000,32'd-22,32'd4956,32'd715,32'd144,32'd-4968,32'd7592,32'd4895,32'd3674,32'd1651,32'd-7299,32'd224,32'd10224,32'd3420,32'd-835,32'd3710,32'd286,32'd-3869,32'd4345,32'd5087,32'd1550,32'd2480,32'd2110,32'd-3464,32'd-5830,32'd2573,32'd6713,32'd2609,32'd7817,32'd3017,32'd5009,32'd-4277,32'd-3461,32'd2680,32'd10009,32'd2912,32'd-770,32'd-2010,32'd-9282,32'd-2390,32'd2172,32'd2050,32'd193,32'd483,32'd5161,32'd8159,32'd-3100,32'd-7294,32'd736,32'd4882,32'd213,32'd-1501,32'd145,32'd4599,32'd1473,32'd3125,32'd4057,32'd3889,32'd2314,32'd-5166,32'd2049,32'd-2396,32'd-3225,32'd4086,32'd3112,32'd-301,32'd2436,32'd6840,32'd-1336,32'd733,32'd5126,32'd-2595,32'd-8237,32'd-10478,32'd3676,32'd-2441,32'd-1494,32'd3588,32'd-2893,32'd42,32'd-5512,32'd-5053,32'd-2692,32'd3764,32'd-226,32'd2332,32'd9360,32'd-181,32'd3908,32'd1093,32'd-1071,32'd2324,32'd6523,32'd1147,32'd4323,32'd4707,32'd1767,32'd6699,32'd7578,32'd-7387,32'd-2341,32'd-689,32'd5175,32'd986,32'd3559,32'd-3576,32'd4157,32'd-4291,32'd3530,32'd-321,32'd1279,32'd4931,32'd8876,32'd8823,32'd1544,32'd6401,32'd579,32'd-3369,32'd-2653,32'd1511,32'd6674,32'd-2219,32'd-1937,32'd-9047,32'd-2727,32'd2125,32'd9428,32'd3457,32'd7460};
    Wx[39]='{32'd52,32'd2357,32'd1258,32'd-1104,32'd205,32'd694,32'd-996,32'd1374,32'd-170,32'd-2656,32'd1164,32'd91,32'd-3745,32'd-852,32'd-1431,32'd606,32'd5620,32'd-3068,32'd-295,32'd2873,32'd-3286,32'd4816,32'd3857,32'd2387,32'd2191,32'd-1256,32'd-1023,32'd-1235,32'd-5449,32'd-2746,32'd-595,32'd-12412,32'd-3354,32'd1196,32'd-159,32'd4096,32'd-3847,32'd1929,32'd-4841,32'd-6127,32'd-4160,32'd-1866,32'd-53,32'd-2963,32'd-7275,32'd-4909,32'd4843,32'd-2385,32'd4299,32'd-2343,32'd-5336,32'd-3369,32'd-1011,32'd-4687,32'd2266,32'd881,32'd1008,32'd-1530,32'd-1276,32'd-784,32'd-3457,32'd-6752,32'd2858,32'd1232,32'd-4536,32'd-72,32'd1108,32'd1010,32'd423,32'd-1452,32'd-2407,32'd-1798,32'd-3940,32'd5483,32'd-1492,32'd-408,32'd825,32'd14,32'd-577,32'd-1279,32'd250,32'd2600,32'd-597,32'd-5195,32'd489,32'd-4978,32'd619,32'd-65,32'd2531,32'd4912,32'd4377,32'd5786,32'd-98,32'd-6713,32'd3759,32'd-960,32'd626,32'd403,32'd-3845,32'd-3913,32'd-3540,32'd4621,32'd-1901,32'd4719,32'd2464,32'd-3176,32'd-5004,32'd-12666,32'd2080,32'd5893,32'd1560,32'd-37,32'd-4975,32'd4780,32'd489,32'd-5522,32'd3847,32'd604,32'd1369,32'd1322,32'd-3249,32'd2700,32'd956,32'd-1472,32'd5087,32'd-2191,32'd-2707,32'd-1292,32'd1721,32'd2406,32'd270,32'd7866,32'd-1247,32'd2138,32'd8,32'd-2729,32'd4743,32'd1315,32'd8925,32'd-6181,32'd3603,32'd8188,32'd5395,32'd4602,32'd4914,32'd-872,32'd859,32'd-10839,32'd2905,32'd1948,32'd6425,32'd13085,32'd14521,32'd3762,32'd2006,32'd8051,32'd-7690,32'd2958,32'd7773,32'd3156,32'd3879,32'd2470,32'd-7436,32'd-1838,32'd7045,32'd1789,32'd-3164,32'd-2462,32'd-608,32'd-1201,32'd-3676,32'd8198,32'd1440,32'd-2486,32'd-1927,32'd7963,32'd-12519,32'd16318,32'd-5102,32'd4797,32'd-5068,32'd1934,32'd3730,32'd-27148,32'd-5683,32'd4519,32'd4169,32'd-2432,32'd1778,32'd9316,32'd-3586,32'd-17031,32'd-336,32'd-559,32'd-5805,32'd-3046,32'd2475,32'd-10107,32'd-1811,32'd-2790,32'd-3364,32'd3903,32'd501,32'd-2702,32'd1104,32'd-274,32'd9326,32'd-5922,32'd3686,32'd800,32'd1549,32'd-237,32'd9223,32'd-242,32'd4938,32'd4719,32'd-3806,32'd-440,32'd-792,32'd1748,32'd-1700,32'd-1679,32'd5258,32'd-159,32'd760,32'd2145,32'd-2998,32'd2587,32'd175,32'd-2429,32'd-1997,32'd12148,32'd11289,32'd7983,32'd-798,32'd760,32'd-1289,32'd-1324,32'd6748,32'd2141,32'd1156,32'd2551,32'd1080,32'd3999,32'd4477,32'd5209,32'd1306,32'd4501,32'd-470,32'd2790,32'd-5410,32'd8041,32'd6538,32'd-4838,32'd1575,32'd-1755,32'd-1761,32'd-447,32'd-2237,32'd2951,32'd2277,32'd2237,32'd143,32'd906,32'd5942,32'd-3562,32'd1804,32'd-11542,32'd728,32'd1217,32'd2651,32'd5581,32'd-2403,32'd7124,32'd-600,32'd4760,32'd5693,32'd1026,32'd-2592,32'd620,32'd-2016,32'd-5888,32'd-3635,32'd6630,32'd-3791,32'd1403,32'd220,32'd3969,32'd-985,32'd2045,32'd7900,32'd-3652,32'd4172,32'd-1010,32'd-7036,32'd-1954,32'd5820,32'd-5615,32'd8359,32'd2449,32'd788,32'd-175,32'd-4819,32'd-2463,32'd2666,32'd10742,32'd10351,32'd-3991,32'd-246,32'd-1993,32'd-10458,32'd-6269,32'd7553,32'd1496,32'd-426,32'd-5297,32'd-1779,32'd-2165,32'd1379,32'd-2221,32'd-2531,32'd-1989,32'd3034,32'd4362,32'd-651,32'd-1039,32'd-2476,32'd2368,32'd-2556,32'd-582,32'd-1248,32'd3410,32'd-3957,32'd-1291,32'd5844,32'd-344,32'd5708,32'd521,32'd-39,32'd-2437,32'd-2634,32'd-693,32'd-2827,32'd-487,32'd-1169,32'd1755,32'd6484,32'd-1286,32'd-2685,32'd-938,32'd-351,32'd273,32'd4221,32'd-4687,32'd7514,32'd1134,32'd-626,32'd2592,32'd-7832,32'd8574,32'd1668,32'd-3862,32'd-4648,32'd-1129,32'd-2741,32'd2795,32'd9555,32'd-3366,32'd9140,32'd4711,32'd-4511,32'd7636,32'd4069,32'd-1794,32'd951,32'd4411,32'd-1927,32'd8603,32'd-5131,32'd-3823,32'd2004,32'd-1044,32'd-7558,32'd4995,32'd990,32'd1623,32'd-97,32'd-421,32'd-3947,32'd17714,32'd4636,32'd-7436,32'd-1198,32'd4809,32'd-5244,32'd-595,32'd7617,32'd5527,32'd1883,32'd2924};
    Wx[40]='{32'd-586,32'd-165,32'd2381,32'd492,32'd-830,32'd3239,32'd5913,32'd755,32'd3110,32'd-1773,32'd-4555,32'd133,32'd-500,32'd3957,32'd3244,32'd5034,32'd-2297,32'd-1275,32'd1021,32'd-2264,32'd-2177,32'd-917,32'd-449,32'd-2425,32'd-2763,32'd3088,32'd3183,32'd2526,32'd3493,32'd-527,32'd4326,32'd-3056,32'd-1934,32'd-5908,32'd4753,32'd-850,32'd2783,32'd1412,32'd-734,32'd-1961,32'd17,32'd1658,32'd-4970,32'd2034,32'd6088,32'd-233,32'd-3527,32'd5375,32'd-5903,32'd570,32'd6279,32'd2587,32'd1883,32'd-2337,32'd38,32'd1041,32'd106,32'd-610,32'd1078,32'd96,32'd-60,32'd3000,32'd-546,32'd3024,32'd2058,32'd-3508,32'd1211,32'd-5742,32'd709,32'd-656,32'd4025,32'd-3264,32'd661,32'd5322,32'd1812,32'd5942,32'd2180,32'd5971,32'd4929,32'd-3286,32'd-1796,32'd-6166,32'd369,32'd-4257,32'd-2973,32'd1148,32'd295,32'd-4406,32'd5390,32'd1251,32'd5507,32'd328,32'd4770,32'd3657,32'd3264,32'd-3168,32'd2680,32'd4645,32'd-1233,32'd-2985,32'd7968,32'd3820,32'd319,32'd3251,32'd-2042,32'd-783,32'd-14296,32'd10966,32'd-4416,32'd5888,32'd2656,32'd9765,32'd7036,32'd17587,32'd56,32'd-5053,32'd24472,32'd10488,32'd-10058,32'd-4956,32'd4841,32'd-13203,32'd6958,32'd-1781,32'd3908,32'd-450,32'd2719,32'd-7451,32'd-3559,32'd798,32'd4104,32'd612,32'd17148,32'd-214,32'd2543,32'd-5322,32'd3066,32'd-997,32'd-12177,32'd-1915,32'd-10000,32'd11289,32'd-13544,32'd-8217,32'd-6625,32'd8588,32'd-7055,32'd9311,32'd-7382,32'd4069,32'd4670,32'd3425,32'd-2259,32'd7553,32'd751,32'd1229,32'd-11181,32'd-1900,32'd-1036,32'd1882,32'd466,32'd-6357,32'd-15498,32'd7294,32'd-13681,32'd7231,32'd-982,32'd-2386,32'd-1934,32'd609,32'd-4338,32'd6674,32'd2475,32'd19980,32'd3071,32'd-9155,32'd1394,32'd-1459,32'd4401,32'd-2117,32'd-3007,32'd-10371,32'd9741,32'd18164,32'd4162,32'd-7045,32'd466,32'd-5434,32'd-1530,32'd4084,32'd-6972,32'd-15478,32'd6499,32'd3979,32'd-12646,32'd-13437,32'd175,32'd4274,32'd-5893,32'd5605,32'd-2020,32'd-4152,32'd1005,32'd-5122,32'd2866,32'd1228,32'd-11376,32'd1303,32'd8740,32'd2156,32'd5048,32'd1501,32'd1088,32'd9785,32'd-4521,32'd-6713,32'd2338,32'd-3791,32'd4836,32'd-3283,32'd1002,32'd3986,32'd-623,32'd-6103,32'd-4296,32'd3681,32'd-4091,32'd-967,32'd-2536,32'd-3808,32'd-5595,32'd3640,32'd-4240,32'd1940,32'd2685,32'd-136,32'd486,32'd2161,32'd1586,32'd12197,32'd3535,32'd1022,32'd817,32'd-4538,32'd-12470,32'd6079,32'd4221,32'd5649,32'd-1993,32'd-4575,32'd10195,32'd3586,32'd909,32'd-5922,32'd-2103,32'd8842,32'd-639,32'd1752,32'd-3281,32'd2646,32'd731,32'd3564,32'd-4326,32'd3828,32'd-6264,32'd-1732,32'd361,32'd2484,32'd3386,32'd3017,32'd-4760,32'd8164,32'd1282,32'd3820,32'd-1325,32'd-3881,32'd11240,32'd-874,32'd-7519,32'd4079,32'd-175,32'd119,32'd3476,32'd-1781,32'd-4050,32'd10449,32'd-700,32'd-2751,32'd-1009,32'd2883,32'd1012,32'd8432,32'd-4809,32'd7192,32'd-4816,32'd4462,32'd-2595,32'd8369,32'd6064,32'd2482,32'd1269,32'd4418,32'd6240,32'd6918,32'd1445,32'd10839,32'd3708,32'd10312,32'd7666,32'd10078,32'd-689,32'd-750,32'd-1789,32'd11728,32'd3149,32'd1959,32'd-6782,32'd9907,32'd-1141,32'd-5834,32'd3811,32'd9326,32'd-4135,32'd-8115,32'd-315,32'd5317,32'd-5532,32'd7451,32'd3864,32'd-6948,32'd1925,32'd635,32'd1434,32'd1226,32'd2358,32'd2668,32'd4511,32'd7416,32'd7539,32'd9438,32'd1258,32'd-3166,32'd2695,32'd8681,32'd3737,32'd695,32'd-4465,32'd9335,32'd8291,32'd5883,32'd11474,32'd2927,32'd8989,32'd-831,32'd-10136,32'd3459,32'd-808,32'd-10107,32'd-4997,32'd2602,32'd-1439,32'd3010,32'd-881,32'd681,32'd14033,32'd5209,32'd-7338,32'd5488,32'd3205,32'd-10429,32'd5302,32'd-234,32'd-3833,32'd148,32'd-5605,32'd-4726,32'd5957,32'd5708,32'd5122,32'd-3493,32'd2408,32'd-1986,32'd-13886,32'd2634,32'd-6640,32'd14609,32'd-4160,32'd-509,32'd-1787,32'd-9843,32'd6967,32'd12656,32'd7338,32'd-5195,32'd1128,32'd6093,32'd4924,32'd-8120,32'd147,32'd4660};
    Wx[41]='{32'd1949,32'd1076,32'd-2386,32'd-3083,32'd-1027,32'd-2474,32'd396,32'd1508,32'd-463,32'd215,32'd-1459,32'd118,32'd-1297,32'd-4768,32'd-3164,32'd-3325,32'd-3471,32'd2098,32'd2683,32'd-3532,32'd715,32'd-3950,32'd-1061,32'd-2600,32'd2563,32'd-2342,32'd-2059,32'd-791,32'd-1030,32'd3376,32'd2663,32'd-3198,32'd-3881,32'd-4223,32'd1650,32'd-2379,32'd-2443,32'd-4277,32'd11191,32'd6166,32'd700,32'd1561,32'd-3723,32'd-4770,32'd-2480,32'd1663,32'd-9326,32'd-2286,32'd-5966,32'd1146,32'd1217,32'd8076,32'd2412,32'd1551,32'd-3449,32'd-2034,32'd-7,32'd2917,32'd-342,32'd4919,32'd2622,32'd-1866,32'd628,32'd-2198,32'd3623,32'd2235,32'd1372,32'd-433,32'd-3388,32'd576,32'd-1507,32'd-28,32'd-1518,32'd-1844,32'd-2132,32'd-1694,32'd1864,32'd828,32'd-3076,32'd2604,32'd690,32'd-1257,32'd-2885,32'd-1436,32'd2998,32'd-4875,32'd-2626,32'd-22,32'd6,32'd-1303,32'd-1870,32'd2132,32'd5556,32'd1962,32'd-1092,32'd924,32'd266,32'd1595,32'd3911,32'd-1943,32'd252,32'd10361,32'd1313,32'd1641,32'd4252,32'd1334,32'd-3183,32'd2298,32'd-5029,32'd-423,32'd-4006,32'd-3129,32'd3845,32'd-8520,32'd-15449,32'd2220,32'd-646,32'd4165,32'd-1706,32'd-2678,32'd1652,32'd-5737,32'd4333,32'd2351,32'd-4262,32'd7163,32'd4335,32'd812,32'd5859,32'd7685,32'd-1343,32'd-1529,32'd16181,32'd-3757,32'd3461,32'd11523,32'd-3876,32'd-4226,32'd16171,32'd-6479,32'd6757,32'd14111,32'd7744,32'd-3505,32'd-14697,32'd-1601,32'd-4682,32'd4084,32'd-6606,32'd-3415,32'd-1446,32'd144,32'd290,32'd-6958,32'd1213,32'd-4763,32'd6196,32'd-3227,32'd-8666,32'd-733,32'd2883,32'd8911,32'd-707,32'd-1929,32'd-17724,32'd724,32'd3952,32'd3303,32'd4868,32'd2076,32'd-13300,32'd-12363,32'd-5649,32'd1597,32'd-3222,32'd9628,32'd-12744,32'd-1390,32'd1461,32'd5981,32'd14970,32'd-138,32'd-7431,32'd7685,32'd-5151,32'd9584,32'd6655,32'd-1663,32'd2932,32'd1267,32'd-7304,32'd-1967,32'd-12685,32'd-3537,32'd2648,32'd-1564,32'd6811,32'd8032,32'd9775,32'd-3093,32'd-880,32'd-2917,32'd930,32'd798,32'd-30,32'd-506,32'd-517,32'd-5922,32'd1251,32'd1878,32'd-2988,32'd1689,32'd-243,32'd-8403,32'd-6074,32'd-4006,32'd5683,32'd-3535,32'd-2126,32'd-374,32'd-141,32'd1320,32'd-1986,32'd-1967,32'd6118,32'd83,32'd-5776,32'd-3168,32'd-9453,32'd-4045,32'd1370,32'd-12324,32'd-2846,32'd-3439,32'd-4189,32'd3395,32'd-2111,32'd-445,32'd-6904,32'd-1284,32'd-597,32'd3674,32'd3967,32'd-1137,32'd-5834,32'd-6113,32'd10205,32'd906,32'd-3203,32'd938,32'd408,32'd-13232,32'd880,32'd-4047,32'd-1634,32'd3552,32'd1298,32'd-769,32'd-1616,32'd-9121,32'd-521,32'd-6723,32'd3774,32'd-352,32'd4248,32'd1557,32'd-1876,32'd-8759,32'd-469,32'd77,32'd-6772,32'd-4177,32'd-2244,32'd-2366,32'd-915,32'd411,32'd5009,32'd2490,32'd-80,32'd-305,32'd-341,32'd-2330,32'd-971,32'd2145,32'd1201,32'd-5175,32'd-4121,32'd-3359,32'd-799,32'd872,32'd-4064,32'd-8217,32'd-6010,32'd-5458,32'd2349,32'd2924,32'd-6791,32'd-2358,32'd420,32'd3503,32'd7353,32'd-1712,32'd-8247,32'd5493,32'd1800,32'd-8164,32'd-10927,32'd-6044,32'd2304,32'd9443,32'd-9111,32'd3696,32'd-7490,32'd-5322,32'd-5390,32'd-681,32'd-6323,32'd-2056,32'd6274,32'd-2456,32'd4626,32'd153,32'd773,32'd-1505,32'd7495,32'd4052,32'd-2286,32'd-478,32'd-22,32'd-5170,32'd5234,32'd-8300,32'd-2675,32'd642,32'd5639,32'd3024,32'd3027,32'd3723,32'd-1221,32'd5688,32'd2729,32'd4802,32'd-2016,32'd3081,32'd-5703,32'd-1387,32'd5966,32'd6953,32'd-3264,32'd2541,32'd-1514,32'd-828,32'd13828,32'd4599,32'd7089,32'd6230,32'd818,32'd-9824,32'd1035,32'd187,32'd-2373,32'd98,32'd1439,32'd3837,32'd7788,32'd611,32'd2629,32'd-6459,32'd-29,32'd-134,32'd5698,32'd-10156,32'd2119,32'd-1218,32'd3684,32'd-170,32'd6025,32'd-4423,32'd640,32'd-2198,32'd1700,32'd-6181,32'd2318,32'd-1643,32'd-4223,32'd-9287,32'd-364,32'd-7158,32'd6665,32'd5566,32'd239,32'd-2829,32'd460,32'd6088,32'd-12285,32'd802,32'd-1128,32'd-5117,32'd2580,32'd-3725};
    Wx[42]='{32'd-1068,32'd3452,32'd-4758,32'd2030,32'd-770,32'd1817,32'd3779,32'd-894,32'd-722,32'd-3166,32'd-2780,32'd727,32'd572,32'd-6967,32'd-354,32'd1269,32'd-10195,32'd1241,32'd626,32'd1856,32'd1147,32'd-344,32'd-60,32'd-1573,32'd236,32'd-1076,32'd2186,32'd-3068,32'd-984,32'd-2446,32'd-1519,32'd-8481,32'd-1029,32'd-5117,32'd1319,32'd2670,32'd-308,32'd1879,32'd-543,32'd-2797,32'd3015,32'd-3613,32'd-544,32'd-1677,32'd5439,32'd2127,32'd-3637,32'd-1882,32'd711,32'd129,32'd-1141,32'd-5522,32'd1323,32'd1892,32'd-2998,32'd-2878,32'd-171,32'd-2131,32'd2541,32'd-2453,32'd-7006,32'd40,32'd4152,32'd-1756,32'd1062,32'd555,32'd1558,32'd-8994,32'd1437,32'd1131,32'd1048,32'd1041,32'd-2990,32'd385,32'd2081,32'd-5478,32'd-638,32'd824,32'd-764,32'd-1044,32'd-2382,32'd-7451,32'd-3957,32'd-1430,32'd3950,32'd-4208,32'd726,32'd-2288,32'd-4167,32'd-70,32'd-3664,32'd713,32'd-1135,32'd-1618,32'd-1938,32'd-20,32'd-5126,32'd126,32'd-1791,32'd-6411,32'd-989,32'd3847,32'd1690,32'd2504,32'd5864,32'd-3012,32'd-4741,32'd-10761,32'd-3063,32'd-3952,32'd-4355,32'd-1914,32'd-355,32'd11796,32'd10478,32'd-4089,32'd-2235,32'd-2495,32'd342,32'd1788,32'd3422,32'd3918,32'd5292,32'd-3188,32'd-3920,32'd2103,32'd-412,32'd-8535,32'd-6206,32'd-1002,32'd-1741,32'd-1934,32'd-22109,32'd-10341,32'd1757,32'd-938,32'd-4003,32'd4904,32'd-5273,32'd-16552,32'd-3874,32'd-13574,32'd-3337,32'd1871,32'd3007,32'd4499,32'd6064,32'd-9409,32'd-4111,32'd687,32'd-4936,32'd573,32'd10673,32'd16855,32'd-1981,32'd8774,32'd-438,32'd1640,32'd-381,32'd1187,32'd2629,32'd9160,32'd5429,32'd-5249,32'd7797,32'd-3259,32'd-5053,32'd1439,32'd-1618,32'd-2871,32'd1577,32'd5605,32'd3754,32'd-5209,32'd2907,32'd-6489,32'd7988,32'd-14208,32'd740,32'd-4770,32'd2478,32'd-686,32'd-4809,32'd-5317,32'd-1318,32'd-3173,32'd3911,32'd-7592,32'd1727,32'd-4829,32'd-592,32'd-1098,32'd-4040,32'd4868,32'd6313,32'd5483,32'd-8901,32'd-13632,32'd440,32'd-22304,32'd-668,32'd1531,32'd-3361,32'd-3244,32'd4824,32'd-513,32'd8203,32'd5981,32'd-338,32'd-2209,32'd-4372,32'd1500,32'd2968,32'd8217,32'd2113,32'd-654,32'd5947,32'd778,32'd-740,32'd492,32'd444,32'd650,32'd1353,32'd-2751,32'd5288,32'd-3186,32'd5307,32'd1287,32'd4980,32'd-5761,32'd1406,32'd5385,32'd-2205,32'd5458,32'd-2451,32'd-134,32'd-1459,32'd1006,32'd-6958,32'd7475,32'd4440,32'd7631,32'd8310,32'd8779,32'd-14560,32'd-560,32'd-1604,32'd-799,32'd-1805,32'd635,32'd-5117,32'd703,32'd-288,32'd1397,32'd-3115,32'd-1890,32'd463,32'd627,32'd-285,32'd-8901,32'd-5595,32'd3376,32'd1233,32'd-2176,32'd-3215,32'd-3835,32'd874,32'd-2407,32'd-1363,32'd3,32'd-3786,32'd-208,32'd-325,32'd-3442,32'd-26,32'd-243,32'd-2612,32'd7485,32'd-4145,32'd-5048,32'd-115,32'd1170,32'd-6577,32'd351,32'd7260,32'd-1993,32'd2944,32'd729,32'd6445,32'd1425,32'd4541,32'd537,32'd1018,32'd1705,32'd6718,32'd-1514,32'd-1462,32'd-11718,32'd-782,32'd2854,32'd-1809,32'd6210,32'd-6845,32'd-1217,32'd7285,32'd144,32'd7202,32'd6523,32'd-4370,32'd-1934,32'd-9501,32'd-3869,32'd-753,32'd8696,32'd-5229,32'd-7275,32'd6166,32'd4052,32'd2949,32'd275,32'd4907,32'd-114,32'd2407,32'd-1953,32'd8872,32'd-3366,32'd3149,32'd-580,32'd49,32'd619,32'd-1459,32'd2763,32'd-5458,32'd777,32'd3737,32'd-3176,32'd-185,32'd4519,32'd-235,32'd3986,32'd7099,32'd-1756,32'd3435,32'd-624,32'd-1437,32'd-1955,32'd-7963,32'd-10000,32'd-2861,32'd-136,32'd2680,32'd-6972,32'd4899,32'd4750,32'd5756,32'd1953,32'd3093,32'd2238,32'd5678,32'd-8691,32'd-2038,32'd1881,32'd-3378,32'd537,32'd-7309,32'd-755,32'd4106,32'd914,32'd11220,32'd6621,32'd-3593,32'd3354,32'd-1501,32'd837,32'd4550,32'd-3461,32'd515,32'd2020,32'd-3652,32'd-7543,32'd-3327,32'd4375,32'd-3044,32'd-5532,32'd-3566,32'd1657,32'd3115,32'd645,32'd-1531,32'd-5571,32'd431,32'd1041,32'd-6850,32'd8940,32'd3139,32'd-5839,32'd-2631,32'd-1464,32'd3308,32'd396};
    Wx[43]='{32'd394,32'd-1755,32'd-3083,32'd-1658,32'd-6074,32'd-704,32'd-5585,32'd-2905,32'd671,32'd3210,32'd-720,32'd1778,32'd-4360,32'd-658,32'd3530,32'd-5136,32'd-6313,32'd-1887,32'd-3498,32'd-777,32'd2416,32'd451,32'd-1545,32'd-324,32'd-3100,32'd-3571,32'd757,32'd2421,32'd-351,32'd-1516,32'd3168,32'd-7709,32'd3190,32'd-5449,32'd125,32'd-2142,32'd1164,32'd-1523,32'd-1577,32'd-2131,32'd-4184,32'd4506,32'd-351,32'd3393,32'd-615,32'd-2663,32'd-814,32'd2089,32'd-1921,32'd-580,32'd-545,32'd-5664,32'd-1575,32'd2893,32'd1817,32'd-4816,32'd1024,32'd3896,32'd-2968,32'd-3220,32'd-642,32'd1956,32'd-1362,32'd-3706,32'd-4084,32'd1517,32'd-847,32'd-8916,32'd-2011,32'd4323,32'd602,32'd-1163,32'd872,32'd1909,32'd171,32'd3056,32'd1303,32'd4077,32'd-1217,32'd-221,32'd-1470,32'd-2663,32'd-4748,32'd-1278,32'd-2519,32'd69,32'd-367,32'd-1052,32'd-354,32'd-1245,32'd-7651,32'd-4692,32'd809,32'd-1441,32'd-5195,32'd-2380,32'd-6176,32'd1073,32'd-1655,32'd-271,32'd757,32'd-2712,32'd1844,32'd-6464,32'd426,32'd636,32'd-4289,32'd-14541,32'd-812,32'd2602,32'd11982,32'd8544,32'd-4423,32'd-5434,32'd-21855,32'd-7543,32'd2376,32'd4694,32'd2275,32'd-2003,32'd2421,32'd-809,32'd7338,32'd1558,32'd-2714,32'd1936,32'd-2117,32'd-5185,32'd-7280,32'd12812,32'd-6972,32'd-6782,32'd7246,32'd3850,32'd-3203,32'd-5986,32'd-410,32'd2248,32'd-3225,32'd5175,32'd-8041,32'd1571,32'd-10703,32'd10039,32'd18281,32'd-2802,32'd-5698,32'd3984,32'd3876,32'd-16308,32'd11083,32'd2612,32'd-3210,32'd-11181,32'd-4987,32'd406,32'd5371,32'd-1298,32'd-3500,32'd-2058,32'd-7128,32'd-3020,32'd26035,32'd-9082,32'd1254,32'd-608,32'd3447,32'd1024,32'd-2141,32'd1135,32'd3408,32'd-8334,32'd2307,32'd-11914,32'd-3520,32'd2849,32'd-3425,32'd1085,32'd2055,32'd3637,32'd-5434,32'd10566,32'd-13300,32'd16816,32'd4279,32'd-6142,32'd-2678,32'd-5913,32'd-3278,32'd188,32'd4555,32'd3920,32'd-3605,32'd-2070,32'd-5170,32'd-1845,32'd-4562,32'd3464,32'd-6337,32'd3913,32'd5712,32'd-9462,32'd-5610,32'd-2102,32'd-202,32'd-1447,32'd3696,32'd1116,32'd-7719,32'd-3449,32'd-1768,32'd-1133,32'd-3569,32'd-2941,32'd1073,32'd-4521,32'd-7363,32'd-867,32'd-5532,32'd-1696,32'd2371,32'd-125,32'd-6347,32'd3395,32'd-3217,32'd-4494,32'd3149,32'd-1791,32'd-910,32'd2452,32'd5849,32'd-3137,32'd-12490,32'd-2451,32'd-2519,32'd1146,32'd2437,32'd3300,32'd-6948,32'd-5209,32'd1202,32'd-10751,32'd2597,32'd-9394,32'd-14599,32'd1240,32'd-2070,32'd-3544,32'd-1408,32'd-5346,32'd1024,32'd-4472,32'd2717,32'd3515,32'd787,32'd7006,32'd-7700,32'd1750,32'd-5654,32'd3308,32'd3337,32'd-3071,32'd-3891,32'd5385,32'd-700,32'd-271,32'd-1414,32'd-5473,32'd-1256,32'd3559,32'd-1833,32'd-2188,32'd5751,32'd-4399,32'd3535,32'd-1636,32'd-2900,32'd-4465,32'd-6835,32'd2111,32'd-1940,32'd-6708,32'd759,32'd-2231,32'd-505,32'd-7641,32'd548,32'd1483,32'd-4462,32'd-1860,32'd2215,32'd2089,32'd-1056,32'd3190,32'd5415,32'd-6884,32'd-5634,32'd1588,32'd2124,32'd-3715,32'd9550,32'd-16845,32'd1397,32'd1304,32'd-3698,32'd31,32'd6406,32'd266,32'd-2272,32'd2734,32'd-6005,32'd182,32'd-7280,32'd-7612,32'd612,32'd-1972,32'd-7666,32'd-809,32'd-6196,32'd8037,32'd9223,32'd3022,32'd-208,32'd3386,32'd3703,32'd-1392,32'd-737,32'd4348,32'd864,32'd-1135,32'd6113,32'd-11923,32'd-9931,32'd687,32'd3613,32'd-2795,32'd-2580,32'd2634,32'd-2304,32'd-10712,32'd-4228,32'd-5800,32'd-865,32'd-2873,32'd-4645,32'd-4648,32'd-7265,32'd154,32'd-606,32'd-2619,32'd-6186,32'd-3488,32'd10751,32'd2983,32'd5883,32'd3483,32'd-1527,32'd3496,32'd-1019,32'd-3977,32'd-1927,32'd-5200,32'd-6616,32'd-1025,32'd1755,32'd4389,32'd-3801,32'd-12099,32'd1939,32'd13037,32'd2602,32'd2462,32'd6689,32'd-49,32'd-301,32'd-625,32'd-4985,32'd7246,32'd5351,32'd1252,32'd550,32'd-4123,32'd2983,32'd-10634,32'd-1652,32'd-3500,32'd-2468,32'd-4616,32'd1889,32'd6152,32'd-2370,32'd4609,32'd2780,32'd-9638,32'd10224,32'd-8276,32'd-5781,32'd-9912,32'd2091,32'd-7543};
    Wx[44]='{32'd1169,32'd5332,32'd172,32'd1384,32'd-1635,32'd606,32'd5708,32'd407,32'd-478,32'd-848,32'd-2026,32'd1743,32'd-2021,32'd-3044,32'd-4599,32'd-1247,32'd-3232,32'd-2497,32'd-3024,32'd767,32'd-2446,32'd1258,32'd4570,32'd-1778,32'd1782,32'd-469,32'd776,32'd-561,32'd-1555,32'd1287,32'd330,32'd-3708,32'd4755,32'd222,32'd-4790,32'd-1896,32'd283,32'd-670,32'd414,32'd-6503,32'd-339,32'd-3037,32'd-2741,32'd-6474,32'd-4802,32'd1932,32'd4216,32'd-6962,32'd-1843,32'd-21,32'd7124,32'd1376,32'd1350,32'd-1811,32'd2929,32'd2990,32'd-2941,32'd-540,32'd577,32'd-22,32'd-66,32'd-207,32'd6469,32'd-1284,32'd1843,32'd-428,32'd-708,32'd-4353,32'd-1062,32'd-1258,32'd-5415,32'd-2155,32'd-1860,32'd-1573,32'd-284,32'd-253,32'd-104,32'd-2856,32'd-1110,32'd4064,32'd-386,32'd-2474,32'd-562,32'd24,32'd4489,32'd-711,32'd630,32'd2856,32'd4257,32'd2087,32'd-1730,32'd1596,32'd162,32'd1739,32'd4616,32'd-2275,32'd-1063,32'd5449,32'd-1848,32'd-2416,32'd1190,32'd-6708,32'd957,32'd-7211,32'd-2565,32'd-482,32'd-2744,32'd-3491,32'd-220,32'd1936,32'd3955,32'd1630,32'd3041,32'd-6459,32'd6259,32'd-1124,32'd-12519,32'd-2236,32'd1949,32'd1401,32'd1635,32'd-83,32'd-3791,32'd2900,32'd1146,32'd-3181,32'd-1942,32'd-1418,32'd-3198,32'd-11708,32'd3886,32'd1850,32'd-9741,32'd2780,32'd-1287,32'd-3615,32'd-2968,32'd-3305,32'd5610,32'd4289,32'd4838,32'd-16826,32'd-1965,32'd-4921,32'd-11298,32'd-3898,32'd-3447,32'd-6943,32'd-4082,32'd-7685,32'd-1198,32'd571,32'd-2453,32'd6875,32'd-2504,32'd6450,32'd1105,32'd42,32'd-4667,32'd-1495,32'd4140,32'd474,32'd6616,32'd711,32'd2174,32'd-2490,32'd-1624,32'd9448,32'd-566,32'd-6513,32'd-5024,32'd-1480,32'd2592,32'd-3666,32'd1428,32'd-16552,32'd-3107,32'd2471,32'd514,32'd3977,32'd-1362,32'd-10156,32'd2858,32'd2746,32'd-468,32'd-697,32'd-1699,32'd1816,32'd1544,32'd-1887,32'd-2900,32'd-18925,32'd-2430,32'd2619,32'd2071,32'd-2768,32'd2653,32'd19052,32'd-5908,32'd2561,32'd638,32'd7934,32'd2463,32'd-3237,32'd1163,32'd110,32'd-5576,32'd131,32'd-1262,32'd869,32'd1840,32'd-1636,32'd-4255,32'd11767,32'd-9589,32'd6831,32'd6323,32'd7456,32'd-5634,32'd969,32'd-556,32'd-4892,32'd4965,32'd-7695,32'd2088,32'd5249,32'd-2246,32'd822,32'd-4389,32'd-5786,32'd-1840,32'd7875,32'd5483,32'd-2675,32'd1262,32'd2873,32'd-1566,32'd-24,32'd5019,32'd-3190,32'd-2252,32'd-2829,32'd4355,32'd3432,32'd-2961,32'd-6445,32'd5268,32'd1568,32'd5747,32'd3288,32'd-992,32'd4353,32'd-1649,32'd12861,32'd243,32'd5258,32'd3955,32'd-1213,32'd-1329,32'd1950,32'd-5068,32'd787,32'd4003,32'd-2622,32'd-2324,32'd-3271,32'd-3430,32'd7631,32'd-740,32'd1475,32'd513,32'd2236,32'd736,32'd3986,32'd2753,32'd11396,32'd187,32'd5009,32'd2081,32'd-1643,32'd-309,32'd-5976,32'd2524,32'd5385,32'd1923,32'd2486,32'd2316,32'd2956,32'd-4370,32'd1666,32'd1678,32'd1358,32'd2127,32'd4296,32'd-1036,32'd1798,32'd-1232,32'd-6059,32'd3542,32'd748,32'd-1865,32'd12958,32'd-2766,32'd1276,32'd2335,32'd1860,32'd-4448,32'd-9975,32'd-5366,32'd3850,32'd-9824,32'd-4257,32'd-3176,32'd-2053,32'd-9790,32'd-2229,32'd3208,32'd1093,32'd-6127,32'd1961,32'd-5781,32'd-1695,32'd4133,32'd-5708,32'd4868,32'd3278,32'd-3767,32'd1145,32'd-3190,32'd697,32'd-7968,32'd3010,32'd-1705,32'd-2744,32'd-6713,32'd1934,32'd-1903,32'd4465,32'd-1125,32'd-5917,32'd-1281,32'd-2368,32'd-1621,32'd-1181,32'd-1396,32'd-5185,32'd3100,32'd-954,32'd4040,32'd-9,32'd5839,32'd-5161,32'd2834,32'd5717,32'd1015,32'd-4726,32'd642,32'd-3259,32'd3872,32'd-2069,32'd-10146,32'd1372,32'd3547,32'd187,32'd-856,32'd-7651,32'd1999,32'd-113,32'd1892,32'd-7709,32'd1296,32'd-6210,32'd-8388,32'd-1262,32'd-7172,32'd6337,32'd4187,32'd28,32'd-3706,32'd-407,32'd348,32'd-3825,32'd-4150,32'd9672,32'd1567,32'd6689,32'd-4724,32'd8530,32'd-1425,32'd-3254,32'd4108,32'd2443,32'd1643,32'd3652,32'd2353,32'd5874,32'd9150,32'd-6923,32'd2211,32'd1666};
    Wx[45]='{32'd-29,32'd-5000,32'd-3706,32'd-3371,32'd1628,32'd-345,32'd-3059,32'd-1054,32'd761,32'd2893,32'd6708,32'd3715,32'd1241,32'd-464,32'd1760,32'd-520,32'd835,32'd5292,32'd2056,32'd-3818,32'd937,32'd-320,32'd-4331,32'd1167,32'd-2359,32'd2335,32'd2430,32'd2384,32'd-2512,32'd-2264,32'd-65,32'd-2449,32'd-2468,32'd937,32'd-1029,32'd1285,32'd345,32'd-296,32'd-8950,32'd5209,32'd-755,32'd2919,32'd-104,32'd2543,32'd2856,32'd-3007,32'd662,32'd8618,32'd1050,32'd-2362,32'd-1947,32'd-850,32'd-55,32'd-5234,32'd2331,32'd-6342,32'd-830,32'd-1612,32'd2141,32'd-1947,32'd1857,32'd1658,32'd-2132,32'd-3811,32'd-2858,32'd-600,32'd-610,32'd121,32'd6835,32'd3388,32'd-997,32'd2573,32'd2497,32'd1607,32'd2165,32'd2514,32'd10097,32'd12,32'd-3505,32'd-2797,32'd1011,32'd3510,32'd-1994,32'd2561,32'd160,32'd1516,32'd157,32'd563,32'd-2619,32'd-408,32'd-1773,32'd-2071,32'd-184,32'd-3417,32'd965,32'd3789,32'd-3020,32'd-1999,32'd-1057,32'd3918,32'd1618,32'd-1467,32'd877,32'd837,32'd6528,32'd-1091,32'd2631,32'd7065,32'd214,32'd-237,32'd-773,32'd-6264,32'd-1296,32'd-11113,32'd-3881,32'd-4841,32'd2775,32'd4111,32'd3190,32'd-5576,32'd-2966,32'd-5698,32'd-128,32'd-8710,32'd4020,32'd-1179,32'd-546,32'd5083,32'd-3774,32'd2016,32'd-3051,32'd-10732,32'd11474,32'd-11816,32'd-1319,32'd-459,32'd6191,32'd541,32'd-19111,32'd640,32'd-4689,32'd4064,32'd-16083,32'd-623,32'd-5053,32'd19287,32'd13457,32'd4721,32'd-3933,32'd-8935,32'd-2279,32'd2088,32'd-4353,32'd7587,32'd-2834,32'd-12070,32'd-5136,32'd4565,32'd-3874,32'd125,32'd-1922,32'd-5561,32'd-4289,32'd-3576,32'd-2044,32'd-764,32'd2246,32'd-3237,32'd197,32'd-2414,32'd9511,32'd-8701,32'd-2863,32'd10390,32'd-1961,32'd19990,32'd-529,32'd8437,32'd14833,32'd-7670,32'd4257,32'd10585,32'd9658,32'd-9008,32'd-6254,32'd-417,32'd-3979,32'd-6831,32'd-3798,32'd-1436,32'd4108,32'd-11044,32'd9067,32'd1900,32'd9755,32'd-7954,32'd5688,32'd11464,32'd4787,32'd-88,32'd393,32'd11357,32'd-3078,32'd998,32'd-2279,32'd328,32'd-3615,32'd5195,32'd4587,32'd2431,32'd-2783,32'd-2006,32'd-2812,32'd-7954,32'd-1151,32'd1838,32'd4956,32'd2504,32'd-2578,32'd-1006,32'd-371,32'd2792,32'd-3251,32'd4531,32'd-1021,32'd-2897,32'd-4509,32'd-1315,32'd1201,32'd222,32'd-1641,32'd-3405,32'd3591,32'd-1496,32'd-7412,32'd-5878,32'd-222,32'd-97,32'd-1529,32'd4777,32'd-900,32'd-1840,32'd10732,32'd-52,32'd4619,32'd-26,32'd2176,32'd-2812,32'd-3298,32'd-3640,32'd-9462,32'd-5644,32'd-5327,32'd-6064,32'd2548,32'd3703,32'd-4655,32'd-1480,32'd-2404,32'd3933,32'd-5073,32'd-6508,32'd429,32'd-3930,32'd5888,32'd-5620,32'd-600,32'd5610,32'd2954,32'd-489,32'd-3745,32'd-5937,32'd2778,32'd-4328,32'd-6665,32'd-955,32'd-9858,32'd-262,32'd2137,32'd-908,32'd2476,32'd-1422,32'd-5698,32'd-9912,32'd-5292,32'd-733,32'd-6005,32'd2192,32'd797,32'd286,32'd4143,32'd2305,32'd-7143,32'd1940,32'd3579,32'd-1328,32'd988,32'd-4487,32'd408,32'd1245,32'd3002,32'd-2709,32'd141,32'd-206,32'd-2766,32'd6132,32'd-9033,32'd11562,32'd6254,32'd-6542,32'd-3581,32'd-2425,32'd3149,32'd-9184,32'd-9790,32'd4797,32'd8754,32'd1713,32'd-942,32'd1856,32'd-296,32'd-3105,32'd-7797,32'd1215,32'd-1171,32'd3078,32'd-2144,32'd3415,32'd-2709,32'd3103,32'd6665,32'd235,32'd-540,32'd7412,32'd5385,32'd-7294,32'd244,32'd3652,32'd934,32'd2399,32'd3930,32'd675,32'd-5122,32'd-7060,32'd3942,32'd-2479,32'd3750,32'd2398,32'd1270,32'd-4040,32'd2839,32'd-4409,32'd-6684,32'd-2025,32'd8222,32'd-4309,32'd3327,32'd8164,32'd899,32'd2097,32'd1235,32'd-334,32'd-1181,32'd4641,32'd-6875,32'd914,32'd800,32'd-1264,32'd25312,32'd7036,32'd-6640,32'd-4465,32'd9868,32'd3295,32'd-563,32'd1087,32'd101,32'd2770,32'd-204,32'd-452,32'd832,32'd-2149,32'd-2305,32'd-19394,32'd-4711,32'd2464,32'd-8247,32'd-106,32'd722,32'd4367,32'd2592,32'd-5366,32'd-6533,32'd-960,32'd-4758,32'd-3542,32'd-286,32'd-251,32'd-5209,32'd6938};
    Wx[46]='{32'd-582,32'd-491,32'd310,32'd-1315,32'd-1761,32'd2119,32'd1201,32'd1461,32'd113,32'd-1035,32'd490,32'd-865,32'd1442,32'd3713,32'd-3476,32'd-1486,32'd-1977,32'd2252,32'd-1729,32'd2822,32'd2895,32'd2298,32'd-569,32'd547,32'd-410,32'd-1931,32'd2792,32'd1302,32'd-36,32'd365,32'd3041,32'd5761,32'd4975,32'd2626,32'd3718,32'd-1322,32'd-2553,32'd401,32'd-1651,32'd-1013,32'd503,32'd2624,32'd2263,32'd-2395,32'd1070,32'd4001,32'd3984,32'd-4643,32'd-269,32'd-2937,32'd3825,32'd4155,32'd3640,32'd4382,32'd-1402,32'd-11152,32'd3229,32'd5361,32'd-106,32'd-901,32'd-2031,32'd2044,32'd-933,32'd1958,32'd1217,32'd-382,32'd2497,32'd3073,32'd-1006,32'd-1900,32'd-1420,32'd944,32'd4748,32'd3471,32'd-205,32'd5195,32'd4130,32'd3256,32'd-2673,32'd3942,32'd1112,32'd4301,32'd16,32'd4174,32'd541,32'd5063,32'd-14,32'd2509,32'd1765,32'd4003,32'd-1068,32'd4357,32'd-814,32'd3916,32'd169,32'd-3386,32'd-2275,32'd3830,32'd2229,32'd-6010,32'd-2861,32'd-9453,32'd-726,32'd3666,32'd1928,32'd-38,32'd616,32'd1343,32'd-21,32'd-2951,32'd-4313,32'd3562,32'd7348,32'd-2438,32'd6025,32'd-836,32'd8256,32'd3115,32'd530,32'd1878,32'd2395,32'd1003,32'd2043,32'd-4550,32'd-3127,32'd1197,32'd944,32'd6230,32'd-13496,32'd-1781,32'd1080,32'd12246,32'd8134,32'd12070,32'd221,32'd773,32'd1489,32'd-1481,32'd-5234,32'd-14628,32'd549,32'd6835,32'd-14550,32'd-5253,32'd-5625,32'd-3669,32'd-13496,32'd10351,32'd-6088,32'd-3142,32'd-7460,32'd-7978,32'd5102,32'd-5424,32'd-373,32'd-14160,32'd1502,32'd-7031,32'd-2900,32'd-2910,32'd-863,32'd-3928,32'd-8710,32'd-2369,32'd14541,32'd-1505,32'd-2161,32'd7734,32'd1247,32'd-7485,32'd-8969,32'd2885,32'd3623,32'd-15117,32'd1934,32'd-1555,32'd-14335,32'd-906,32'd-5776,32'd-3229,32'd2305,32'd6801,32'd-1802,32'd-1794,32'd3867,32'd-11474,32'd1090,32'd10126,32'd-55,32'd4575,32'd-2115,32'd-9448,32'd266,32'd-70,32'd-7265,32'd1063,32'd-2093,32'd9370,32'd-3833,32'd2344,32'd-787,32'd4978,32'd1069,32'd-41,32'd1657,32'd-1533,32'd-6450,32'd-2086,32'd-1949,32'd2780,32'd-4013,32'd-689,32'd-2337,32'd4130,32'd-8413,32'd-1616,32'd-4838,32'd397,32'd-1040,32'd-1223,32'd1560,32'd-2133,32'd-1547,32'd-4660,32'd-2056,32'd-3959,32'd-1148,32'd85,32'd-2607,32'd-4589,32'd-6630,32'd-5170,32'd-569,32'd-415,32'd-2465,32'd-3806,32'd1873,32'd1170,32'd-1665,32'd-1617,32'd1297,32'd-8916,32'd-4421,32'd1295,32'd3398,32'd1679,32'd-9086,32'd-1563,32'd-1663,32'd1151,32'd-6435,32'd7021,32'd1254,32'd4570,32'd394,32'd5151,32'd-2288,32'd654,32'd-2988,32'd4511,32'd-2299,32'd-6274,32'd2514,32'd-1550,32'd-3759,32'd3066,32'd858,32'd-4238,32'd934,32'd-3334,32'd4699,32'd2170,32'd1644,32'd-1520,32'd1682,32'd-1021,32'd3395,32'd3984,32'd1059,32'd2519,32'd1955,32'd-496,32'd7309,32'd-8779,32'd-660,32'd-4777,32'd-2893,32'd2239,32'd-5297,32'd3195,32'd-4152,32'd3198,32'd-5234,32'd-643,32'd2519,32'd4567,32'd2744,32'd751,32'd168,32'd2678,32'd8198,32'd7016,32'd-194,32'd-2534,32'd-3103,32'd4348,32'd2717,32'd-1198,32'd5595,32'd-928,32'd-3005,32'd-1378,32'd-735,32'd4335,32'd-3586,32'd-2885,32'd-3625,32'd-2402,32'd1436,32'd-1157,32'd3310,32'd-2553,32'd-2197,32'd-2666,32'd-54,32'd-2900,32'd-1623,32'd1635,32'd-3835,32'd3359,32'd-2277,32'd967,32'd-3999,32'd427,32'd-5771,32'd-1551,32'd-3955,32'd-6635,32'd-6137,32'd-2072,32'd567,32'd-1745,32'd-285,32'd-2301,32'd-949,32'd626,32'd5644,32'd481,32'd2105,32'd-3386,32'd-643,32'd4768,32'd4882,32'd2670,32'd-11435,32'd-6191,32'd-57,32'd-5932,32'd-2011,32'd-630,32'd-5170,32'd-2775,32'd3947,32'd1385,32'd-3974,32'd-5009,32'd7055,32'd5688,32'd-11074,32'd-5468,32'd4812,32'd4562,32'd-2534,32'd-4279,32'd-3896,32'd3515,32'd563,32'd-962,32'd1938,32'd2661,32'd3928,32'd3034,32'd-2868,32'd6401,32'd-833,32'd-1069,32'd-1586,32'd-2524,32'd-6284,32'd6191,32'd-7275,32'd-4248,32'd-1145,32'd7133,32'd9829,32'd4223,32'd1922,32'd2687,32'd946,32'd2702};
    Wx[47]='{32'd-2420,32'd-7260,32'd-2692,32'd1049,32'd-1883,32'd1707,32'd-4045,32'd-6572,32'd1113,32'd-996,32'd242,32'd-4003,32'd-8618,32'd-3469,32'd-4599,32'd-5517,32'd-9838,32'd-2347,32'd-5815,32'd-623,32'd76,32'd-1933,32'd-549,32'd-4348,32'd-2949,32'd-4174,32'd-7954,32'd-6572,32'd-8334,32'd2661,32'd-1965,32'd-7153,32'd-3776,32'd736,32'd-7338,32'd-4580,32'd-3566,32'd88,32'd-2543,32'd-2122,32'd-4118,32'd2213,32'd-3930,32'd-2357,32'd577,32'd-4960,32'd202,32'd-5810,32'd-624,32'd-955,32'd-8427,32'd4345,32'd5092,32'd-2536,32'd2430,32'd-17998,32'd-2001,32'd-2211,32'd-2639,32'd-6503,32'd-7817,32'd-4726,32'd-2121,32'd-2819,32'd-1405,32'd-1677,32'd-2553,32'd-4123,32'd503,32'd1087,32'd-1479,32'd-1306,32'd-844,32'd-286,32'd3261,32'd-4501,32'd-8974,32'd1585,32'd799,32'd-8671,32'd-4406,32'd-4899,32'd-3867,32'd-1296,32'd1630,32'd-8925,32'd2097,32'd-2949,32'd-3825,32'd858,32'd-449,32'd-8442,32'd-5722,32'd2309,32'd-7451,32'd-6210,32'd-8159,32'd-4687,32'd-4816,32'd-5947,32'd5107,32'd-5219,32'd-1606,32'd3806,32'd-2868,32'd-1563,32'd-5229,32'd125,32'd-4191,32'd5346,32'd3850,32'd2597,32'd-2460,32'd0,32'd17861,32'd-9770,32'd-6699,32'd2773,32'd-873,32'd292,32'd-815,32'd938,32'd7436,32'd-334,32'd-4807,32'd61,32'd-6723,32'd1390,32'd4572,32'd1082,32'd1093,32'd-4746,32'd-966,32'd-963,32'd-2221,32'd-12402,32'd-4458,32'd-2863,32'd-5517,32'd11230,32'd6064,32'd-1029,32'd-2546,32'd-13583,32'd-2459,32'd5820,32'd-10429,32'd2822,32'd-5395,32'd-5830,32'd-551,32'd-870,32'd-5322,32'd13535,32'd-1944,32'd-3295,32'd2507,32'd-262,32'd-2226,32'd-5791,32'd2534,32'd-15322,32'd-7656,32'd1741,32'd1738,32'd-1611,32'd-89,32'd13320,32'd-3496,32'd740,32'd4416,32'd4045,32'd6250,32'd-15224,32'd6967,32'd-12792,32'd936,32'd-6972,32'd14667,32'd1983,32'd-1245,32'd-2697,32'd16552,32'd-6484,32'd5952,32'd-7968,32'd-6547,32'd-6069,32'd-149,32'd-439,32'd-7602,32'd2148,32'd5034,32'd3020,32'd-17548,32'd-12968,32'd-3471,32'd-16591,32'd-12636,32'd-810,32'd-652,32'd4003,32'd-2587,32'd-2666,32'd-1735,32'd2052,32'd-6411,32'd5581,32'd2827,32'd-1937,32'd-11,32'd-1206,32'd3359,32'd1351,32'd-2883,32'd3986,32'd1425,32'd-4382,32'd-2384,32'd-443,32'd-2032,32'd-2736,32'd1312,32'd-1395,32'd1870,32'd-817,32'd6069,32'd241,32'd1057,32'd-4465,32'd-2492,32'd973,32'd5327,32'd-3488,32'd4575,32'd-3757,32'd4670,32'd-293,32'd-592,32'd7109,32'd-629,32'd3586,32'd4157,32'd2055,32'd6137,32'd13525,32'd5654,32'd545,32'd1232,32'd2712,32'd5673,32'd3566,32'd825,32'd1230,32'd-424,32'd8037,32'd-53,32'd1331,32'd-135,32'd1661,32'd-2792,32'd1123,32'd3054,32'd-1329,32'd-10449,32'd5009,32'd265,32'd6621,32'd2283,32'd6635,32'd-3444,32'd3652,32'd-2016,32'd1898,32'd922,32'd-53,32'd1497,32'd2521,32'd4260,32'd-747,32'd-306,32'd1218,32'd453,32'd5180,32'd7695,32'd-1427,32'd-994,32'd2734,32'd3293,32'd846,32'd2517,32'd8583,32'd3867,32'd8027,32'd-5073,32'd180,32'd2084,32'd-4609,32'd696,32'd334,32'd3872,32'd4699,32'd3469,32'd312,32'd-1276,32'd-1026,32'd-2376,32'd4943,32'd-3928,32'd-1103,32'd-9858,32'd-6782,32'd-1311,32'd-1328,32'd5561,32'd3793,32'd-834,32'd-12578,32'd-3012,32'd-5678,32'd7758,32'd1379,32'd-6411,32'd-13437,32'd4521,32'd-3645,32'd-4113,32'd-1636,32'd-5004,32'd-1956,32'd-3022,32'd991,32'd1776,32'd5434,32'd-1221,32'd-1997,32'd-2971,32'd6152,32'd4775,32'd-1778,32'd-3918,32'd-2012,32'd-922,32'd5263,32'd4909,32'd4040,32'd-4760,32'd-162,32'd8281,32'd-3410,32'd1341,32'd2463,32'd5693,32'd416,32'd5063,32'd-4548,32'd8178,32'd-190,32'd-3916,32'd-12421,32'd-1606,32'd-2236,32'd8593,32'd-3679,32'd-7158,32'd8437,32'd-4265,32'd4470,32'd7939,32'd399,32'd-560,32'd-7685,32'd-12041,32'd-4326,32'd1335,32'd-6860,32'd-6660,32'd-1002,32'd-1745,32'd-8959,32'd-2915,32'd4987,32'd-8403,32'd2065,32'd-1744,32'd2360,32'd-2768,32'd-859,32'd-1168,32'd-1343,32'd-3745,32'd-1696,32'd-1901,32'd9550,32'd10527,32'd3850,32'd-2053,32'd1135,32'd-1619,32'd-8354};
    Wx[48]='{32'd-537,32'd-2158,32'd2563,32'd398,32'd-1657,32'd-793,32'd2030,32'd-173,32'd-2357,32'd-2795,32'd3591,32'd593,32'd3439,32'd2617,32'd57,32'd9716,32'd-2098,32'd-3781,32'd-1480,32'd-2888,32'd916,32'd1032,32'd503,32'd-848,32'd3044,32'd-294,32'd2188,32'd788,32'd-346,32'd-1281,32'd-385,32'd-2751,32'd6850,32'd1406,32'd2285,32'd-562,32'd4228,32'd3059,32'd-778,32'd-1458,32'd-869,32'd-1089,32'd6762,32'd1450,32'd338,32'd2978,32'd10429,32'd1583,32'd-1158,32'd2375,32'd-1004,32'd3803,32'd-956,32'd-957,32'd-1113,32'd6665,32'd-109,32'd-1561,32'd297,32'd-1408,32'd2963,32'd5356,32'd4863,32'd3710,32'd6762,32'd-1590,32'd2844,32'd-1025,32'd-2609,32'd-2944,32'd3779,32'd2321,32'd3483,32'd1665,32'd-891,32'd1110,32'd6962,32'd1740,32'd-1204,32'd-219,32'd1613,32'd8076,32'd1997,32'd1759,32'd-7641,32'd1614,32'd-1697,32'd318,32'd-1433,32'd-515,32'd-50,32'd331,32'd3496,32'd2138,32'd5791,32'd-2658,32'd1794,32'd1979,32'd2770,32'd1072,32'd7250,32'd-2208,32'd820,32'd-118,32'd2114,32'd322,32'd-6855,32'd2568,32'd-4792,32'd432,32'd6962,32'd-1395,32'd5571,32'd8027,32'd-3273,32'd513,32'd425,32'd5092,32'd1517,32'd-500,32'd1867,32'd1511,32'd-4716,32'd-5820,32'd-649,32'd5346,32'd-610,32'd3,32'd-9589,32'd-6147,32'd4221,32'd9116,32'd-2,32'd-7836,32'd-6489,32'd-112,32'd1353,32'd5366,32'd5742,32'd-8085,32'd940,32'd-13232,32'd5317,32'd-7294,32'd-13388,32'd-10615,32'd-7333,32'd-1766,32'd-5629,32'd4094,32'd3886,32'd3701,32'd-1730,32'd-2697,32'd1683,32'd4992,32'd-1669,32'd2963,32'd-5107,32'd-1372,32'd-6074,32'd9482,32'd-3569,32'd5439,32'd-10878,32'd81,32'd-5991,32'd7929,32'd-258,32'd283,32'd-3041,32'd-5659,32'd2580,32'd1986,32'd-1400,32'd8652,32'd9384,32'd-574,32'd10917,32'd-3034,32'd-3188,32'd-4230,32'd1168,32'd2790,32'd-7460,32'd-22929,32'd7597,32'd12265,32'd1862,32'd817,32'd-1983,32'd-3630,32'd4182,32'd5297,32'd-6079,32'd-68,32'd-4672,32'd3542,32'd2479,32'd-13134,32'd-1553,32'd-8208,32'd-1669,32'd-1668,32'd1667,32'd-93,32'd-4809,32'd-12197,32'd364,32'd-459,32'd-6015,32'd-80,32'd-2661,32'd-3950,32'd-3901,32'd-8588,32'd4934,32'd-8325,32'd3708,32'd-1590,32'd1006,32'd-880,32'd-1658,32'd-2575,32'd-6406,32'd-2639,32'd-596,32'd-2275,32'd-4399,32'd-5927,32'd-5688,32'd-8525,32'd-8227,32'd-10478,32'd-8842,32'd3593,32'd1566,32'd-1546,32'd456,32'd-2288,32'd-3881,32'd-2692,32'd-7426,32'd-9326,32'd-10390,32'd1701,32'd7983,32'd-4384,32'd-541,32'd-3432,32'd3103,32'd-2183,32'd-4709,32'd-5405,32'd-5200,32'd-1512,32'd4265,32'd-2309,32'd-4929,32'd5581,32'd88,32'd-4284,32'd-690,32'd3854,32'd-13457,32'd-3195,32'd-1799,32'd-2060,32'd408,32'd-4653,32'd-3801,32'd6010,32'd2592,32'd-429,32'd-2568,32'd-7158,32'd7861,32'd-10498,32'd-8281,32'd2592,32'd2968,32'd4108,32'd-8598,32'd-3417,32'd-1689,32'd-1317,32'd-3225,32'd-3830,32'd7500,32'd2495,32'd117,32'd-3959,32'd-6596,32'd6440,32'd3586,32'd-4731,32'd-7045,32'd-6186,32'd-8955,32'd-10410,32'd-1098,32'd1762,32'd161,32'd5893,32'd-1033,32'd-12968,32'd-83,32'd-4714,32'd1583,32'd2534,32'd4736,32'd452,32'd2396,32'd348,32'd-6713,32'd-1106,32'd-1051,32'd2176,32'd5380,32'd-1734,32'd-7402,32'd-520,32'd4711,32'd-305,32'd4396,32'd5590,32'd-3525,32'd-4716,32'd-473,32'd-4375,32'd1794,32'd1582,32'd104,32'd1227,32'd-2678,32'd3833,32'd-5708,32'd-2829,32'd-4101,32'd-6660,32'd6547,32'd-1156,32'd886,32'd4721,32'd-5981,32'd1894,32'd-7065,32'd-4824,32'd-2883,32'd6567,32'd5717,32'd-7216,32'd-5683,32'd81,32'd-9135,32'd502,32'd8139,32'd-3032,32'd4057,32'd234,32'd-87,32'd973,32'd7246,32'd-3647,32'd-139,32'd-7622,32'd-422,32'd-3107,32'd-5185,32'd-6191,32'd3693,32'd7475,32'd2095,32'd1333,32'd-2381,32'd-3603,32'd1505,32'd3076,32'd-3732,32'd358,32'd-1535,32'd4975,32'd-5029,32'd-606,32'd-14785,32'd4055,32'd-11884,32'd88,32'd3208,32'd-4355,32'd7080,32'd-35,32'd-2978,32'd9819,32'd10927,32'd-6376,32'd-1503,32'd-13271,32'd-2666,32'd-3691};
    Wx[49]='{32'd145,32'd9926,32'd-215,32'd-316,32'd2229,32'd-1645,32'd-361,32'd-175,32'd-143,32'd4741,32'd12080,32'd5556,32'd-3552,32'd-2841,32'd-1688,32'd-3129,32'd1463,32'd6220,32'd-1087,32'd-2753,32'd3732,32'd4167,32'd-1826,32'd2729,32'd974,32'd-2868,32'd400,32'd-849,32'd1645,32'd335,32'd-2054,32'd1309,32'd4785,32'd4567,32'd-4411,32'd3264,32'd-5517,32'd-3769,32'd1169,32'd-349,32'd1903,32'd5805,32'd-6308,32'd5083,32'd-6181,32'd485,32'd1987,32'd7026,32'd1844,32'd-994,32'd1052,32'd952,32'd2103,32'd182,32'd4782,32'd1894,32'd8037,32'd4455,32'd4074,32'd-2810,32'd-747,32'd1311,32'd-4338,32'd-191,32'd1743,32'd-1391,32'd4174,32'd1694,32'd745,32'd4025,32'd-1529,32'd-45,32'd-4499,32'd739,32'd-192,32'd-761,32'd-129,32'd1092,32'd-2238,32'd177,32'd3518,32'd5317,32'd3620,32'd3110,32'd4633,32'd5361,32'd-1098,32'd1287,32'd-695,32'd-222,32'd1049,32'd6005,32'd-659,32'd-1842,32'd4648,32'd1010,32'd-3808,32'd4208,32'd841,32'd2340,32'd-1419,32'd14179,32'd2207,32'd4750,32'd-1925,32'd1610,32'd-1205,32'd-5678,32'd-850,32'd-7651,32'd2668,32'd-4389,32'd-5249,32'd14082,32'd16582,32'd909,32'd4672,32'd-8159,32'd2646,32'd2290,32'd-1678,32'd-1097,32'd-4003,32'd1062,32'd-2152,32'd1401,32'd-1093,32'd-4069,32'd-1458,32'd-2100,32'd-481,32'd-3959,32'd17861,32'd-9291,32'd-1370,32'd529,32'd8208,32'd2452,32'd-1600,32'd12001,32'd456,32'd858,32'd-18623,32'd-172,32'd15253,32'd5043,32'd12578,32'd9150,32'd-1091,32'd226,32'd3972,32'd-2415,32'd7749,32'd5488,32'd4133,32'd-10517,32'd12412,32'd1149,32'd-206,32'd446,32'd3693,32'd6523,32'd-9555,32'd-3664,32'd8608,32'd-2514,32'd3110,32'd-10234,32'd-2141,32'd-49,32'd706,32'd-15859,32'd-5903,32'd-1522,32'd-558,32'd-5053,32'd-4919,32'd5825,32'd-3701,32'd1336,32'd497,32'd1680,32'd-4479,32'd-2531,32'd-2270,32'd-10625,32'd2875,32'd-4321,32'd-4321,32'd-2291,32'd-975,32'd-5566,32'd-10732,32'd-1422,32'd5825,32'd-8764,32'd-3974,32'd678,32'd4174,32'd-2675,32'd-3398,32'd9731,32'd-2012,32'd838,32'd-2215,32'd-158,32'd6718,32'd-759,32'd1224,32'd6826,32'd-6318,32'd-168,32'd1560,32'd-2646,32'd-3825,32'd1241,32'd-502,32'd1511,32'd-1345,32'd2595,32'd1445,32'd-1657,32'd-1000,32'd-4294,32'd3129,32'd-3918,32'd-2778,32'd1055,32'd-990,32'd1896,32'd-3242,32'd-4775,32'd-5859,32'd1475,32'd-4335,32'd-2025,32'd-1571,32'd-4836,32'd-7231,32'd-914,32'd-4501,32'd-5258,32'd1437,32'd10673,32'd11357,32'd897,32'd1462,32'd-4714,32'd-3049,32'd-418,32'd-11992,32'd-7338,32'd2261,32'd4504,32'd-2619,32'd-4702,32'd-5429,32'd-1046,32'd-938,32'd7475,32'd162,32'd-6079,32'd2944,32'd-8935,32'd58,32'd1762,32'd1329,32'd10048,32'd-1843,32'd5195,32'd1666,32'd-2609,32'd-2493,32'd-1623,32'd-163,32'd-4375,32'd-7446,32'd-7275,32'd1304,32'd-127,32'd-1499,32'd2883,32'd1682,32'd-2795,32'd-750,32'd-6684,32'd1142,32'd-3012,32'd-978,32'd-2059,32'd-1141,32'd-624,32'd-3994,32'd-2607,32'd-5585,32'd-730,32'd375,32'd-9438,32'd4489,32'd1372,32'd-4404,32'd9023,32'd4050,32'd-4970,32'd-7636,32'd5878,32'd3666,32'd1765,32'd9057,32'd4787,32'd-2169,32'd4042,32'd386,32'd2724,32'd492,32'd4099,32'd12363,32'd-7509,32'd-3808,32'd-831,32'd9980,32'd-4709,32'd-3266,32'd1145,32'd-527,32'd22,32'd1114,32'd2340,32'd1163,32'd2878,32'd-2279,32'd6982,32'd-3522,32'd2636,32'd165,32'd-4436,32'd6025,32'd4245,32'd-2017,32'd-6577,32'd5200,32'd-487,32'd172,32'd-1247,32'd-3759,32'd1038,32'd16132,32'd-3066,32'd-2059,32'd-3063,32'd-603,32'd1658,32'd-4914,32'd-1328,32'd-114,32'd3476,32'd3374,32'd4978,32'd5024,32'd3271,32'd3093,32'd-1013,32'd-254,32'd1356,32'd-1087,32'd2619,32'd4672,32'd1849,32'd6166,32'd8798,32'd7133,32'd1314,32'd4792,32'd-66,32'd4387,32'd1331,32'd1647,32'd-4667,32'd-1708,32'd4741,32'd1058,32'd7197,32'd3630,32'd-5161,32'd9277,32'd-3376,32'd4721,32'd-6459,32'd-59,32'd-1774,32'd2218,32'd-3149,32'd-4548,32'd7949,32'd-4064,32'd971,32'd-6821,32'd13779,32'd2685,32'd6059};
    Wx[50]='{32'd-8,32'd5322,32'd-4401,32'd2883,32'd2114,32'd941,32'd5688,32'd5224,32'd1192,32'd2961,32'd10195,32'd-2517,32'd5620,32'd1824,32'd-2866,32'd-1058,32'd4118,32'd2137,32'd-853,32'd1126,32'd-2476,32'd-126,32'd1749,32'd214,32'd1844,32'd1560,32'd-208,32'd-800,32'd-622,32'd1145,32'd-2770,32'd5048,32'd-4086,32'd-569,32'd-1245,32'd4462,32'd4770,32'd1791,32'd-2861,32'd188,32'd2795,32'd-447,32'd-242,32'd-3125,32'd-1821,32'd4433,32'd7187,32'd12832,32'd419,32'd-731,32'd33,32'd-619,32'd2073,32'd739,32'd1550,32'd2580,32'd-2032,32'd-5463,32'd1552,32'd-6308,32'd-5346,32'd369,32'd-2498,32'd1032,32'd-3547,32'd3278,32'd961,32'd-974,32'd-157,32'd-1851,32'd4099,32'd3066,32'd-4946,32'd2364,32'd357,32'd-2169,32'd3818,32'd4025,32'd1150,32'd5839,32'd-171,32'd7792,32'd-3352,32'd5156,32'd2453,32'd1325,32'd599,32'd-1324,32'd-1094,32'd4160,32'd3090,32'd327,32'd2285,32'd-52,32'd4653,32'd3361,32'd5390,32'd3464,32'd1052,32'd2407,32'd-2670,32'd4145,32'd1856,32'd-6083,32'd-1932,32'd2529,32'd-1340,32'd-318,32'd-328,32'd-2478,32'd-194,32'd-1538,32'd-3969,32'd-3164,32'd11845,32'd2963,32'd11396,32'd1953,32'd4985,32'd2641,32'd-154,32'd-4672,32'd875,32'd-7563,32'd1507,32'd-4938,32'd775,32'd-2778,32'd-2047,32'd-8720,32'd3986,32'd-2946,32'd-5283,32'd14785,32'd5166,32'd6030,32'd-698,32'd5053,32'd2778,32'd-7631,32'd3161,32'd-979,32'd-7636,32'd-1512,32'd-5000,32'd-7304,32'd11601,32'd-5961,32'd1330,32'd-4008,32'd8330,32'd1578,32'd4792,32'd11640,32'd-3352,32'd3176,32'd-6660,32'd3166,32'd3283,32'd4426,32'd-2254,32'd728,32'd8212,32'd-6655,32'd-12978,32'd531,32'd-2058,32'd12792,32'd525,32'd-2370,32'd3796,32'd11279,32'd59,32'd-9804,32'd1878,32'd-1750,32'd458,32'd8569,32'd2885,32'd3178,32'd-2744,32'd8032,32'd-3603,32'd-5986,32'd4770,32'd-2934,32'd2958,32'd-3864,32'd5664,32'd2307,32'd-5761,32'd-7377,32'd-3981,32'd2087,32'd10234,32'd1159,32'd-902,32'd17031,32'd-1223,32'd-5068,32'd-228,32'd-21074,32'd-2324,32'd787,32'd-5571,32'd455,32'd3208,32'd-1663,32'd2286,32'd343,32'd-4873,32'd4975,32'd-1083,32'd2893,32'd5771,32'd-6318,32'd8305,32'd4365,32'd-302,32'd5869,32'd-2033,32'd-1023,32'd2880,32'd-1658,32'd2393,32'd3496,32'd5458,32'd1784,32'd1525,32'd-4399,32'd1842,32'd-2778,32'd-111,32'd3430,32'd-1754,32'd6313,32'd-5590,32'd55,32'd-8603,32'd50,32'd892,32'd5961,32'd5439,32'd7861,32'd7524,32'd878,32'd-3952,32'd-697,32'd-434,32'd1180,32'd-1512,32'd-2062,32'd-2836,32'd8417,32'd1248,32'd1159,32'd3212,32'd-4816,32'd1430,32'd1038,32'd-3728,32'd4479,32'd5317,32'd-892,32'd-5947,32'd-572,32'd-2685,32'd-3740,32'd-1221,32'd-1791,32'd7919,32'd-5195,32'd1061,32'd-1455,32'd1406,32'd1871,32'd-933,32'd6650,32'd5991,32'd6923,32'd-5092,32'd-12636,32'd2451,32'd554,32'd4584,32'd-6748,32'd1279,32'd-814,32'd1781,32'd6215,32'd-1927,32'd-4306,32'd3872,32'd-5375,32'd7587,32'd-2308,32'd1132,32'd-27,32'd2406,32'd2707,32'd354,32'd-3330,32'd-6987,32'd3308,32'd-6567,32'd-377,32'd149,32'd-755,32'd446,32'd-16,32'd3571,32'd2973,32'd-140,32'd3742,32'd4880,32'd-3598,32'd1677,32'd14423,32'd-740,32'd2631,32'd-798,32'd2093,32'd2111,32'd3364,32'd191,32'd509,32'd-942,32'd4028,32'd635,32'd-2166,32'd-603,32'd1028,32'd9399,32'd4814,32'd3505,32'd1707,32'd3588,32'd-3547,32'd-2047,32'd3874,32'd-1857,32'd12236,32'd961,32'd4770,32'd6040,32'd1441,32'd-3112,32'd664,32'd-1922,32'd886,32'd-1975,32'd-3676,32'd1522,32'd4504,32'd928,32'd-858,32'd1673,32'd-8208,32'd1091,32'd7368,32'd-1285,32'd1994,32'd500,32'd-1705,32'd4589,32'd4797,32'd-5913,32'd1147,32'd5219,32'd-1345,32'd4445,32'd1883,32'd1262,32'd10039,32'd1240,32'd-8256,32'd-1389,32'd10117,32'd378,32'd-5356,32'd-3244,32'd-2391,32'd-7656,32'd4013,32'd8657,32'd501,32'd2012,32'd-6474,32'd-1802,32'd7954,32'd2697,32'd6967,32'd859,32'd-5512,32'd8759,32'd-9301,32'd6289,32'd-908,32'd1508,32'd5786};
    Wx[51]='{32'd362,32'd-661,32'd112,32'd-1336,32'd-1534,32'd-1273,32'd2604,32'd899,32'd-311,32'd-1596,32'd9018,32'd1429,32'd-3205,32'd1763,32'd1442,32'd-5639,32'd-1306,32'd932,32'd-664,32'd-1667,32'd132,32'd-1317,32'd108,32'd-2081,32'd3662,32'd-1251,32'd-255,32'd-1227,32'd2995,32'd2517,32'd3166,32'd3605,32'd2687,32'd-2448,32'd2205,32'd5239,32'd-717,32'd370,32'd-6513,32'd1981,32'd-446,32'd1838,32'd1115,32'd971,32'd1108,32'd-1662,32'd11923,32'd2697,32'd-508,32'd-1452,32'd1278,32'd382,32'd1270,32'd-1884,32'd-1379,32'd3562,32'd2568,32'd4467,32'd3750,32'd797,32'd-236,32'd-1434,32'd1411,32'd2403,32'd1553,32'd3049,32'd-583,32'd10429,32'd169,32'd493,32'd-2137,32'd2359,32'd-4494,32'd3657,32'd-714,32'd-4516,32'd-1566,32'd-94,32'd-877,32'd3354,32'd-1456,32'd10410,32'd4277,32'd10341,32'd-1745,32'd-472,32'd2534,32'd644,32'd2269,32'd-23,32'd-1553,32'd2839,32'd-809,32'd2827,32'd2156,32'd1024,32'd-260,32'd391,32'd-1029,32'd-483,32'd1132,32'd11718,32'd2873,32'd-679,32'd-7167,32'd910,32'd2290,32'd-2167,32'd3854,32'd-8476,32'd9233,32'd3781,32'd-781,32'd7465,32'd7387,32'd-12919,32'd-6259,32'd-3513,32'd-7792,32'd258,32'd-4143,32'd3547,32'd1938,32'd7119,32'd1224,32'd-8447,32'd4916,32'd1657,32'd5874,32'd-2341,32'd115,32'd8715,32'd-9785,32'd2293,32'd548,32'd4414,32'd7524,32'd1230,32'd-5844,32'd7490,32'd-2283,32'd-1834,32'd-11230,32'd6240,32'd-10068,32'd11728,32'd-952,32'd-4033,32'd-5791,32'd4846,32'd10634,32'd3940,32'd4794,32'd-3229,32'd4843,32'd3312,32'd14648,32'd742,32'd7490,32'd-1091,32'd262,32'd5668,32'd3405,32'd-1876,32'd15771,32'd-3684,32'd-749,32'd10458,32'd228,32'd-904,32'd-12773,32'd-2709,32'd-20,32'd-12734,32'd2775,32'd11611,32'd-1320,32'd2491,32'd-15175,32'd5468,32'd-734,32'd17412,32'd-1202,32'd-398,32'd-5107,32'd-8959,32'd101,32'd-7646,32'd-640,32'd1673,32'd-3063,32'd1572,32'd-4626,32'd1728,32'd-4543,32'd2432,32'd3002,32'd-6381,32'd-4973,32'd2004,32'd891,32'd-982,32'd1824,32'd4897,32'd252,32'd-1589,32'd3166,32'd-1441,32'd412,32'd1387,32'd-3215,32'd1949,32'd-2281,32'd-4460,32'd-117,32'd-2402,32'd3691,32'd4328,32'd1533,32'd2036,32'd3139,32'd-2756,32'd-3537,32'd-3955,32'd4301,32'd2517,32'd5029,32'd-886,32'd-3254,32'd3205,32'd-890,32'd-542,32'd6430,32'd3295,32'd5351,32'd-3552,32'd2358,32'd2983,32'd-1622,32'd-3806,32'd579,32'd-10156,32'd-6611,32'd5102,32'd-9418,32'd-5239,32'd-14482,32'd3125,32'd-2080,32'd-1793,32'd637,32'd1978,32'd5839,32'd-12197,32'd-8173,32'd-7783,32'd-2871,32'd3686,32'd313,32'd-913,32'd280,32'd5996,32'd-619,32'd-5869,32'd7133,32'd114,32'd3518,32'd1990,32'd-2152,32'd-56,32'd4851,32'd928,32'd-5317,32'd-7207,32'd-33,32'd6591,32'd420,32'd6196,32'd-4543,32'd-1383,32'd1043,32'd2915,32'd-270,32'd-1588,32'd4978,32'd-2683,32'd3081,32'd6738,32'd-3688,32'd1844,32'd4812,32'd718,32'd2741,32'd258,32'd-4,32'd-2917,32'd-2617,32'd13310,32'd-2492,32'd2741,32'd2437,32'd-1945,32'd-8115,32'd-643,32'd-372,32'd-622,32'd1755,32'd-2089,32'd2430,32'd-5454,32'd-244,32'd-1350,32'd-864,32'd-2310,32'd3291,32'd-1666,32'd6191,32'd1418,32'd1262,32'd2932,32'd9741,32'd-2131,32'd-1173,32'd1424,32'd9184,32'd-339,32'd5976,32'd4262,32'd3571,32'd2010,32'd-4138,32'd2382,32'd7519,32'd2778,32'd3591,32'd-3186,32'd1152,32'd7788,32'd1279,32'd-4052,32'd1020,32'd-3754,32'd-2583,32'd565,32'd-4326,32'd-9199,32'd3422,32'd858,32'd-6196,32'd-2648,32'd-478,32'd-1951,32'd-5073,32'd-2709,32'd-2347,32'd-1368,32'd-1907,32'd-8334,32'd5302,32'd-962,32'd-4414,32'd-2807,32'd7055,32'd-3669,32'd770,32'd8037,32'd89,32'd-110,32'd-3408,32'd11337,32'd-2314,32'd-1159,32'd5917,32'd-687,32'd4162,32'd3632,32'd7397,32'd384,32'd-6635,32'd1114,32'd3684,32'd379,32'd1003,32'd50,32'd12636,32'd-8525,32'd9433,32'd-1159,32'd-3146,32'd-3500,32'd7514,32'd6401,32'd-4,32'd17177,32'd2243,32'd-469,32'd6083,32'd9375,32'd2551,32'd-3002};
    Wx[52]='{32'd-1489,32'd1262,32'd-2768,32'd-1322,32'd1990,32'd-26,32'd-5673,32'd-7514,32'd-2502,32'd-2702,32'd-2851,32'd2541,32'd-2114,32'd-2399,32'd-3547,32'd-1708,32'd459,32'd-2854,32'd145,32'd1162,32'd4914,32'd-626,32'd-1444,32'd0,32'd767,32'd-1756,32'd2150,32'd887,32'd2797,32'd1683,32'd410,32'd4375,32'd-295,32'd2351,32'd-4116,32'd-3049,32'd-2412,32'd3471,32'd2897,32'd-1290,32'd-1018,32'd-1817,32'd2492,32'd2133,32'd2198,32'd3691,32'd4279,32'd-8540,32'd-1051,32'd895,32'd-4697,32'd4777,32'd1979,32'd1334,32'd1883,32'd2003,32'd481,32'd-367,32'd-1577,32'd2543,32'd5029,32'd-4904,32'd4003,32'd-1323,32'd-4379,32'd-2349,32'd-2509,32'd-1842,32'd253,32'd-18,32'd-1000,32'd-292,32'd7177,32'd-3415,32'd2380,32'd-1668,32'd5600,32'd1303,32'd1914,32'd534,32'd-1373,32'd446,32'd1910,32'd-1531,32'd3881,32'd346,32'd2153,32'd3476,32'd-3049,32'd1038,32'd-4841,32'd-8559,32'd-4536,32'd4729,32'd-91,32'd-208,32'd-1052,32'd-2873,32'd-53,32'd-1253,32'd-1950,32'd-2199,32'd1093,32'd-4421,32'd5361,32'd475,32'd5991,32'd-12822,32'd165,32'd-3657,32'd-2692,32'd-2922,32'd277,32'd-11718,32'd5097,32'd-16582,32'd-11845,32'd5961,32'd4067,32'd3217,32'd3635,32'd-4245,32'd6171,32'd-2602,32'd-949,32'd4294,32'd-8652,32'd-624,32'd-14580,32'd6748,32'd-185,32'd5014,32'd-13242,32'd5209,32'd-2355,32'd-2170,32'd-5131,32'd4089,32'd6318,32'd-5712,32'd935,32'd-1734,32'd7836,32'd903,32'd7324,32'd-7597,32'd-15644,32'd-8120,32'd4252,32'd1257,32'd-3679,32'd4809,32'd6269,32'd-5039,32'd5659,32'd-2381,32'd9086,32'd-2653,32'd6035,32'd-4416,32'd-6772,32'd-16376,32'd6030,32'd-6469,32'd7958,32'd2125,32'd-664,32'd-7524,32'd-1627,32'd3642,32'd4138,32'd288,32'd1962,32'd19667,32'd390,32'd-306,32'd-10517,32'd9985,32'd-2116,32'd5883,32'd-10458,32'd-9370,32'd4333,32'd14560,32'd9916,32'd-5830,32'd-1347,32'd6660,32'd2502,32'd-1790,32'd15107,32'd10595,32'd378,32'd1867,32'd-11806,32'd9082,32'd-9687,32'd-8168,32'd-6718,32'd-3132,32'd-3107,32'd-13564,32'd-2590,32'd35,32'd-158,32'd1296,32'd-4401,32'd-1220,32'd-1300,32'd-2039,32'd-8710,32'd427,32'd251,32'd501,32'd2346,32'd-4042,32'd-181,32'd-1558,32'd-1878,32'd-445,32'd-21,32'd1524,32'd-7114,32'd4672,32'd-2937,32'd-4531,32'd1511,32'd-673,32'd961,32'd-2966,32'd788,32'd-1503,32'd-2985,32'd-7431,32'd-1205,32'd2739,32'd498,32'd1716,32'd-202,32'd-6997,32'd2680,32'd-3823,32'd3752,32'd-5922,32'd-199,32'd-4887,32'd3388,32'd-1234,32'd-1396,32'd-3764,32'd-2170,32'd-8085,32'd-2182,32'd-2249,32'd-3708,32'd-5092,32'd-971,32'd2724,32'd-6323,32'd-183,32'd256,32'd125,32'd-156,32'd4978,32'd-10136,32'd-4699,32'd-2060,32'd-9311,32'd-3332,32'd-755,32'd4777,32'd622,32'd6225,32'd214,32'd1408,32'd2915,32'd-2785,32'd-5683,32'd-2624,32'd3120,32'd-565,32'd3400,32'd5092,32'd1903,32'd-3286,32'd2731,32'd2341,32'd-3034,32'd-734,32'd-1916,32'd-606,32'd1933,32'd-1868,32'd2131,32'd-9501,32'd1424,32'd-2636,32'd-3449,32'd-1206,32'd-5063,32'd-2177,32'd-143,32'd-207,32'd1726,32'd1182,32'd-559,32'd-254,32'd3381,32'd-4399,32'd-1651,32'd-1551,32'd-1915,32'd-3366,32'd-1566,32'd-4550,32'd-5185,32'd-8613,32'd7622,32'd-7421,32'd354,32'd7080,32'd4033,32'd-5161,32'd-2990,32'd4223,32'd-4724,32'd-3269,32'd-3771,32'd-106,32'd-1796,32'd291,32'd2266,32'd-10458,32'd-10146,32'd4138,32'd4667,32'd1319,32'd3547,32'd-10048,32'd-10878,32'd-5517,32'd-10185,32'd7089,32'd-4326,32'd1469,32'd-4763,32'd-4650,32'd6005,32'd1307,32'd4240,32'd-9951,32'd-7773,32'd2724,32'd1655,32'd-826,32'd-663,32'd-1237,32'd5463,32'd-4365,32'd-2556,32'd2697,32'd-7265,32'd-3459,32'd-4697,32'd-12021,32'd-316,32'd-10146,32'd1569,32'd-847,32'd-11113,32'd-3876,32'd-6650,32'd4504,32'd-5043,32'd-1580,32'd4892,32'd-5595,32'd-1671,32'd2517,32'd-2075,32'd1610,32'd-5439,32'd-1137,32'd331,32'd2438,32'd-6152,32'd-4858,32'd-7504,32'd-5478,32'd3813,32'd1531,32'd7080,32'd-5693,32'd-5346,32'd-2340,32'd6015,32'd-194,32'd-8144,32'd-5449,32'd-1710};
    Wx[53]='{32'd117,32'd2116,32'd-330,32'd-1658,32'd1151,32'd-2064,32'd-4123,32'd-3442,32'd1547,32'd455,32'd-5747,32'd-922,32'd-1849,32'd1729,32'd1118,32'd-7744,32'd3833,32'd3190,32'd-503,32'd1308,32'd1293,32'd1194,32'd974,32'd1538,32'd0,32'd-1531,32'd1596,32'd-1490,32'd-3002,32'd-3256,32'd-376,32'd-1127,32'd2941,32'd3300,32'd-3781,32'd3112,32'd1282,32'd-2093,32'd-4396,32'd3608,32'd1751,32'd2712,32'd1437,32'd-3347,32'd-900,32'd368,32'd-3522,32'd-759,32'd1525,32'd-3039,32'd-820,32'd897,32'd1721,32'd-2807,32'd405,32'd8823,32'd-128,32'd3493,32'd411,32'd3291,32'd79,32'd-2032,32'd-675,32'd1964,32'd-2934,32'd2258,32'd-1136,32'd-4909,32'd3215,32'd745,32'd-6918,32'd-8247,32'd4416,32'd-2683,32'd-2851,32'd495,32'd12236,32'd-1370,32'd-3781,32'd1462,32'd-2432,32'd-5893,32'd-856,32'd2878,32'd3725,32'd4555,32'd-1781,32'd-1386,32'd-2498,32'd-1407,32'd-5649,32'd-948,32'd-137,32'd1158,32'd-954,32'd-1262,32'd2047,32'd-939,32'd2126,32'd4260,32'd2045,32'd20371,32'd3244,32'd-2000,32'd4428,32'd3349,32'd-1502,32'd5126,32'd1995,32'd15,32'd-5043,32'd-3083,32'd14,32'd-2194,32'd9394,32'd-2707,32'd-7910,32'd-3251,32'd388,32'd-2758,32'd-4,32'd1650,32'd143,32'd4064,32'd-187,32'd-769,32'd2088,32'd6284,32'd-23984,32'd3640,32'd-244,32'd12099,32'd-6840,32'd16572,32'd-535,32'd-3251,32'd-2990,32'd3500,32'd-5117,32'd-4592,32'd-1843,32'd-17880,32'd-13066,32'd6215,32'd11806,32'd-771,32'd373,32'd2448,32'd10507,32'd14677,32'd-11845,32'd-3120,32'd11240,32'd7031,32'd-2519,32'd-1541,32'd7011,32'd25,32'd2186,32'd1034,32'd3845,32'd7070,32'd-8691,32'd-2758,32'd8139,32'd-1495,32'd-2427,32'd6762,32'd1502,32'd130,32'd2012,32'd-4877,32'd-2568,32'd2222,32'd-6376,32'd17900,32'd1334,32'd-388,32'd6567,32'd-3791,32'd327,32'd-5131,32'd-5717,32'd3071,32'd-9213,32'd-1,32'd4533,32'd-20449,32'd2075,32'd-702,32'd3305,32'd-2954,32'd-4001,32'd1216,32'd3994,32'd8530,32'd-1754,32'd-6152,32'd7963,32'd-23867,32'd-3295,32'd-2332,32'd-1627,32'd-1126,32'd-3166,32'd-1444,32'd5498,32'd1282,32'd-3081,32'd378,32'd-3806,32'd3659,32'd-1849,32'd1685,32'd9663,32'd-7236,32'd-10058,32'd4650,32'd668,32'd1213,32'd3046,32'd953,32'd-1128,32'd-916,32'd-3049,32'd816,32'd-1213,32'd1839,32'd-535,32'd1243,32'd-6777,32'd2451,32'd9755,32'd7773,32'd6372,32'd-2509,32'd-299,32'd2741,32'd3669,32'd2685,32'd-1,32'd7216,32'd-4797,32'd4094,32'd9912,32'd-1810,32'd7060,32'd6982,32'd-2080,32'd7905,32'd-10683,32'd1646,32'd6860,32'd513,32'd2792,32'd-2497,32'd3771,32'd4394,32'd340,32'd-4594,32'd634,32'd2302,32'd830,32'd-4050,32'd15380,32'd3481,32'd2319,32'd-1953,32'd-709,32'd1845,32'd3439,32'd1490,32'd2734,32'd53,32'd-2077,32'd3386,32'd-4338,32'd2902,32'd1713,32'd-5883,32'd861,32'd3640,32'd-2712,32'd5664,32'd2110,32'd-8564,32'd-3991,32'd4858,32'd-3942,32'd3486,32'd3347,32'd-276,32'd-969,32'd5903,32'd7050,32'd5332,32'd7207,32'd-12822,32'd3769,32'd3864,32'd65,32'd-392,32'd-10429,32'd2272,32'd-3005,32'd-3203,32'd-481,32'd6513,32'd-2091,32'd-6821,32'd-4772,32'd2012,32'd-5893,32'd3034,32'd4182,32'd-3930,32'd2089,32'd6127,32'd3305,32'd6611,32'd6181,32'd930,32'd-7890,32'd304,32'd-6816,32'd-2142,32'd-352,32'd4299,32'd2521,32'd8798,32'd-2344,32'd3881,32'd871,32'd5942,32'd6176,32'd-2958,32'd8188,32'd3891,32'd1944,32'd676,32'd4953,32'd3330,32'd-3110,32'd-9589,32'd3801,32'd-1453,32'd7729,32'd8476,32'd-3791,32'd-1657,32'd1329,32'd508,32'd-7949,32'd-281,32'd-3430,32'd-273,32'd4279,32'd1464,32'd-265,32'd1901,32'd1258,32'd-1579,32'd7866,32'd-3168,32'd-6347,32'd-4536,32'd-319,32'd-1086,32'd-5976,32'd-2230,32'd-1357,32'd-3352,32'd7016,32'd-1553,32'd-2222,32'd4248,32'd4162,32'd5415,32'd-4750,32'd2089,32'd-1495,32'd5341,32'd-2595,32'd-1920,32'd-10136,32'd1734,32'd-7954,32'd6381,32'd-676,32'd9868,32'd2187,32'd-470,32'd-5664,32'd-4499,32'd-2756,32'd1905,32'd4604,32'd3586,32'd5874,32'd5283};
    Wx[54]='{32'd-2885,32'd-5112,32'd-1523,32'd3850,32'd225,32'd-3244,32'd1015,32'd404,32'd-3740,32'd1507,32'd-3132,32'd-1119,32'd-3059,32'd2944,32'd-3444,32'd-2553,32'd6269,32'd1665,32'd1030,32'd-177,32'd1083,32'd1724,32'd4492,32'd899,32'd3398,32'd4597,32'd2052,32'd-997,32'd1361,32'd1887,32'd-1149,32'd-829,32'd-3085,32'd623,32'd1937,32'd255,32'd-1185,32'd-1683,32'd-5771,32'd3107,32'd891,32'd-1448,32'd-3945,32'd-1188,32'd2095,32'd583,32'd-8173,32'd841,32'd2609,32'd-1191,32'd9956,32'd-1624,32'd5351,32'd2125,32'd2597,32'd7358,32'd-2478,32'd478,32'd979,32'd8935,32'd-513,32'd2238,32'd2780,32'd2800,32'd-327,32'd1420,32'd-976,32'd-834,32'd-1322,32'd-980,32'd-4125,32'd2012,32'd1932,32'd1888,32'd1107,32'd-2105,32'd-1734,32'd243,32'd-6357,32'd-2673,32'd-268,32'd4682,32'd-3920,32'd-6147,32'd2316,32'd-6147,32'd97,32'd-1247,32'd3796,32'd2344,32'd228,32'd-3295,32'd877,32'd-1589,32'd-2932,32'd-1759,32'd9033,32'd-3754,32'd-911,32'd3681,32'd-399,32'd-4475,32'd2124,32'd521,32'd-8208,32'd827,32'd-8789,32'd-5292,32'd5546,32'd196,32'd-9790,32'd6567,32'd-6928,32'd2009,32'd4086,32'd12412,32'd9799,32'd-633,32'd4770,32'd4914,32'd-2095,32'd4814,32'd-820,32'd-3105,32'd657,32'd-116,32'd-3215,32'd1026,32'd11464,32'd3571,32'd2489,32'd10117,32'd-4765,32'd-3669,32'd2705,32'd-4174,32'd878,32'd4250,32'd8642,32'd-11181,32'd4814,32'd-6806,32'd146,32'd-2792,32'd-17460,32'd-6899,32'd7314,32'd-13886,32'd8217,32'd-3103,32'd5595,32'd16035,32'd10087,32'd3925,32'd-4912,32'd4704,32'd8530,32'd-1726,32'd-10253,32'd-1044,32'd964,32'd1412,32'd17753,32'd7377,32'd2211,32'd468,32'd2022,32'd-18701,32'd2368,32'd-3066,32'd4746,32'd4401,32'd7114,32'd-8789,32'd-3395,32'd-1058,32'd2648,32'd1032,32'd13808,32'd-3127,32'd-4240,32'd137,32'd-1987,32'd-14375,32'd2149,32'd-6323,32'd2445,32'd-1303,32'd4816,32'd1359,32'd-6181,32'd441,32'd-3891,32'd2257,32'd1210,32'd3383,32'd4343,32'd-1370,32'd-3393,32'd12089,32'd2543,32'd-2524,32'd-1263,32'd-9018,32'd-2447,32'd-1098,32'd-964,32'd-1506,32'd3408,32'd-2556,32'd-4526,32'd2199,32'd2646,32'd5283,32'd4704,32'd-6459,32'd-10771,32'd-1226,32'd-3710,32'd-382,32'd976,32'd2352,32'd-2602,32'd-2795,32'd-3752,32'd-399,32'd2427,32'd-3137,32'd-4743,32'd5170,32'd734,32'd1239,32'd2111,32'd-8803,32'd-5810,32'd-4472,32'd-3642,32'd-2883,32'd-2070,32'd2736,32'd742,32'd7929,32'd-3122,32'd-3483,32'd1293,32'd-9213,32'd-6660,32'd1057,32'd1462,32'd7216,32'd-3720,32'd-4409,32'd4089,32'd-5361,32'd3796,32'd1547,32'd-4362,32'd2536,32'd-2590,32'd48,32'd-560,32'd-1922,32'd-5385,32'd1137,32'd-520,32'd-191,32'd-2683,32'd-4929,32'd588,32'd-3142,32'd14,32'd-5664,32'd-2756,32'd-3295,32'd-1821,32'd-6865,32'd-3935,32'd-2360,32'd1986,32'd-2490,32'd-535,32'd-9160,32'd-71,32'd-2053,32'd-293,32'd-9062,32'd1843,32'd5112,32'd-4802,32'd4067,32'd-4660,32'd-12519,32'd-5688,32'd4594,32'd-6259,32'd-5239,32'd2690,32'd1396,32'd3266,32'd-2374,32'd2083,32'd836,32'd-41,32'd-5556,32'd-3510,32'd-694,32'd3830,32'd2812,32'd292,32'd-10957,32'd-9848,32'd3615,32'd-901,32'd6928,32'd2135,32'd-2500,32'd-1973,32'd3200,32'd-5566,32'd-4042,32'd-5058,32'd3056,32'd1931,32'd428,32'd-1546,32'd-2861,32'd2149,32'd-6918,32'd3535,32'd1907,32'd1911,32'd2239,32'd3627,32'd-7636,32'd248,32'd-2773,32'd-3239,32'd-5527,32'd1497,32'd9057,32'd1049,32'd5541,32'd-2089,32'd-7304,32'd6679,32'd-4172,32'd-4020,32'd-4812,32'd-1844,32'd363,32'd-826,32'd-9970,32'd1206,32'd-5034,32'd2824,32'd1361,32'd-4260,32'd-5942,32'd1256,32'd-1027,32'd-1359,32'd780,32'd-382,32'd719,32'd-2271,32'd5126,32'd-6684,32'd-5869,32'd6586,32'd-5336,32'd1506,32'd-8110,32'd3090,32'd3115,32'd-5424,32'd-133,32'd-1333,32'd-3420,32'd-897,32'd-3403,32'd-3220,32'd-829,32'd3366,32'd-4228,32'd4086,32'd-4565,32'd5537,32'd4680,32'd2624,32'd6630,32'd-3256,32'd1386,32'd758,32'd-5683,32'd-3974,32'd-1279,32'd8349,32'd3979,32'd-2778,32'd-560};
    Wx[55]='{32'd-334,32'd-960,32'd667,32'd1856,32'd-2719,32'd-3935,32'd1132,32'd-3737,32'd927,32'd2570,32'd4230,32'd201,32'd-242,32'd-4494,32'd449,32'd2421,32'd-2973,32'd-1025,32'd-2373,32'd233,32'd-2131,32'd137,32'd-3686,32'd-62,32'd-1538,32'd-812,32'd-5224,32'd-2000,32'd-5722,32'd-1093,32'd-128,32'd-3627,32'd-936,32'd-1689,32'd-5937,32'd5981,32'd-5151,32'd-2585,32'd-7397,32'd-2993,32'd1186,32'd-3281,32'd314,32'd-505,32'd-1839,32'd224,32'd6733,32'd-4650,32'd-1939,32'd-1557,32'd-2458,32'd-1502,32'd-3498,32'd2937,32'd2893,32'd-3955,32'd-100,32'd1845,32'd3332,32'd-464,32'd-3830,32'd-3657,32'd-3537,32'd-4824,32'd-83,32'd1712,32'd-1644,32'd-5693,32'd-5058,32'd-2155,32'd60,32'd-1015,32'd-2238,32'd-3571,32'd-2462,32'd-3576,32'd-5737,32'd-3867,32'd-2238,32'd-2080,32'd1113,32'd4077,32'd2934,32'd-4775,32'd-6181,32'd679,32'd-102,32'd397,32'd720,32'd1647,32'd-1572,32'd-1170,32'd-260,32'd-3315,32'd-1579,32'd-3022,32'd-2802,32'd-1028,32'd-4841,32'd-2578,32'd718,32'd15283,32'd-1741,32'd-1215,32'd-5517,32'd1927,32'd-3745,32'd9248,32'd-6577,32'd-5810,32'd14033,32'd5332,32'd-1012,32'd-15068,32'd5668,32'd9096,32'd-6416,32'd796,32'd2690,32'd-375,32'd-928,32'd-2135,32'd2100,32'd-3464,32'd1965,32'd1973,32'd6376,32'd5229,32'd687,32'd-1022,32'd884,32'd582,32'd-7099,32'd4245,32'd3049,32'd3527,32'd1242,32'd2321,32'd1927,32'd-5214,32'd4025,32'd616,32'd-137,32'd3107,32'd-15576,32'd-3151,32'd5483,32'd-1811,32'd526,32'd-6474,32'd1971,32'd-8198,32'd-12119,32'd9272,32'd-7246,32'd6835,32'd3881,32'd423,32'd-8310,32'd1172,32'd2995,32'd15117,32'd946,32'd-1478,32'd-8461,32'd-1654,32'd-2213,32'd-138,32'd1232,32'd156,32'd898,32'd-5205,32'd-2705,32'd-5405,32'd-2012,32'd3674,32'd1264,32'd1644,32'd13564,32'd8906,32'd6000,32'd6816,32'd-3952,32'd-1605,32'd-79,32'd15517,32'd-3769,32'd-2648,32'd-521,32'd376,32'd-1574,32'd-5502,32'd-4577,32'd-2061,32'd804,32'd-14941,32'd2160,32'd-2293,32'd1318,32'd4208,32'd1922,32'd7368,32'd-1759,32'd1084,32'd1129,32'd-1697,32'd4147,32'd8403,32'd-2988,32'd-1956,32'd1918,32'd-2624,32'd-718,32'd-7358,32'd2917,32'd-1787,32'd1519,32'd1566,32'd-2006,32'd784,32'd-2541,32'd-3527,32'd-828,32'd-793,32'd5527,32'd-1209,32'd3408,32'd-1492,32'd2479,32'd1890,32'd-2476,32'd6782,32'd-2438,32'd2966,32'd3659,32'd3654,32'd-2171,32'd910,32'd3574,32'd8652,32'd-4077,32'd-6225,32'd-253,32'd-5185,32'd-2310,32'd-617,32'd2934,32'd5034,32'd-2407,32'd3559,32'd2971,32'd3181,32'd-6845,32'd1983,32'd-778,32'd8686,32'd5332,32'd-653,32'd680,32'd-5878,32'd589,32'd-9516,32'd5786,32'd5009,32'd8056,32'd3891,32'd-2404,32'd18378,32'd-480,32'd1466,32'd-4853,32'd883,32'd-2624,32'd-2766,32'd-1461,32'd2047,32'd3315,32'd-1680,32'd1004,32'd-593,32'd-289,32'd2587,32'd-4226,32'd7607,32'd3740,32'd4555,32'd-955,32'd3637,32'd-5039,32'd895,32'd-2285,32'd42,32'd-3471,32'd-3540,32'd9936,32'd4455,32'd-4050,32'd8105,32'd-1871,32'd5727,32'd-496,32'd-2174,32'd-5864,32'd-1938,32'd1167,32'd-2861,32'd-2900,32'd1352,32'd-4580,32'd2270,32'd-6416,32'd-3361,32'd6347,32'd-1483,32'd1994,32'd-1518,32'd3793,32'd-5112,32'd3188,32'd4160,32'd2166,32'd-3930,32'd-3708,32'd3334,32'd2592,32'd494,32'd-2758,32'd-488,32'd-10839,32'd-1870,32'd-401,32'd5898,32'd924,32'd-471,32'd-5380,32'd3547,32'd2381,32'd1827,32'd3896,32'd2121,32'd-1723,32'd-189,32'd-7729,32'd-2280,32'd-2287,32'd5693,32'd12529,32'd96,32'd-1518,32'd1239,32'd-1514,32'd1229,32'd-9487,32'd-572,32'd-571,32'd9067,32'd2687,32'd1538,32'd5507,32'd1439,32'd-4453,32'd-5126,32'd1783,32'd2897,32'd1190,32'd9096,32'd1850,32'd2788,32'd447,32'd3239,32'd2038,32'd1541,32'd-6015,32'd858,32'd-2915,32'd2215,32'd3408,32'd-4382,32'd-6982,32'd3300,32'd-4562,32'd2834,32'd-2158,32'd-1715,32'd-10732,32'd8339,32'd-3295,32'd7885,32'd429,32'd-5390,32'd1511,32'd5454,32'd-3029,32'd-9658,32'd693,32'd2006,32'd-4602,32'd7763,32'd-5000,32'd1170};
    Wx[56]='{32'd-4067,32'd6372,32'd1017,32'd2,32'd-1558,32'd739,32'd-2320,32'd7436,32'd-746,32'd-2919,32'd-4890,32'd-1329,32'd3691,32'd-4963,32'd-4714,32'd4206,32'd-7753,32'd-5166,32'd2213,32'd-369,32'd2558,32'd1186,32'd-2480,32'd-3369,32'd1412,32'd1511,32'd-374,32'd2252,32'd-1936,32'd1417,32'd2185,32'd2281,32'd2100,32'd-2763,32'd3266,32'd-1378,32'd5795,32'd669,32'd2087,32'd-6225,32'd4509,32'd-7172,32'd1838,32'd2265,32'd8686,32'd-697,32'd2810,32'd-1519,32'd896,32'd-1959,32'd4301,32'd1293,32'd-4401,32'd795,32'd1517,32'd-1816,32'd2558,32'd2431,32'd-5205,32'd4794,32'd-1856,32'd-142,32'd3796,32'd0,32'd6157,32'd-3420,32'd1505,32'd-689,32'd-4235,32'd-2841,32'd-1619,32'd-8105,32'd2180,32'd-5219,32'd2254,32'd1906,32'd-11250,32'd2929,32'd4326,32'd-2902,32'd-1417,32'd-5644,32'd1466,32'd-2100,32'd979,32'd5737,32'd-853,32'd1153,32'd5507,32'd965,32'd4089,32'd2174,32'd-2386,32'd-1314,32'd4670,32'd3818,32'd784,32'd-8466,32'd-4401,32'd621,32'd1439,32'd-18535,32'd-5083,32'd-3503,32'd-170,32'd-1322,32'd7700,32'd-8056,32'd-3576,32'd-1101,32'd1748,32'd-564,32'd4543,32'd604,32'd11074,32'd9902,32'd-6787,32'd-18,32'd-1212,32'd-1706,32'd668,32'd2897,32'd15322,32'd5009,32'd-497,32'd2316,32'd-7817,32'd1702,32'd9311,32'd7104,32'd-292,32'd12021,32'd-905,32'd-13789,32'd4409,32'd-8217,32'd-1016,32'd324,32'd622,32'd2069,32'd3452,32'd-10742,32'd1672,32'd9365,32'd14169,32'd-9326,32'd-5253,32'd2983,32'd-6499,32'd-1034,32'd-744,32'd-13974,32'd-4296,32'd-4125,32'd54,32'd9370,32'd3972,32'd-1364,32'd-2066,32'd2556,32'd3918,32'd5258,32'd-7700,32'd1523,32'd7875,32'd1634,32'd-1365,32'd-6166,32'd2165,32'd264,32'd8242,32'd1601,32'd-3779,32'd191,32'd-246,32'd2115,32'd-788,32'd14697,32'd290,32'd9428,32'd1017,32'd14160,32'd-12031,32'd3227,32'd303,32'd15966,32'd4047,32'd132,32'd-1667,32'd330,32'd3391,32'd-348,32'd8002,32'd1734,32'd-1440,32'd461,32'd-9589,32'd-17500,32'd-9775,32'd6142,32'd1041,32'd840,32'd4638,32'd-245,32'd3549,32'd-1680,32'd4116,32'd7539,32'd1976,32'd-3984,32'd374,32'd-1810,32'd-74,32'd1982,32'd-80,32'd3664,32'd1464,32'd436,32'd-2995,32'd568,32'd-385,32'd1872,32'd864,32'd4521,32'd2084,32'd-183,32'd-1182,32'd-4311,32'd-1064,32'd2312,32'd-1065,32'd-3486,32'd6123,32'd-7368,32'd-837,32'd-2905,32'd-2690,32'd2423,32'd-6020,32'd-3569,32'd2484,32'd-1656,32'd2442,32'd-1206,32'd-11435,32'd-6914,32'd-4252,32'd4465,32'd5439,32'd-1224,32'd2108,32'd-2159,32'd-914,32'd-8051,32'd2932,32'd2824,32'd-1196,32'd2163,32'd-1157,32'd-4025,32'd2070,32'd9814,32'd19,32'd4401,32'd6020,32'd-4216,32'd714,32'd15927,32'd-2346,32'd-1451,32'd-993,32'd3564,32'd-3364,32'd-1311,32'd6362,32'd8388,32'd-3608,32'd-8286,32'd4179,32'd2183,32'd969,32'd-6450,32'd4006,32'd2609,32'd1162,32'd-1800,32'd2211,32'd-835,32'd277,32'd-233,32'd6455,32'd2371,32'd5517,32'd2205,32'd13447,32'd1385,32'd-1392,32'd4458,32'd4582,32'd8466,32'd1472,32'd-2797,32'd243,32'd-6162,32'd7944,32'd12646,32'd-117,32'd4511,32'd2191,32'd2481,32'd-9970,32'd-5234,32'd-1815,32'd4680,32'd6596,32'd-9741,32'd662,32'd-14228,32'd1402,32'd-855,32'd5175,32'd-1238,32'd-128,32'd-1441,32'd2888,32'd-2749,32'd128,32'd-8339,32'd-1207,32'd-132,32'd-3300,32'd-3967,32'd10273,32'd-12509,32'd1939,32'd-4958,32'd-1072,32'd6430,32'd-2379,32'd-11464,32'd-2081,32'd-3679,32'd-3623,32'd3010,32'd269,32'd-7187,32'd1549,32'd-1353,32'd3881,32'd-663,32'd3811,32'd-1071,32'd-252,32'd-3684,32'd166,32'd7060,32'd-1794,32'd6611,32'd-2683,32'd-2373,32'd-1585,32'd-2058,32'd-423,32'd-4240,32'd-2406,32'd3996,32'd299,32'd-2274,32'd10947,32'd3583,32'd-8720,32'd1052,32'd450,32'd-11757,32'd5380,32'd-399,32'd-437,32'd-9355,32'd-3142,32'd-2578,32'd8129,32'd-1793,32'd-3837,32'd3083,32'd616,32'd-4980,32'd1093,32'd121,32'd3342,32'd235,32'd4396,32'd-9765,32'd-570,32'd6596,32'd7470,32'd7612,32'd180,32'd7841,32'd2067,32'd3090};
    Wx[57]='{32'd-2132,32'd-4680,32'd71,32'd863,32'd760,32'd9,32'd841,32'd1237,32'd-1582,32'd-282,32'd-8784,32'd-1182,32'd2602,32'd-1617,32'd7524,32'd-7084,32'd-1363,32'd-3073,32'd-2213,32'd-3540,32'd-2166,32'd3894,32'd841,32'd-3566,32'd1799,32'd1828,32'd-2624,32'd-2138,32'd-6206,32'd3410,32'd397,32'd-4047,32'd141,32'd-1872,32'd1202,32'd3222,32'd-848,32'd6240,32'd2446,32'd230,32'd-1715,32'd-675,32'd1948,32'd1481,32'd-2115,32'd188,32'd9819,32'd2447,32'd-1155,32'd-1561,32'd-1076,32'd2188,32'd-1313,32'd3957,32'd-715,32'd744,32'd-2316,32'd-5009,32'd2255,32'd-1639,32'd-3889,32'd-5458,32'd8354,32'd-2426,32'd-4421,32'd-1462,32'd-1939,32'd-8276,32'd-2164,32'd1162,32'd1622,32'd-1685,32'd-3093,32'd5205,32'd581,32'd3518,32'd-2080,32'd187,32'd3496,32'd452,32'd-1795,32'd-867,32'd1250,32'd-3049,32'd-2817,32'd-6660,32'd1405,32'd-1596,32'd-946,32'd-727,32'd2915,32'd1910,32'd761,32'd-5708,32'd-8583,32'd-300,32'd2089,32'd617,32'd-2958,32'd3002,32'd287,32'd-5600,32'd722,32'd4707,32'd-3686,32'd-411,32'd-9067,32'd-7309,32'd-181,32'd1767,32'd10029,32'd1340,32'd-3310,32'd9926,32'd-10771,32'd-4101,32'd-3701,32'd2432,32'd-285,32'd-2617,32'd-723,32'd3889,32'd-5214,32'd-1320,32'd1470,32'd-3415,32'd3203,32'd2156,32'd-4096,32'd-13593,32'd4667,32'd4858,32'd-4018,32'd3427,32'd-4604,32'd4045,32'd-3554,32'd2922,32'd-9570,32'd-1571,32'd6635,32'd-6586,32'd-1555,32'd7109,32'd-3254,32'd2495,32'd-2335,32'd-4516,32'd-6313,32'd-688,32'd14189,32'd-7788,32'd1756,32'd4499,32'd1499,32'd16035,32'd-10419,32'd2534,32'd-1796,32'd-897,32'd5034,32'd-4841,32'd-6284,32'd-932,32'd6806,32'd63,32'd5195,32'd-5346,32'd-1274,32'd-959,32'd196,32'd-4479,32'd2156,32'd-14902,32'd559,32'd-4357,32'd-7353,32'd-2185,32'd4401,32'd-526,32'd4033,32'd-12216,32'd-5468,32'd-4350,32'd915,32'd10146,32'd-1639,32'd7880,32'd-4848,32'd1860,32'd-3591,32'd-3408,32'd-6464,32'd-1324,32'd-4841,32'd2758,32'd3725,32'd12578,32'd-781,32'd-8754,32'd-484,32'd-8906,32'd-2536,32'd-6489,32'd-1416,32'd704,32'd-1998,32'd3957,32'd2841,32'd-1276,32'd-3498,32'd10,32'd3015,32'd-6518,32'd-295,32'd220,32'd-1596,32'd-3764,32'd1748,32'd2108,32'd-443,32'd-2775,32'd955,32'd-2949,32'd-5454,32'd-86,32'd2147,32'd625,32'd10908,32'd-3479,32'd1291,32'd3801,32'd-1173,32'd1483,32'd-4064,32'd13,32'd2702,32'd5419,32'd3830,32'd-3295,32'd3908,32'd-2829,32'd689,32'd-2058,32'd8022,32'd4238,32'd8598,32'd-667,32'd-3049,32'd-5854,32'd-3100,32'd33,32'd-704,32'd1751,32'd-1145,32'd276,32'd-3981,32'd-4233,32'd-5551,32'd-273,32'd911,32'd-691,32'd-2465,32'd4216,32'd-662,32'd3000,32'd3854,32'd34,32'd-332,32'd2420,32'd-3747,32'd3505,32'd-10224,32'd-7119,32'd-903,32'd1180,32'd10244,32'd-4797,32'd2563,32'd363,32'd2038,32'd1787,32'd-2183,32'd7187,32'd134,32'd-5136,32'd1077,32'd1417,32'd-1859,32'd-980,32'd41,32'd-4506,32'd-7421,32'd-3684,32'd-9799,32'd-4484,32'd2617,32'd-3215,32'd150,32'd-6142,32'd-30,32'd3610,32'd7568,32'd2580,32'd-2714,32'd-1405,32'd-683,32'd-3525,32'd-4809,32'd304,32'd-14677,32'd4440,32'd4389,32'd2524,32'd4958,32'd-5014,32'd2546,32'd-681,32'd4455,32'd-6669,32'd867,32'd-2418,32'd3405,32'd-690,32'd-2106,32'd-4409,32'd2849,32'd-2749,32'd1148,32'd5732,32'd845,32'd1154,32'd8925,32'd2866,32'd6630,32'd1593,32'd-1557,32'd1870,32'd4360,32'd-3701,32'd4755,32'd-1383,32'd-4111,32'd9521,32'd5981,32'd4125,32'd-9326,32'd-5073,32'd2927,32'd-115,32'd11240,32'd257,32'd2208,32'd5991,32'd-556,32'd-1110,32'd-5551,32'd-4689,32'd-1036,32'd919,32'd1885,32'd-1324,32'd553,32'd-212,32'd386,32'd4453,32'd1507,32'd-254,32'd811,32'd-3918,32'd1248,32'd-3740,32'd-9614,32'd-3129,32'd-762,32'd-3864,32'd1975,32'd135,32'd6337,32'd66,32'd-296,32'd8486,32'd-679,32'd10693,32'd-2932,32'd-3232,32'd-1678,32'd8491,32'd375,32'd700,32'd3320,32'd6352,32'd-7006,32'd-5278,32'd345,32'd-336,32'd3195,32'd-8422,32'd-5336,32'd2863};
    Wx[58]='{32'd-912,32'd-7055,32'd1208,32'd-1329,32'd-1910,32'd-1749,32'd4938,32'd4689,32'd-2121,32'd3974,32'd-1154,32'd4016,32'd3452,32'd1095,32'd3041,32'd2116,32'd-1583,32'd2152,32'd4072,32'd1871,32'd-1608,32'd2563,32'd-78,32'd-804,32'd-2580,32'd2548,32'd2124,32'd953,32'd739,32'd-3046,32'd-3666,32'd2408,32'd-1912,32'd661,32'd-791,32'd1536,32'd-3269,32'd4133,32'd6,32'd-1420,32'd4560,32'd148,32'd1138,32'd1080,32'd9257,32'd2927,32'd1479,32'd3549,32'd4565,32'd-606,32'd8432,32'd4882,32'd700,32'd1577,32'd-355,32'd65,32'd4348,32'd4665,32'd3300,32'd3166,32'd-2402,32'd352,32'd9697,32'd2301,32'd2259,32'd2143,32'd-813,32'd7294,32'd-685,32'd-471,32'd517,32'd-2631,32'd-2352,32'd-247,32'd-314,32'd446,32'd3586,32'd-2980,32'd273,32'd3508,32'd2023,32'd272,32'd1998,32'd-263,32'd-5102,32'd3366,32'd-1838,32'd-424,32'd-359,32'd5375,32'd1281,32'd2276,32'd4316,32'd-3684,32'd-330,32'd1538,32'd-1716,32'd-4279,32'd858,32'd2128,32'd-1436,32'd-136,32'd1391,32'd-336,32'd3395,32'd-41,32'd-6616,32'd7553,32'd3630,32'd715,32'd-1190,32'd-1246,32'd2619,32'd6479,32'd2229,32'd6821,32'd-11259,32'd-3388,32'd164,32'd-1380,32'd-143,32'd5039,32'd3320,32'd8310,32'd4526,32'd2807,32'd7802,32'd821,32'd-5327,32'd-3710,32'd6728,32'd-1091,32'd-5229,32'd5043,32'd-746,32'd13085,32'd-4797,32'd1871,32'd-15810,32'd3835,32'd442,32'd9379,32'd9013,32'd13740,32'd27832,32'd-13037,32'd11728,32'd5136,32'd2900,32'd-2841,32'd1441,32'd-15244,32'd1929,32'd-258,32'd-5400,32'd4152,32'd-2365,32'd-4108,32'd6015,32'd4765,32'd2805,32'd13925,32'd-5366,32'd5131,32'd-240,32'd869,32'd526,32'd11093,32'd5004,32'd-1898,32'd-5937,32'd-7978,32'd-2033,32'd-1712,32'd1995,32'd-5249,32'd1235,32'd-7690,32'd-11064,32'd3276,32'd-7485,32'd-5527,32'd-14453,32'd-3569,32'd-2080,32'd4165,32'd2932,32'd3449,32'd-1986,32'd6123,32'd-591,32'd-14013,32'd-8608,32'd-2578,32'd-7666,32'd7265,32'd2333,32'd-5419,32'd2110,32'd10351,32'd661,32'd-7436,32'd1770,32'd1469,32'd80,32'd-1645,32'd2080,32'd-3906,32'd2531,32'd2436,32'd-864,32'd-207,32'd-2575,32'd-6064,32'd1078,32'd-7773,32'd2156,32'd-1207,32'd2198,32'd6147,32'd-1468,32'd-2331,32'd78,32'd-1608,32'd-223,32'd-3002,32'd-602,32'd1267,32'd1463,32'd2922,32'd13,32'd-4362,32'd-5390,32'd-2536,32'd-1485,32'd6713,32'd-1850,32'd2592,32'd-5639,32'd-5107,32'd-4660,32'd-8969,32'd-2033,32'd6254,32'd-3291,32'd-1705,32'd-14853,32'd-6054,32'd-1126,32'd-4497,32'd-7534,32'd-6538,32'd2172,32'd-1511,32'd1715,32'd-3403,32'd-3652,32'd2360,32'd954,32'd-7270,32'd2902,32'd-2978,32'd-3947,32'd-85,32'd4106,32'd3759,32'd-4230,32'd-6669,32'd-3085,32'd-6616,32'd2517,32'd-406,32'd-6196,32'd-3366,32'd-650,32'd-3945,32'd-8066,32'd-4616,32'd3979,32'd305,32'd-2216,32'd-1638,32'd-4399,32'd-5092,32'd-3037,32'd950,32'd404,32'd-1203,32'd725,32'd2966,32'd6674,32'd-1453,32'd-5776,32'd-8110,32'd1873,32'd-116,32'd-549,32'd-6606,32'd5800,32'd-1791,32'd-1142,32'd1888,32'd-1260,32'd-5747,32'd-1232,32'd-1846,32'd9257,32'd-6210,32'd-1120,32'd7597,32'd2983,32'd6445,32'd5048,32'd-506,32'd444,32'd-4826,32'd8886,32'd4580,32'd9912,32'd7065,32'd-8432,32'd-6894,32'd462,32'd4228,32'd-6235,32'd-1430,32'd1192,32'd-8198,32'd5825,32'd4523,32'd-712,32'd-3571,32'd-5385,32'd-3735,32'd1986,32'd4960,32'd-5922,32'd-4670,32'd-14101,32'd-2656,32'd4626,32'd-2553,32'd-2656,32'd5483,32'd-3974,32'd1904,32'd-2695,32'd4279,32'd-8178,32'd-167,32'd6416,32'd2128,32'd-6254,32'd-6547,32'd-661,32'd-4355,32'd-7167,32'd3312,32'd-195,32'd1787,32'd3234,32'd3715,32'd-2069,32'd3181,32'd-508,32'd-8198,32'd1329,32'd-5620,32'd-3352,32'd-1872,32'd-1717,32'd532,32'd-54,32'd-1726,32'd3513,32'd-2392,32'd-3789,32'd1163,32'd3303,32'd5166,32'd-728,32'd2531,32'd1906,32'd1661,32'd-7216,32'd-5507,32'd-32,32'd3237,32'd1248,32'd6909,32'd11269,32'd-2087,32'd-1956,32'd12324,32'd-3339,32'd-6025,32'd-8471,32'd-1613,32'd2058,32'd3081};
    Wx[59]='{32'd-1990,32'd-8383,32'd-4753,32'd682,32'd296,32'd398,32'd2171,32'd-2347,32'd-740,32'd2670,32'd-1413,32'd858,32'd-2491,32'd245,32'd1243,32'd-4548,32'd11953,32'd4902,32'd3640,32'd-1254,32'd746,32'd-1566,32'd-2680,32'd-2086,32'd-2449,32'd-962,32'd2517,32'd1026,32'd-2141,32'd-3566,32'd-2409,32'd-5761,32'd536,32'd-3962,32'd-8164,32'd4135,32'd-2154,32'd-3383,32'd-3225,32'd-198,32'd-2475,32'd-9570,32'd-4570,32'd289,32'd138,32'd-2476,32'd-4335,32'd3100,32'd-1300,32'd-1396,32'd-2651,32'd-1649,32'd-181,32'd-1169,32'd-3781,32'd-5854,32'd-3552,32'd5000,32'd1680,32'd-3034,32'd-7763,32'd8759,32'd-3413,32'd-2033,32'd-875,32'd5234,32'd132,32'd-7055,32'd-1353,32'd3532,32'd20,32'd-9931,32'd727,32'd-7329,32'd-78,32'd-2083,32'd5532,32'd-449,32'd731,32'd2215,32'd5986,32'd-1239,32'd1407,32'd-4453,32'd-1506,32'd318,32'd-662,32'd-2673,32'd-34,32'd-2895,32'd913,32'd-4702,32'd-1833,32'd4013,32'd-2459,32'd-3811,32'd1741,32'd-5229,32'd7143,32'd-759,32'd-3547,32'd10625,32'd3166,32'd5522,32'd7597,32'd455,32'd-4047,32'd-996,32'd3430,32'd-2424,32'd-9702,32'd-6982,32'd2700,32'd12216,32'd1210,32'd9765,32'd845,32'd-6801,32'd2038,32'd-4663,32'd1220,32'd-5747,32'd1262,32'd4274,32'd-5971,32'd-2775,32'd5820,32'd4907,32'd-10498,32'd-3229,32'd-3212,32'd-618,32'd4155,32'd-10781,32'd-2229,32'd2595,32'd-4055,32'd2648,32'd-4299,32'd-1560,32'd-3750,32'd5273,32'd-10332,32'd13095,32'd1665,32'd569,32'd692,32'd4675,32'd823,32'd-9570,32'd-3508,32'd-7299,32'd-10224,32'd3408,32'd-7124,32'd-8,32'd7851,32'd368,32'd2565,32'd-3964,32'd-617,32'd4670,32'd9775,32'd-5317,32'd-2430,32'd-4140,32'd-2036,32'd1307,32'd5922,32'd735,32'd-1124,32'd-9936,32'd-6352,32'd6923,32'd-759,32'd11201,32'd13144,32'd10927,32'd5566,32'd-1816,32'd9726,32'd4433,32'd-8046,32'd-13964,32'd-8886,32'd-5556,32'd2924,32'd-2729,32'd-5244,32'd-253,32'd-10810,32'd4936,32'd-8574,32'd2233,32'd16767,32'd-6582,32'd4694,32'd431,32'd6347,32'd-8676,32'd-1087,32'd1942,32'd-2824,32'd5302,32'd-394,32'd1376,32'd8398,32'd2197,32'd351,32'd10107,32'd5776,32'd2117,32'd-2343,32'd3544,32'd5122,32'd61,32'd-4033,32'd7236,32'd-1268,32'd-363,32'd1671,32'd35,32'd-3188,32'd-7133,32'd-29,32'd2268,32'd-2741,32'd3449,32'd4699,32'd-10039,32'd-507,32'd5971,32'd4187,32'd9116,32'd2408,32'd1588,32'd-3078,32'd-1490,32'd-827,32'd2890,32'd-1079,32'd-3183,32'd5844,32'd449,32'd38,32'd-1134,32'd-4655,32'd461,32'd-8037,32'd2196,32'd-9702,32'd4206,32'd2727,32'd6230,32'd3364,32'd2583,32'd2493,32'd809,32'd2988,32'd6376,32'd720,32'd-3525,32'd4194,32'd-2380,32'd-6503,32'd3269,32'd358,32'd1291,32'd834,32'd4206,32'd-31,32'd7363,32'd-3110,32'd-2746,32'd-1654,32'd-3869,32'd1232,32'd-1237,32'd7939,32'd232,32'd-933,32'd-6513,32'd-621,32'd1071,32'd-7934,32'd5405,32'd-5673,32'd2783,32'd1102,32'd-22,32'd-2768,32'd-4902,32'd4865,32'd1470,32'd9809,32'd6230,32'd-1951,32'd-542,32'd1413,32'd7807,32'd-7250,32'd944,32'd1452,32'd1013,32'd-3300,32'd-6127,32'd12871,32'd-2062,32'd1611,32'd7001,32'd-2089,32'd3061,32'd-7348,32'd11826,32'd-2127,32'd4221,32'd8881,32'd7333,32'd11572,32'd-939,32'd-1484,32'd-678,32'd-2474,32'd-1507,32'd-9633,32'd2607,32'd4296,32'd1064,32'd-761,32'd-287,32'd3105,32'd-1501,32'd-4309,32'd3676,32'd-5009,32'd1264,32'd3464,32'd-1050,32'd-2998,32'd8041,32'd3708,32'd1806,32'd-462,32'd9204,32'd-755,32'd7241,32'd1461,32'd9370,32'd-9550,32'd-1945,32'd6362,32'd5878,32'd3547,32'd1893,32'd7998,32'd1579,32'd899,32'd-4755,32'd5712,32'd569,32'd-3403,32'd5693,32'd-2680,32'd827,32'd-2692,32'd-4545,32'd11318,32'd399,32'd-5781,32'd5927,32'd471,32'd3605,32'd2592,32'd-989,32'd12031,32'd-2454,32'd-2072,32'd3674,32'd-1779,32'd-154,32'd3059,32'd9252,32'd5864,32'd1138,32'd-11357,32'd-1614,32'd-4072,32'd2312,32'd-5585,32'd967,32'd-141,32'd-4123,32'd-5131,32'd14951,32'd-698,32'd-723,32'd476,32'd3933,32'd4318,32'd7216};
    Wx[60]='{32'd784,32'd-1481,32'd2177,32'd1282,32'd-458,32'd-2575,32'd-1320,32'd-2836,32'd4060,32'd3269,32'd5385,32'd807,32'd-2496,32'd6435,32'd-3925,32'd1126,32'd-6489,32'd242,32'd1693,32'd545,32'd489,32'd-3681,32'd-5859,32'd1672,32'd-2272,32'd-1125,32'd1768,32'd193,32'd1824,32'd1054,32'd-2156,32'd-2369,32'd1262,32'd-141,32'd-1932,32'd1982,32'd-2700,32'd1755,32'd-2073,32'd-2220,32'd-1842,32'd-3225,32'd-3327,32'd1231,32'd-1827,32'd2583,32'd2270,32'd-480,32'd938,32'd-1405,32'd-1033,32'd-4113,32'd-5141,32'd-4030,32'd5341,32'd-2264,32'd-1006,32'd5937,32'd-2073,32'd-5800,32'd3850,32'd-1063,32'd-8945,32'd-142,32'd-676,32'd3415,32'd-367,32'd-3957,32'd-46,32'd1555,32'd-4030,32'd-7656,32'd1245,32'd-1298,32'd-736,32'd-1010,32'd-1373,32'd-4025,32'd-4855,32'd-3796,32'd-510,32'd555,32'd-5810,32'd-2031,32'd-3110,32'd-9648,32'd-3125,32'd3051,32'd1345,32'd3293,32'd-2233,32'd1921,32'd-2390,32'd-4138,32'd-6391,32'd-2305,32'd-2442,32'd-4182,32'd3945,32'd-3911,32'd-1043,32'd13798,32'd-3088,32'd-3403,32'd-1001,32'd4990,32'd5297,32'd1369,32'd-2467,32'd811,32'd430,32'd7275,32'd-721,32'd7475,32'd9565,32'd11406,32'd-3757,32'd4108,32'd-1271,32'd1878,32'd-1121,32'd-1892,32'd-423,32'd9770,32'd4313,32'd-5131,32'd-2358,32'd-1483,32'd-1842,32'd-4357,32'd7026,32'd-10654,32'd-32,32'd1593,32'd-4943,32'd-2109,32'd5146,32'd-387,32'd-2326,32'd8413,32'd-4130,32'd20625,32'd-1213,32'd4570,32'd11386,32'd-13115,32'd4584,32'd6875,32'd-6455,32'd1547,32'd-7353,32'd835,32'd5180,32'd-6538,32'd-3989,32'd-7177,32'd-789,32'd-3757,32'd6528,32'd6342,32'd-181,32'd5039,32'd-18603,32'd-4582,32'd10468,32'd1412,32'd-2805,32'd-12275,32'd698,32'd-2851,32'd7299,32'd1683,32'd-5131,32'd4509,32'd60,32'd14960,32'd4440,32'd-1754,32'd-7104,32'd-883,32'd-1618,32'd5024,32'd8378,32'd12636,32'd-5234,32'd-3024,32'd2421,32'd4438,32'd-646,32'd-1778,32'd-3586,32'd-10195,32'd401,32'd-99,32'd22539,32'd-6572,32'd-4318,32'd9750,32'd7333,32'd-12861,32'd-822,32'd6323,32'd4353,32'd1749,32'd99,32'd-2370,32'd5175,32'd5595,32'd-8076,32'd2141,32'd5683,32'd-2418,32'd367,32'd8173,32'd-4301,32'd5639,32'd-200,32'd7470,32'd1243,32'd-80,32'd4614,32'd57,32'd-2081,32'd1090,32'd811,32'd-354,32'd-2476,32'd1157,32'd1815,32'd3024,32'd-3244,32'd1210,32'd-673,32'd3647,32'd-2565,32'd1801,32'd-5288,32'd-1694,32'd10917,32'd6542,32'd1966,32'd2052,32'd2041,32'd-2846,32'd3269,32'd1917,32'd-13671,32'd-7353,32'd2442,32'd2917,32'd3686,32'd1455,32'd-639,32'd773,32'd2561,32'd-2322,32'd897,32'd4670,32'd-6308,32'd5976,32'd4250,32'd3662,32'd2546,32'd5610,32'd-1434,32'd921,32'd-968,32'd-125,32'd3498,32'd817,32'd4572,32'd2448,32'd3771,32'd4645,32'd-2492,32'd9116,32'd8354,32'd1872,32'd1885,32'd-8227,32'd-4633,32'd279,32'd447,32'd-2154,32'd-3195,32'd4609,32'd-3215,32'd-4523,32'd-5312,32'd-1357,32'd-4294,32'd7460,32'd9633,32'd-3786,32'd7602,32'd1342,32'd-1757,32'd-778,32'd-393,32'd-1990,32'd-2070,32'd-5942,32'd3295,32'd115,32'd-1745,32'd-12255,32'd2524,32'd-4555,32'd3344,32'd5156,32'd11005,32'd-1014,32'd898,32'd3637,32'd-1719,32'd5581,32'd1043,32'd3837,32'd-12294,32'd498,32'd-3098,32'd-2086,32'd-7622,32'd4348,32'd-2363,32'd3208,32'd3022,32'd3583,32'd-2915,32'd892,32'd-1160,32'd-5151,32'd-11425,32'd-29,32'd5605,32'd5317,32'd1777,32'd-1497,32'd-3852,32'd2678,32'd976,32'd4880,32'd931,32'd6640,32'd1203,32'd4567,32'd-1152,32'd-1337,32'd-13408,32'd-132,32'd4333,32'd3471,32'd-6191,32'd-3837,32'd4938,32'd10244,32'd-3093,32'd10087,32'd-1105,32'd651,32'd-661,32'd-3298,32'd-2137,32'd7890,32'd1304,32'd-1781,32'd-2766,32'd3215,32'd-507,32'd-7006,32'd-5639,32'd-128,32'd901,32'd2851,32'd-86,32'd2514,32'd2541,32'd-92,32'd827,32'd-2420,32'd1095,32'd6889,32'd2447,32'd-8579,32'd-7485,32'd774,32'd-2108,32'd-457,32'd458,32'd1088,32'd1981,32'd4570,32'd1212,32'd-2846,32'd-3798,32'd83,32'd-8168,32'd2802,32'd5888,32'd-3779};
    Wx[61]='{32'd1846,32'd-3222,32'd1066,32'd1682,32'd-1350,32'd972,32'd-3073,32'd-2454,32'd-8085,32'd1235,32'd1353,32'd-765,32'd-603,32'd-2304,32'd-584,32'd4721,32'd3012,32'd-1729,32'd-4743,32'd1927,32'd585,32'd-924,32'd-1295,32'd-4272,32'd1904,32'd-315,32'd-3056,32'd2761,32'd330,32'd3598,32'd4794,32'd-5439,32'd4309,32'd805,32'd2656,32'd-991,32'd544,32'd-2512,32'd5668,32'd4704,32'd2105,32'd3227,32'd3608,32'd-465,32'd7553,32'd2695,32'd-5473,32'd1574,32'd-4375,32'd937,32'd-2235,32'd-2066,32'd1782,32'd5053,32'd-520,32'd567,32'd3500,32'd2320,32'd-115,32'd-54,32'd-2832,32'd186,32'd-575,32'd1050,32'd2683,32'd-2888,32'd-2369,32'd1392,32'd989,32'd299,32'd-1927,32'd8598,32'd-5800,32'd996,32'd-1467,32'd-5405,32'd2438,32'd407,32'd75,32'd-2575,32'd-2030,32'd-7416,32'd2243,32'd-3254,32'd-1289,32'd-2800,32'd288,32'd3728,32'd-1021,32'd-1001,32'd-1013,32'd-1273,32'd158,32'd1520,32'd809,32'd11,32'd2113,32'd7929,32'd419,32'd-88,32'd-2980,32'd11718,32'd-2291,32'd1051,32'd-3388,32'd-200,32'd-5766,32'd-12001,32'd841,32'd-834,32'd12636,32'd1801,32'd5898,32'd7299,32'd1102,32'd4006,32'd9101,32'd2015,32'd2225,32'd3701,32'd-989,32'd5410,32'd-3291,32'd2663,32'd-5981,32'd4072,32'd-900,32'd-9106,32'd7988,32'd-7031,32'd1610,32'd-6196,32'd1429,32'd5800,32'd-680,32'd-2335,32'd1160,32'd3049,32'd-11621,32'd1160,32'd-4372,32'd-8427,32'd-6420,32'd-13007,32'd1416,32'd673,32'd-6674,32'd4160,32'd-2171,32'd-10908,32'd15498,32'd-495,32'd7329,32'd1501,32'd227,32'd975,32'd9858,32'd2199,32'd-1461,32'd-7509,32'd1165,32'd4636,32'd1817,32'd-3139,32'd6865,32'd-2932,32'd-1090,32'd5932,32'd-466,32'd847,32'd-6782,32'd-6962,32'd284,32'd-18818,32'd-3815,32'd-17041,32'd-8554,32'd4641,32'd328,32'd-3127,32'd-3671,32'd9809,32'd2888,32'd3342,32'd-2692,32'd5952,32'd-1159,32'd10644,32'd3610,32'd-1656,32'd-1253,32'd6381,32'd-14404,32'd-1735,32'd-6362,32'd4836,32'd-2481,32'd-1807,32'd950,32'd9946,32'd310,32'd-7299,32'd170,32'd-5029,32'd-2093,32'd-1106,32'd856,32'd-4174,32'd-1915,32'd-4333,32'd-4033,32'd1607,32'd-2839,32'd-4992,32'd-2517,32'd-9370,32'd3378,32'd-7729,32'd-4272,32'd1624,32'd1566,32'd813,32'd-1844,32'd-7719,32'd-5419,32'd-4406,32'd-3549,32'd-379,32'd-11523,32'd298,32'd-930,32'd-6455,32'd-1474,32'd-8325,32'd1055,32'd-3515,32'd-5234,32'd812,32'd-5458,32'd-3137,32'd-4780,32'd11210,32'd-8945,32'd3522,32'd-734,32'd-1596,32'd-1873,32'd-3500,32'd640,32'd-2912,32'd-11582,32'd-1895,32'd-2,32'd-2880,32'd-6088,32'd932,32'd-5112,32'd-4514,32'd3381,32'd-5361,32'd-9,32'd-5717,32'd-4091,32'd-4128,32'd-11503,32'd-3928,32'd-148,32'd-4082,32'd-306,32'd-1832,32'd-2580,32'd7968,32'd-1373,32'd-4824,32'd-3979,32'd-11416,32'd-657,32'd-6538,32'd-6772,32'd-1751,32'd-3291,32'd56,32'd-276,32'd-1013,32'd1633,32'd-3789,32'd-1839,32'd-5151,32'd1667,32'd-902,32'd5825,32'd-679,32'd-11494,32'd1170,32'd-1846,32'd858,32'd-1254,32'd-10781,32'd-5058,32'd-2700,32'd7998,32'd-575,32'd-4431,32'd-3850,32'd-6054,32'd-438,32'd-4738,32'd9838,32'd758,32'd-138,32'd-2401,32'd-3122,32'd4636,32'd-211,32'd-2670,32'd2416,32'd1899,32'd2102,32'd-5112,32'd2338,32'd3447,32'd-257,32'd3918,32'd-1943,32'd1220,32'd-684,32'd-6323,32'd3808,32'd2423,32'd-106,32'd4765,32'd434,32'd-336,32'd-136,32'd-1373,32'd-4816,32'd2773,32'd2722,32'd-706,32'd913,32'd-4533,32'd1943,32'd9985,32'd5498,32'd708,32'd910,32'd1091,32'd-3684,32'd-7182,32'd526,32'd-1524,32'd-11035,32'd386,32'd-269,32'd-4392,32'd3767,32'd-3635,32'd-8779,32'd20,32'd2305,32'd-3408,32'd-834,32'd-1070,32'd7231,32'd-779,32'd-14443,32'd-3127,32'd205,32'd-3549,32'd-1497,32'd1154,32'd5454,32'd-4885,32'd-9291,32'd-4763,32'd-7431,32'd4689,32'd-5981,32'd-1280,32'd-793,32'd-4897,32'd-4523,32'd-6503,32'd-4746,32'd-5463,32'd6113,32'd-272,32'd-1512,32'd-879,32'd-4372,32'd-3928,32'd149,32'd-8095,32'd8725,32'd3771,32'd-1857,32'd-786,32'd-8662,32'd-3940,32'd-163};
    Wx[62]='{32'd1567,32'd6640,32'd-4350,32'd-4843,32'd932,32'd1246,32'd3288,32'd-3261,32'd1307,32'd729,32'd429,32'd-1517,32'd737,32'd-4445,32'd3046,32'd-3073,32'd-1122,32'd1180,32'd545,32'd2418,32'd704,32'd1232,32'd-3110,32'd-2263,32'd-1026,32'd-961,32'd793,32'd225,32'd3203,32'd-794,32'd681,32'd-1866,32'd3020,32'd2983,32'd-803,32'd-4836,32'd-718,32'd-1904,32'd-3825,32'd-2414,32'd260,32'd2683,32'd5532,32'd-2658,32'd-2978,32'd-1303,32'd-7412,32'd-4294,32'd-6923,32'd-3056,32'd-4753,32'd7822,32'd1441,32'd520,32'd363,32'd-5175,32'd-7216,32'd1184,32'd2565,32'd-1724,32'd-2366,32'd-59,32'd-1655,32'd-1643,32'd2758,32'd1690,32'd3310,32'd-2379,32'd-4467,32'd-984,32'd1885,32'd-7622,32'd-1634,32'd6074,32'd87,32'd-188,32'd-12255,32'd-1319,32'd-2451,32'd-4621,32'd-975,32'd-13466,32'd-3395,32'd-5708,32'd5449,32'd3764,32'd2020,32'd-1414,32'd-623,32'd1920,32'd1390,32'd-623,32'd-1547,32'd-1353,32'd-2702,32'd1740,32'd1585,32'd-667,32'd-6396,32'd70,32'd4995,32'd15273,32'd3959,32'd-3007,32'd-1268,32'd-1975,32'd-5019,32'd11210,32'd3349,32'd-47,32'd536,32'd-4113,32'd246,32'd12792,32'd842,32'd-1555,32'd20761,32'd2509,32'd-3178,32'd456,32'd-2073,32'd-6049,32'd10185,32'd-2304,32'd955,32'd-2318,32'd-3315,32'd-4589,32'd17871,32'd-1923,32'd2277,32'd-1422,32'd3474,32'd-1635,32'd653,32'd381,32'd3571,32'd-11025,32'd1762,32'd4565,32'd15751,32'd-1473,32'd5039,32'd-794,32'd8750,32'd3981,32'd-4626,32'd-3444,32'd1613,32'd11992,32'd2312,32'd14384,32'd19033,32'd2770,32'd6240,32'd-642,32'd13388,32'd-307,32'd9541,32'd-2106,32'd4155,32'd-2077,32'd-3076,32'd-332,32'd880,32'd4792,32'd-1414,32'd-11513,32'd-4389,32'd-1447,32'd-7636,32'd440,32'd-3327,32'd426,32'd4165,32'd-12939,32'd-9780,32'd1033,32'd-19765,32'd-5136,32'd3105,32'd10097,32'd-7895,32'd1474,32'd2846,32'd1756,32'd368,32'd-9287,32'd-810,32'd2403,32'd-789,32'd394,32'd-14121,32'd-1137,32'd-8627,32'd-10566,32'd1909,32'd-7675,32'd-4265,32'd-17519,32'd4499,32'd3356,32'd-1596,32'd-4807,32'd-757,32'd2302,32'd4770,32'd4016,32'd397,32'd-2944,32'd-9008,32'd5942,32'd-1939,32'd-1499,32'd-5541,32'd2277,32'd1285,32'd-1035,32'd1049,32'd303,32'd513,32'd-578,32'd561,32'd-4614,32'd-3117,32'd-1494,32'd-6953,32'd2111,32'd3571,32'd-3942,32'd-5024,32'd-8144,32'd9418,32'd3198,32'd-3862,32'd-4453,32'd2229,32'd288,32'd787,32'd700,32'd991,32'd-7968,32'd-1582,32'd-543,32'd1182,32'd1865,32'd7788,32'd-6513,32'd2697,32'd-661,32'd1484,32'd-2188,32'd5107,32'd-1287,32'd-1862,32'd2895,32'd6215,32'd3666,32'd-12519,32'd-243,32'd-4621,32'd-4411,32'd-2239,32'd-7407,32'd1831,32'd-1398,32'd2976,32'd338,32'd-3291,32'd971,32'd-5278,32'd-1354,32'd905,32'd-3378,32'd1644,32'd839,32'd-3828,32'd2954,32'd-1551,32'd-6635,32'd590,32'd152,32'd4545,32'd2539,32'd-654,32'd-4846,32'd-320,32'd-111,32'd-1589,32'd4750,32'd6347,32'd3798,32'd-1212,32'd1994,32'd424,32'd-227,32'd-3256,32'd1730,32'd5083,32'd1845,32'd3352,32'd2687,32'd-7822,32'd-1378,32'd-5078,32'd9716,32'd1137,32'd-4584,32'd-3098,32'd-797,32'd-15390,32'd131,32'd808,32'd-8266,32'd3728,32'd-1967,32'd-256,32'd-4970,32'd-3879,32'd-14394,32'd-627,32'd223,32'd-5703,32'd-5776,32'd-272,32'd-1263,32'd-3115,32'd5288,32'd-1790,32'd-2521,32'd-4821,32'd-14140,32'd3510,32'd-1413,32'd-1779,32'd-6821,32'd-2314,32'd7475,32'd-1807,32'd-1807,32'd-3198,32'd-11210,32'd-2729,32'd552,32'd-2810,32'd-3579,32'd-1685,32'd-9125,32'd142,32'd1932,32'd-1549,32'd235,32'd-3388,32'd-1965,32'd-4633,32'd-8154,32'd-2469,32'd-2059,32'd-9130,32'd-4602,32'd1778,32'd-6948,32'd-2155,32'd-457,32'd1871,32'd5722,32'd3999,32'd-1280,32'd5786,32'd-8916,32'd-4987,32'd-12021,32'd802,32'd-7412,32'd-71,32'd-2700,32'd-12177,32'd-12314,32'd-648,32'd-3427,32'd1063,32'd-8066,32'd-11113,32'd2983,32'd5302,32'd-5229,32'd393,32'd-2929,32'd4523,32'd1016,32'd3598,32'd2468,32'd-3251,32'd2346,32'd-596,32'd4211,32'd3759,32'd5375,32'd-1552,32'd-2939};
    Wx[63]='{32'd1256,32'd2656,32'd51,32'd-3034,32'd2639,32'd3413,32'd-2587,32'd2415,32'd-919,32'd-751,32'd2502,32'd-1591,32'd32,32'd-1087,32'd-1894,32'd-278,32'd-4631,32'd-505,32'd-1406,32'd-996,32'd-3186,32'd-4201,32'd-3618,32'd-6215,32'd-832,32'd-5556,32'd1789,32'd-944,32'd-1595,32'd153,32'd750,32'd-5537,32'd-3420,32'd-1408,32'd2348,32'd-588,32'd1052,32'd-3847,32'd-1865,32'd1892,32'd-1605,32'd1119,32'd-2188,32'd-1385,32'd-1496,32'd2303,32'd-7924,32'd95,32'd-5361,32'd553,32'd-7939,32'd1402,32'd-3061,32'd1579,32'd1096,32'd2673,32'd-962,32'd-957,32'd2077,32'd-6713,32'd-821,32'd3002,32'd-6757,32'd-3459,32'd-4890,32'd-3610,32'd-2819,32'd2568,32'd-451,32'd1069,32'd-567,32'd-798,32'd4345,32'd-1708,32'd1216,32'd-2995,32'd-6933,32'd-971,32'd-901,32'd-972,32'd1320,32'd-3369,32'd-3823,32'd-2739,32'd2648,32'd-164,32'd918,32'd1890,32'd2159,32'd-3093,32'd-681,32'd-3618,32'd-6840,32'd4721,32'd-4938,32'd-9584,32'd3254,32'd3732,32'd-2230,32'd-5791,32'd4948,32'd4746,32'd-1161,32'd-3886,32'd-85,32'd-1381,32'd-2434,32'd-1311,32'd-2912,32'd-575,32'd15644,32'd192,32'd892,32'd-2966,32'd-13603,32'd-5747,32'd8261,32'd83,32'd-2712,32'd-1962,32'd-1662,32'd-2204,32'd3520,32'd2512,32'd-8920,32'd-5092,32'd2012,32'd2165,32'd6958,32'd-1777,32'd304,32'd-4755,32'd10830,32'd5322,32'd-3859,32'd4025,32'd-2259,32'd-4643,32'd17109,32'd-7592,32'd6479,32'd2061,32'd5854,32'd-3488,32'd-17919,32'd-601,32'd-23808,32'd6489,32'd-5078,32'd5180,32'd-2980,32'd-14208,32'd-544,32'd3798,32'd2824,32'd-5053,32'd8613,32'd985,32'd-17167,32'd-3725,32'd-6811,32'd4030,32'd1121,32'd-3693,32'd-1348,32'd-1740,32'd192,32'd6352,32'd2183,32'd2995,32'd-2089,32'd-6777,32'd-2070,32'd-4272,32'd-504,32'd-603,32'd-11035,32'd-33,32'd12636,32'd2391,32'd8466,32'd-9062,32'd-10234,32'd12255,32'd6088,32'd-15214,32'd-1876,32'd6914,32'd1168,32'd1441,32'd-3618,32'd9296,32'd-4353,32'd3376,32'd-9921,32'd-6074,32'd4724,32'd4270,32'd-3623,32'd-9594,32'd60,32'd-5175,32'd275,32'd1291,32'd1541,32'd79,32'd-4572,32'd-5000,32'd-1933,32'd-1921,32'd-1713,32'd-2060,32'd-3234,32'd2795,32'd851,32'd8505,32'd13017,32'd-3510,32'd1646,32'd-502,32'd-1868,32'd-2773,32'd2414,32'd-162,32'd-3527,32'd-957,32'd-9028,32'd-75,32'd527,32'd1077,32'd335,32'd-4965,32'd-4514,32'd-3498,32'd10273,32'd-5253,32'd1837,32'd-1175,32'd-7153,32'd1600,32'd1540,32'd6210,32'd-5043,32'd-7822,32'd2878,32'd8798,32'd4028,32'd600,32'd-2524,32'd1257,32'd13496,32'd576,32'd-2800,32'd-8481,32'd-3869,32'd-8168,32'd1765,32'd3107,32'd-10292,32'd2475,32'd1791,32'd-1091,32'd2541,32'd2064,32'd-11650,32'd1367,32'd581,32'd547,32'd2279,32'd1252,32'd5678,32'd2027,32'd1302,32'd-2301,32'd2059,32'd5703,32'd4680,32'd1749,32'd2534,32'd6064,32'd2631,32'd-2023,32'd4824,32'd-989,32'd993,32'd5424,32'd-898,32'd1414,32'd-2166,32'd2371,32'd-720,32'd4912,32'd4172,32'd9619,32'd-99,32'd3720,32'd3078,32'd-1168,32'd-6547,32'd438,32'd10087,32'd4143,32'd6582,32'd3994,32'd4731,32'd6372,32'd-4826,32'd-2761,32'd1350,32'd1162,32'd-5649,32'd1071,32'd-3864,32'd-3640,32'd-872,32'd-3366,32'd-403,32'd-7558,32'd-2329,32'd-7851,32'd-4694,32'd-1249,32'd-2756,32'd-7397,32'd-2183,32'd1704,32'd-8818,32'd3022,32'd-1265,32'd-4711,32'd-786,32'd-6875,32'd5000,32'd-2001,32'd-1934,32'd-1552,32'd-2399,32'd-2731,32'd-5415,32'd-4968,32'd-1485,32'd-538,32'd-3251,32'd-1237,32'd-2524,32'd5688,32'd-2983,32'd-672,32'd1540,32'd-1580,32'd-3383,32'd-2412,32'd-900,32'd748,32'd-125,32'd-4182,32'd6870,32'd-5981,32'd-5908,32'd-899,32'd-2973,32'd248,32'd-4055,32'd3188,32'd4768,32'd-3869,32'd2624,32'd-7836,32'd5019,32'd-5981,32'd5502,32'd-2480,32'd237,32'd-2331,32'd-439,32'd-49,32'd-1246,32'd-5971,32'd-4233,32'd3310,32'd1348,32'd-3535,32'd-5014,32'd-206,32'd-754,32'd6352,32'd-760,32'd-460,32'd1024,32'd-4670,32'd-2282,32'd1124,32'd-838,32'd21445,32'd21250,32'd-1763,32'd5820,32'd-1065,32'd-6684,32'd-186};
    Wx[64]='{32'd894,32'd5019,32'd-1356,32'd-1984,32'd-650,32'd1312,32'd5263,32'd339,32'd-4267,32'd-242,32'd-4074,32'd-4704,32'd-8369,32'd-1722,32'd1329,32'd-5527,32'd-4982,32'd-1105,32'd-552,32'd283,32'd-622,32'd-3083,32'd-5205,32'd59,32'd-3757,32'd4404,32'd845,32'd-1023,32'd-1706,32'd26,32'd-921,32'd5966,32'd-5527,32'd-1209,32'd-6489,32'd2639,32'd1859,32'd1205,32'd-122,32'd665,32'd66,32'd763,32'd6811,32'd3161,32'd-4575,32'd-4230,32'd1400,32'd-2641,32'd-2827,32'd-1992,32'd-712,32'd5791,32'd-2431,32'd2084,32'd-1821,32'd-4548,32'd-1490,32'd2268,32'd1893,32'd-6108,32'd-5112,32'd1372,32'd-3002,32'd-1794,32'd3903,32'd-3210,32'd-152,32'd-1436,32'd-395,32'd-219,32'd-2797,32'd2941,32'd-5913,32'd222,32'd-1688,32'd-3483,32'd-4870,32'd-3093,32'd-1077,32'd584,32'd-1330,32'd7514,32'd4130,32'd4074,32'd-855,32'd-9023,32'd-3344,32'd-3256,32'd-5014,32'd-662,32'd426,32'd5825,32'd-4848,32'd4345,32'd-5615,32'd-693,32'd592,32'd-4394,32'd-3552,32'd-3723,32'd802,32'd6547,32'd2541,32'd-7294,32'd3376,32'd-643,32'd-7265,32'd-2512,32'd7172,32'd-4643,32'd-11318,32'd-474,32'd-9350,32'd215,32'd5410,32'd4072,32'd3920,32'd2204,32'd-1450,32'd-141,32'd527,32'd453,32'd8100,32'd5971,32'd-2086,32'd-206,32'd-213,32'd2331,32'd6791,32'd-14570,32'd5087,32'd21562,32'd-934,32'd1237,32'd364,32'd4892,32'd9067,32'd8916,32'd-6176,32'd21777,32'd-7329,32'd5566,32'd6499,32'd-15654,32'd6899,32'd12333,32'd3369,32'd-1816,32'd-1959,32'd-2180,32'd16044,32'd-13408,32'd-364,32'd-4619,32'd2174,32'd-657,32'd-4187,32'd-3974,32'd8159,32'd-4782,32'd-4521,32'd14091,32'd9301,32'd12578,32'd-18212,32'd2075,32'd-2858,32'd1474,32'd-3127,32'd2252,32'd-656,32'd5537,32'd1483,32'd3366,32'd2281,32'd-4389,32'd-6801,32'd-443,32'd7104,32'd8750,32'd-2067,32'd-14628,32'd3583,32'd-4938,32'd-47,32'd8032,32'd3984,32'd11933,32'd9863,32'd2211,32'd-2775,32'd180,32'd3369,32'd2344,32'd-6733,32'd-2551,32'd4309,32'd-6884,32'd1142,32'd12988,32'd-445,32'd-7680,32'd-983,32'd4199,32'd-2578,32'd1359,32'd-1580,32'd-2374,32'd-553,32'd-2919,32'd4848,32'd4143,32'd-397,32'd4255,32'd819,32'd9990,32'd11621,32'd2949,32'd2321,32'd-231,32'd304,32'd-838,32'd-622,32'd-2104,32'd1695,32'd5751,32'd2543,32'd1578,32'd5966,32'd-9755,32'd2375,32'd5551,32'd7866,32'd-1605,32'd1514,32'd1677,32'd-988,32'd3686,32'd3562,32'd-794,32'd3376,32'd6953,32'd5048,32'd-7358,32'd4338,32'd3801,32'd2028,32'd950,32'd-4934,32'd-3305,32'd6074,32'd-5,32'd2622,32'd2327,32'd1937,32'd-2451,32'd1848,32'd7446,32'd-5649,32'd8569,32'd1334,32'd8984,32'd-549,32'd-3386,32'd-1307,32'd-1844,32'd3056,32'd-207,32'd2049,32'd2524,32'd6225,32'd-2309,32'd-3071,32'd-1693,32'd1773,32'd2971,32'd11826,32'd10566,32'd-3012,32'd919,32'd-4016,32'd3630,32'd4243,32'd-468,32'd-3024,32'd8706,32'd-1315,32'd2171,32'd-1157,32'd-514,32'd-4597,32'd4084,32'd958,32'd1337,32'd-2064,32'd-6655,32'd349,32'd2939,32'd1400,32'd4873,32'd-6357,32'd508,32'd1739,32'd8247,32'd624,32'd6674,32'd6948,32'd-5771,32'd-2624,32'd-3461,32'd288,32'd979,32'd-2270,32'd12695,32'd7563,32'd5043,32'd1408,32'd2670,32'd-3015,32'd-9355,32'd8457,32'd-1549,32'd-2447,32'd-301,32'd-4201,32'd3527,32'd4086,32'd529,32'd2155,32'd-5932,32'd-3308,32'd-3493,32'd910,32'd7314,32'd-5092,32'd5976,32'd-3249,32'd2729,32'd3908,32'd-924,32'd-6992,32'd7485,32'd939,32'd2180,32'd1361,32'd-4108,32'd-1678,32'd-3830,32'd-1914,32'd2038,32'd3256,32'd4975,32'd8017,32'd160,32'd1040,32'd-1340,32'd1193,32'd-723,32'd-4455,32'd-4406,32'd-3320,32'd-737,32'd-4001,32'd939,32'd-1912,32'd-4453,32'd5502,32'd8789,32'd-64,32'd5874,32'd-617,32'd-1771,32'd1673,32'd1638,32'd-5122,32'd3029,32'd12001,32'd219,32'd-338,32'd-2371,32'd-3706,32'd2768,32'd-2106,32'd3383,32'd-2890,32'd9321,32'd-4460,32'd90,32'd-2641,32'd-9418,32'd1154,32'd-962,32'd1516,32'd5219,32'd-725,32'd-4123,32'd4536,32'd-1147,32'd-1868,32'd6123};
    Wx[65]='{32'd171,32'd-2905,32'd-655,32'd4196,32'd1851,32'd3647,32'd308,32'd-1613,32'd1400,32'd-90,32'd2282,32'd847,32'd1962,32'd5888,32'd-301,32'd-2434,32'd6835,32'd2391,32'd-2170,32'd-1197,32'd267,32'd165,32'd523,32'd1500,32'd-3522,32'd-2460,32'd1785,32'd-3715,32'd-1606,32'd-1342,32'd-996,32'd240,32'd-3837,32'd3725,32'd3774,32'd788,32'd1614,32'd-4,32'd3991,32'd-925,32'd745,32'd1834,32'd-2607,32'd121,32'd5595,32'd-584,32'd7026,32'd-1795,32'd121,32'd3,32'd-2512,32'd3251,32'd-142,32'd2861,32'd-2717,32'd-6313,32'd3334,32'd87,32'd-921,32'd-2915,32'd-2839,32'd-2181,32'd3359,32'd1002,32'd4091,32'd-3435,32'd375,32'd-1417,32'd2438,32'd-2692,32'd1964,32'd3112,32'd368,32'd158,32'd-2131,32'd5097,32'd6665,32'd3957,32'd3493,32'd994,32'd1485,32'd9511,32'd1322,32'd7792,32'd-2344,32'd-307,32'd-414,32'd317,32'd738,32'd-2768,32'd-202,32'd-1834,32'd-427,32'd-125,32'd937,32'd-2692,32'd-560,32'd9135,32'd-288,32'd4501,32'd1306,32'd1162,32'd-2370,32'd-1955,32'd-1424,32'd-5317,32'd-7880,32'd-5693,32'd930,32'd-4335,32'd-8950,32'd-10712,32'd4577,32'd5869,32'd9228,32'd-9589,32'd6650,32'd5805,32'd241,32'd1600,32'd2061,32'd-6630,32'd-3188,32'd-7636,32'd-1962,32'd2583,32'd-1116,32'd-1774,32'd-2814,32'd-2406,32'd76,32'd-7177,32'd1203,32'd12919,32'd960,32'd-6049,32'd8422,32'd-3366,32'd-294,32'd-7309,32'd-71,32'd-13652,32'd-7153,32'd-8515,32'd-15087,32'd-6250,32'd6796,32'd-580,32'd-3403,32'd-2131,32'd-811,32'd8789,32'd-842,32'd-12597,32'd2604,32'd-9086,32'd-5942,32'd2060,32'd4995,32'd-2036,32'd-2509,32'd-2861,32'd-11533,32'd666,32'd-6020,32'd5473,32'd-1001,32'd-384,32'd-2929,32'd-304,32'd5708,32'd7280,32'd3200,32'd2646,32'd1038,32'd11386,32'd6567,32'd-6435,32'd2692,32'd-6645,32'd-3188,32'd1004,32'd-145,32'd1065,32'd-1256,32'd5502,32'd3869,32'd-1069,32'd-1770,32'd701,32'd-495,32'd-11005,32'd5371,32'd2442,32'd-14599,32'd-5434,32'd-864,32'd5517,32'd-1166,32'd-7934,32'd594,32'd-5380,32'd-312,32'd948,32'd-2358,32'd803,32'd-7724,32'd-10937,32'd-2368,32'd-1556,32'd4287,32'd-1059,32'd-1939,32'd-3117,32'd1895,32'd5854,32'd-207,32'd3969,32'd5327,32'd-3200,32'd805,32'd-1204,32'd224,32'd1743,32'd385,32'd-3195,32'd1760,32'd1632,32'd-2154,32'd3149,32'd-2066,32'd1713,32'd100,32'd-564,32'd-6284,32'd572,32'd-1552,32'd-3010,32'd671,32'd2403,32'd3649,32'd-8793,32'd-6269,32'd-2260,32'd-7495,32'd479,32'd8037,32'd3017,32'd2912,32'd-333,32'd-3210,32'd2164,32'd-2529,32'd-195,32'd-4382,32'd-3808,32'd5278,32'd-3913,32'd2421,32'd3134,32'd2514,32'd-704,32'd2072,32'd-9770,32'd-13281,32'd-3913,32'd1898,32'd7363,32'd1928,32'd-1602,32'd-5332,32'd1928,32'd3718,32'd-894,32'd-2763,32'd-5258,32'd-2263,32'd-8720,32'd-2216,32'd-623,32'd-2619,32'd368,32'd5371,32'd-3159,32'd2176,32'd-3139,32'd-985,32'd-5776,32'd-6240,32'd-1234,32'd2536,32'd-5375,32'd-4602,32'd2309,32'd4724,32'd2587,32'd160,32'd-2944,32'd-3405,32'd-3503,32'd3520,32'd3039,32'd5234,32'd4675,32'd-4895,32'd2851,32'd2619,32'd3417,32'd-6127,32'd-8618,32'd5458,32'd-651,32'd-5864,32'd2117,32'd-2617,32'd4233,32'd-4853,32'd11171,32'd787,32'd1145,32'd-4226,32'd-1154,32'd3195,32'd-2690,32'd-458,32'd-2707,32'd-5874,32'd-2678,32'd-5947,32'd1970,32'd-15,32'd6909,32'd-14628,32'd394,32'd-4157,32'd-3706,32'd4130,32'd-2993,32'd2044,32'd-195,32'd-640,32'd-6528,32'd4887,32'd-2299,32'd-2052,32'd-1420,32'd2778,32'd4458,32'd6406,32'd3486,32'd-2810,32'd-5527,32'd1287,32'd-337,32'd-2135,32'd-3271,32'd6147,32'd14130,32'd-902,32'd6308,32'd1003,32'd-2266,32'd3352,32'd-4831,32'd555,32'd-2753,32'd-7641,32'd4401,32'd-338,32'd-8251,32'd-2178,32'd3547,32'd950,32'd-1739,32'd-4069,32'd-5463,32'd-12890,32'd-3063,32'd-2004,32'd-6269,32'd1295,32'd200,32'd3039,32'd2512,32'd1572,32'd2437,32'd-1345,32'd-4338,32'd-3142,32'd3317,32'd-1257,32'd-8251,32'd-2700,32'd5327,32'd4235,32'd1427,32'd4589,32'd712,32'd-11181,32'd-4589};
    Wx[66]='{32'd1850,32'd-1746,32'd-1229,32'd-2398,32'd3195,32'd-1928,32'd-4069,32'd-83,32'd2237,32'd4680,32'd1414,32'd-2573,32'd664,32'd-8422,32'd6215,32'd-1937,32'd6220,32'd-3051,32'd887,32'd979,32'd118,32'd5419,32'd4050,32'd2602,32'd751,32'd-3247,32'd1854,32'd-1845,32'd-120,32'd-4995,32'd964,32'd-5839,32'd-944,32'd3754,32'd1647,32'd3251,32'd1499,32'd1571,32'd-5380,32'd-4458,32'd451,32'd2073,32'd2386,32'd3090,32'd1119,32'd-5659,32'd5815,32'd-886,32'd1716,32'd-1325,32'd-1262,32'd651,32'd992,32'd-20,32'd6445,32'd4514,32'd458,32'd-2296,32'd2302,32'd3752,32'd1768,32'd23,32'd2507,32'd3291,32'd1649,32'd2375,32'd-417,32'd-7333,32'd313,32'd-2521,32'd-214,32'd-3457,32'd1247,32'd-5297,32'd2315,32'd642,32'd-4899,32'd-3537,32'd-423,32'd-1525,32'd-1205,32'd1835,32'd2875,32'd1910,32'd2729,32'd-3750,32'd2963,32'd2232,32'd1342,32'd-51,32'd-1849,32'd-852,32'd-2005,32'd-4711,32'd8134,32'd884,32'd-2076,32'd-4741,32'd-1979,32'd-2941,32'd4804,32'd4948,32'd849,32'd7099,32'd11503,32'd-968,32'd830,32'd-4067,32'd-7050,32'd-583,32'd-12421,32'd-858,32'd1013,32'd-10419,32'd-1694,32'd-6293,32'd-11318,32'd4604,32'd-3232,32'd-1856,32'd-512,32'd2469,32'd3000,32'd-1143,32'd-453,32'd-216,32'd-2376,32'd-1066,32'd916,32'd2890,32'd-3737,32'd-24121,32'd-10957,32'd-2175,32'd1430,32'd3249,32'd725,32'd-758,32'd10156,32'd1000,32'd242,32'd5834,32'd5083,32'd4580,32'd1066,32'd9375,32'd-3835,32'd-6396,32'd7011,32'd6318,32'd-9155,32'd-1036,32'd3173,32'd908,32'd3244,32'd9916,32'd5043,32'd3305,32'd-3217,32'd2792,32'd-376,32'd1760,32'd-2834,32'd-6118,32'd-398,32'd-1169,32'd5952,32'd-7612,32'd1783,32'd2866,32'd-786,32'd8305,32'd5371,32'd-4006,32'd844,32'd12148,32'd-5019,32'd1051,32'd925,32'd4775,32'd-5991,32'd-4274,32'd-2385,32'd-16240,32'd-980,32'd-20859,32'd-228,32'd-1448,32'd-5214,32'd-547,32'd-3391,32'd10371,32'd4575,32'd-1776,32'd-12949,32'd1505,32'd2281,32'd-11162,32'd-3769,32'd-1511,32'd1866,32'd-766,32'd-4909,32'd1864,32'd4133,32'd-897,32'd943,32'd-6215,32'd2988,32'd2763,32'd-6298,32'd-2849,32'd1412,32'd1771,32'd5063,32'd-1810,32'd-4104,32'd-7832,32'd-527,32'd-3435,32'd-1307,32'd163,32'd361,32'd-2224,32'd-303,32'd-5639,32'd-2371,32'd-1949,32'd6147,32'd5903,32'd3012,32'd-1446,32'd2558,32'd-4121,32'd6386,32'd773,32'd955,32'd-1262,32'd-7626,32'd3771,32'd383,32'd5371,32'd-5346,32'd2271,32'd2922,32'd-188,32'd-2888,32'd352,32'd883,32'd-4514,32'd1248,32'd-7055,32'd848,32'd3300,32'd-5571,32'd-7709,32'd1179,32'd-3420,32'd-6679,32'd-5644,32'd5849,32'd60,32'd-2326,32'd4062,32'd-626,32'd513,32'd-2221,32'd10722,32'd-3205,32'd-3605,32'd6196,32'd-6035,32'd-950,32'd-5102,32'd115,32'd-4851,32'd-9116,32'd-6953,32'd-5043,32'd5375,32'd-4216,32'd-11582,32'd-1217,32'd-4802,32'd-1542,32'd-11503,32'd-556,32'd1033,32'd5859,32'd-2238,32'd3686,32'd-5605,32'd269,32'd-2055,32'd-4216,32'd686,32'd7841,32'd-544,32'd4499,32'd-3093,32'd2880,32'd-2900,32'd175,32'd-2893,32'd2883,32'd895,32'd-2680,32'd1300,32'd1490,32'd3781,32'd-8671,32'd-541,32'd6108,32'd-190,32'd-148,32'd949,32'd1977,32'd-8745,32'd9912,32'd485,32'd4855,32'd2663,32'd-1203,32'd-1678,32'd4101,32'd-9389,32'd-1403,32'd879,32'd-4072,32'd849,32'd-1014,32'd-506,32'd-1091,32'd-3764,32'd133,32'd4758,32'd6083,32'd8095,32'd-9003,32'd-4655,32'd6474,32'd-912,32'd-1032,32'd-7490,32'd-588,32'd-2739,32'd8647,32'd29,32'd1950,32'd-1719,32'd-4921,32'd856,32'd-9047,32'd-2054,32'd1306,32'd-1022,32'd2739,32'd-668,32'd-993,32'd-1641,32'd1413,32'd-1389,32'd2583,32'd5776,32'd-9946,32'd3220,32'd-8935,32'd585,32'd7324,32'd-7294,32'd241,32'd-10253,32'd2476,32'd-2644,32'd3752,32'd7338,32'd-6132,32'd-698,32'd467,32'd8447,32'd-3217,32'd-2736,32'd2032,32'd-14062,32'd-4335,32'd-13339,32'd48,32'd502,32'd1710,32'd4035,32'd3518,32'd-9023,32'd-476,32'd-10283,32'd-4274,32'd-4011,32'd4672,32'd8032,32'd616,32'd-528};
    Wx[67]='{32'd-890,32'd304,32'd-2296,32'd-1171,32'd243,32'd233,32'd-1962,32'd-3945,32'd-1751,32'd-2924,32'd-2452,32'd107,32'd-1882,32'd-1562,32'd1619,32'd-1007,32'd-438,32'd-4174,32'd-5327,32'd1624,32'd2739,32'd2517,32'd1652,32'd-1056,32'd-1649,32'd2448,32'd-4184,32'd193,32'd68,32'd471,32'd930,32'd-4204,32'd316,32'd0,32'd-5800,32'd-1230,32'd-2277,32'd466,32'd1264,32'd-1379,32'd-236,32'd4035,32'd3457,32'd-3732,32'd2934,32'd130,32'd4055,32'd484,32'd1849,32'd897,32'd-1542,32'd3112,32'd2575,32'd196,32'd2136,32'd4296,32'd3664,32'd-2071,32'd-1232,32'd-1171,32'd-1008,32'd6137,32'd1533,32'd-3327,32'd-3134,32'd558,32'd598,32'd-5043,32'd733,32'd2387,32'd6616,32'd4458,32'd-2136,32'd-1926,32'd-3532,32'd-2519,32'd-5468,32'd1292,32'd3789,32'd-5737,32'd-4465,32'd3461,32'd-446,32'd-3166,32'd1481,32'd-2763,32'd1072,32'd2368,32'd466,32'd3647,32'd-1915,32'd823,32'd-681,32'd486,32'd-2629,32'd-742,32'd-256,32'd3845,32'd-1733,32'd-2180,32'd-2039,32'd2365,32'd-2912,32'd9926,32'd2685,32'd-2248,32'd-192,32'd-10556,32'd2434,32'd4577,32'd2150,32'd956,32'd-953,32'd-107,32'd-3745,32'd2248,32'd-10634,32'd4521,32'd-796,32'd1682,32'd1533,32'd-2570,32'd1260,32'd-175,32'd-509,32'd946,32'd-975,32'd-3476,32'd-3962,32'd3842,32'd2196,32'd1161,32'd-1058,32'd7890,32'd-1479,32'd-12080,32'd-1245,32'd3276,32'd-20566,32'd-6704,32'd-5141,32'd-6416,32'd-9541,32'd-6103,32'd1225,32'd5483,32'd-14423,32'd3598,32'd-5087,32'd-3325,32'd10839,32'd-10419,32'd5576,32'd4284,32'd589,32'd1802,32'd3098,32'd-3093,32'd4621,32'd-844,32'd-4279,32'd5668,32'd8940,32'd-3830,32'd12890,32'd101,32'd984,32'd-14277,32'd-887,32'd-11,32'd-11777,32'd5395,32'd4755,32'd-5405,32'd-103,32'd5244,32'd-4660,32'd-2194,32'd317,32'd1346,32'd-2415,32'd-6533,32'd-4250,32'd7905,32'd3059,32'd-3725,32'd-1962,32'd2403,32'd-4660,32'd1582,32'd3193,32'd-19707,32'd9423,32'd-888,32'd-13583,32'd8627,32'd-8442,32'd-3684,32'd-4257,32'd652,32'd1115,32'd-7666,32'd-619,32'd-2590,32'd2661,32'd457,32'd-1644,32'd-632,32'd-5761,32'd-1505,32'd-3605,32'd-708,32'd285,32'd4460,32'd-2305,32'd-132,32'd3876,32'd3325,32'd3090,32'd-2653,32'd2519,32'd-3103,32'd332,32'd1751,32'd-2379,32'd-2978,32'd4978,32'd-435,32'd-3664,32'd-9594,32'd1441,32'd358,32'd567,32'd-4311,32'd4118,32'd-4418,32'd5883,32'd1309,32'd-7973,32'd-1812,32'd2070,32'd-1000,32'd-3105,32'd283,32'd7954,32'd700,32'd-1545,32'd-321,32'd68,32'd-3881,32'd-3032,32'd-12753,32'd4091,32'd-3454,32'd311,32'd-7553,32'd-7519,32'd1961,32'd-1103,32'd1582,32'd-1428,32'd-7788,32'd-5029,32'd-498,32'd524,32'd-3881,32'd-258,32'd6093,32'd4682,32'd-1094,32'd-1401,32'd1477,32'd1987,32'd-2032,32'd-593,32'd8784,32'd-4077,32'd309,32'd-6362,32'd1385,32'd-1074,32'd-6118,32'd2956,32'd3002,32'd594,32'd-3889,32'd2170,32'd959,32'd-1544,32'd-1472,32'd2963,32'd5380,32'd-1473,32'd2048,32'd-7373,32'd-5620,32'd1218,32'd614,32'd2191,32'd-4743,32'd5693,32'd-1785,32'd7968,32'd-1301,32'd4245,32'd6665,32'd-1478,32'd-1602,32'd-8823,32'd-2949,32'd-8886,32'd-518,32'd2519,32'd7543,32'd-934,32'd-812,32'd-2121,32'd1658,32'd-5625,32'd-2946,32'd4973,32'd-1665,32'd-3381,32'd352,32'd-2297,32'd-434,32'd-4606,32'd-558,32'd-6889,32'd-1925,32'd51,32'd-4118,32'd-840,32'd-5942,32'd-13798,32'd-4187,32'd-5512,32'd891,32'd-6718,32'd-13242,32'd1805,32'd-1693,32'd-1106,32'd1181,32'd4536,32'd-2486,32'd-9492,32'd2076,32'd9814,32'd-2663,32'd924,32'd-3186,32'd10390,32'd-1542,32'd8164,32'd5395,32'd-6357,32'd4938,32'd1170,32'd-1359,32'd-2880,32'd-3937,32'd-5771,32'd-1374,32'd-2529,32'd7568,32'd-2500,32'd7910,32'd-1428,32'd-5546,32'd37,32'd-2531,32'd-7602,32'd-5444,32'd-4504,32'd-2758,32'd-5639,32'd3974,32'd-5654,32'd-1021,32'd-949,32'd1728,32'd5449,32'd-2719,32'd1645,32'd1833,32'd3325,32'd-399,32'd-2364,32'd7153,32'd-1842,32'd6884,32'd-7622,32'd-6967,32'd3801,32'd-1981,32'd-339,32'd-1480,32'd-147,32'd-6254};
    Wx[68]='{32'd1229,32'd-4042,32'd-192,32'd-2424,32'd938,32'd-953,32'd5932,32'd4494,32'd1971,32'd2152,32'd2734,32'd-1038,32'd5410,32'd-541,32'd4338,32'd5981,32'd5458,32'd440,32'd308,32'd-2775,32'd-348,32'd-366,32'd1042,32'd80,32'd1077,32'd2086,32'd3100,32'd589,32'd4086,32'd-562,32'd1580,32'd5541,32'd6591,32'd5766,32'd1374,32'd-4477,32'd5473,32'd-3122,32'd734,32'd1667,32'd3120,32'd14,32'd2707,32'd1257,32'd-2844,32'd4052,32'd5922,32'd5107,32'd4675,32'd2795,32'd2773,32'd1492,32'd2290,32'd363,32'd-125,32'd5585,32'd1351,32'd1479,32'd3017,32'd4951,32'd363,32'd787,32'd-1564,32'd750,32'd14462,32'd297,32'd1716,32'd4660,32'd-196,32'd-2043,32'd-1494,32'd6904,32'd3806,32'd-5864,32'd1242,32'd487,32'd1018,32'd3090,32'd-185,32'd1668,32'd326,32'd1907,32'd1071,32'd6401,32'd1145,32'd3879,32'd-811,32'd315,32'd-920,32'd2998,32'd3525,32'd-530,32'd-3781,32'd2973,32'd5590,32'd-455,32'd1740,32'd4838,32'd3293,32'd6499,32'd344,32'd6577,32'd2780,32'd-5317,32'd-9218,32'd344,32'd-1826,32'd3825,32'd-1381,32'd3054,32'd-5053,32'd-2756,32'd2797,32'd-16162,32'd-883,32'd-1257,32'd-13330,32'd5126,32'd-122,32'd236,32'd-855,32'd-3293,32'd-1428,32'd-3208,32'd443,32'd-2739,32'd-4377,32'd-302,32'd-1734,32'd3010,32'd125,32'd-1326,32'd6684,32'd-3662,32'd1734,32'd-3403,32'd-3408,32'd123,32'd17324,32'd12363,32'd-1063,32'd-15546,32'd4282,32'd2551,32'd4877,32'd-3769,32'd482,32'd-249,32'd10703,32'd-5532,32'd-16025,32'd33,32'd-2054,32'd-9741,32'd-998,32'd3640,32'd3977,32'd357,32'd692,32'd4040,32'd-5371,32'd711,32'd2454,32'd-4008,32'd-4394,32'd-701,32'd4353,32'd-3127,32'd2724,32'd-2270,32'd5512,32'd1944,32'd-681,32'd-7211,32'd-659,32'd-10458,32'd8657,32'd-3566,32'd1052,32'd4755,32'd-4411,32'd-2934,32'd13574,32'd-698,32'd-1346,32'd-7124,32'd-1300,32'd-5878,32'd-792,32'd-3979,32'd-7353,32'd-2729,32'd13662,32'd157,32'd-2441,32'd4392,32'd227,32'd18300,32'd-5004,32'd12578,32'd969,32'd-5273,32'd936,32'd-582,32'd-2427,32'd-416,32'd-3540,32'd-3659,32'd-1232,32'd-698,32'd-2946,32'd1739,32'd-5678,32'd583,32'd-1160,32'd-6875,32'd-1079,32'd-2386,32'd-1301,32'd469,32'd-1882,32'd-274,32'd-5751,32'd7397,32'd1601,32'd-709,32'd5209,32'd2749,32'd3518,32'd-7416,32'd5756,32'd-63,32'd4020,32'd-5493,32'd-3693,32'd-1352,32'd-3906,32'd-2271,32'd-1124,32'd-7602,32'd1212,32'd162,32'd158,32'd848,32'd-9599,32'd-7416,32'd-10048,32'd-131,32'd3798,32'd-930,32'd-354,32'd-8691,32'd1739,32'd-4291,32'd-1713,32'd-8325,32'd-624,32'd128,32'd-1536,32'd-7329,32'd3234,32'd5786,32'd-3869,32'd70,32'd2514,32'd-1199,32'd841,32'd-1273,32'd-888,32'd-3627,32'd-6645,32'd-6503,32'd2399,32'd969,32'd1516,32'd-1937,32'd-5747,32'd2624,32'd-2507,32'd-1666,32'd-1367,32'd-4331,32'd-413,32'd-7421,32'd404,32'd-691,32'd708,32'd1386,32'd6743,32'd2238,32'd2426,32'd1406,32'd6103,32'd4201,32'd7275,32'd-889,32'd-1171,32'd-3159,32'd-4807,32'd883,32'd3847,32'd-859,32'd2529,32'd2435,32'd-1170,32'd-1635,32'd-3234,32'd-4104,32'd6879,32'd-2250,32'd6694,32'd2043,32'd666,32'd-2788,32'd-3098,32'd1407,32'd529,32'd2509,32'd1707,32'd1531,32'd-9697,32'd3420,32'd-1787,32'd3054,32'd7094,32'd588,32'd4753,32'd-3188,32'd6499,32'd-7519,32'd-584,32'd2470,32'd5195,32'd628,32'd-7900,32'd-1824,32'd-978,32'd-5585,32'd1111,32'd3251,32'd-586,32'd1353,32'd6044,32'd-3674,32'd77,32'd-3522,32'd-11611,32'd3244,32'd-621,32'd-1163,32'd-1030,32'd-4584,32'd5830,32'd-456,32'd-4753,32'd4060,32'd6713,32'd-571,32'd4804,32'd-7055,32'd-1441,32'd2600,32'd-4553,32'd1353,32'd3413,32'd4970,32'd3483,32'd1330,32'd12666,32'd-4060,32'd-1495,32'd-8896,32'd3522,32'd3259,32'd2749,32'd-2369,32'd6440,32'd4274,32'd-7973,32'd-373,32'd-2209,32'd201,32'd4184,32'd-9399,32'd2607,32'd-1271,32'd2836,32'd-2971,32'd1097,32'd-4853,32'd6840,32'd-671,32'd4367,32'd-3791,32'd1270,32'd-1185,32'd3120,32'd1445,32'd3933,32'd-3515};
    Wx[69]='{32'd-1447,32'd-2595,32'd1517,32'd-339,32'd-855,32'd-330,32'd427,32'd-1160,32'd-2905,32'd-2519,32'd-7836,32'd-125,32'd-437,32'd6538,32'd-2399,32'd57,32'd-3576,32'd-6059,32'd-3203,32'd-3046,32'd-1901,32'd1741,32'd-3049,32'd-964,32'd1519,32'd-2734,32'd206,32'd-2629,32'd-3151,32'd-916,32'd-1187,32'd-7768,32'd-294,32'd-3618,32'd-4645,32'd-192,32'd1062,32'd-2922,32'd2224,32'd-1887,32'd-378,32'd-1593,32'd-550,32'd10878,32'd-4982,32'd-2336,32'd9335,32'd1341,32'd-4738,32'd-2656,32'd2252,32'd-10205,32'd-4692,32'd639,32'd-3422,32'd-6953,32'd1710,32'd-2241,32'd-2836,32'd-1007,32'd-3476,32'd-3852,32'd1840,32'd-5581,32'd1207,32'd-4587,32'd1271,32'd2319,32'd-1293,32'd891,32'd-659,32'd619,32'd134,32'd-2456,32'd-414,32'd-3178,32'd2626,32'd3815,32'd-1358,32'd141,32'd1527,32'd4638,32'd38,32'd-1119,32'd-4819,32'd-5893,32'd-505,32'd970,32'd-183,32'd-375,32'd1089,32'd-1391,32'd2731,32'd651,32'd-4558,32'd-3356,32'd344,32'd-7651,32'd-3920,32'd-1793,32'd-1319,32'd-741,32'd-5712,32'd-1271,32'd-2573,32'd1728,32'd748,32'd-2374,32'd-3447,32'd-1850,32'd-1185,32'd-2225,32'd1473,32'd794,32'd-2766,32'd-572,32'd5214,32'd9750,32'd-3200,32'd1577,32'd-2644,32'd1801,32'd3239,32'd-6303,32'd-4960,32'd6596,32'd943,32'd-419,32'd-6445,32'd-536,32'd1507,32'd4780,32'd11191,32'd6845,32'd350,32'd2814,32'd284,32'd6796,32'd3093,32'd-19433,32'd-4392,32'd595,32'd5834,32'd381,32'd5698,32'd-13212,32'd13671,32'd-557,32'd-7998,32'd2885,32'd3093,32'd-3146,32'd-1611,32'd-9443,32'd-3549,32'd17939,32'd-6899,32'd1350,32'd-8095,32'd4233,32'd4414,32'd9345,32'd1162,32'd6875,32'd7329,32'd4096,32'd3928,32'd5917,32'd-9,32'd250,32'd5263,32'd14726,32'd2609,32'd3483,32'd341,32'd-2120,32'd5986,32'd-3996,32'd-141,32'd-1229,32'd-38,32'd-4541,32'd6147,32'd16660,32'd4604,32'd-4599,32'd2365,32'd8691,32'd-2052,32'd289,32'd-7246,32'd11757,32'd12666,32'd-45,32'd-12382,32'd-2408,32'd-1839,32'd-871,32'd3269,32'd8701,32'd1857,32'd2406,32'd3615,32'd-3095,32'd46,32'd-136,32'd-234,32'd3527,32'd1268,32'd-5849,32'd-869,32'd-1413,32'd4621,32'd-3708,32'd-1771,32'd4450,32'd814,32'd-7690,32'd2729,32'd128,32'd-1519,32'd68,32'd549,32'd5610,32'd712,32'd-888,32'd4672,32'd-1364,32'd4003,32'd-5024,32'd-764,32'd-2770,32'd-6689,32'd-8676,32'd3999,32'd-5649,32'd-2108,32'd4260,32'd-406,32'd-438,32'd-572,32'd-3916,32'd2370,32'd-5576,32'd4328,32'd6459,32'd10361,32'd-2492,32'd325,32'd-1772,32'd919,32'd6811,32'd5888,32'd-11601,32'd-1068,32'd-4072,32'd-6845,32'd2500,32'd-2447,32'd-2059,32'd1943,32'd2666,32'd-1612,32'd5048,32'd-6748,32'd3200,32'd-1503,32'd-4191,32'd-4035,32'd-95,32'd-3559,32'd-8178,32'd-2800,32'd-2480,32'd1019,32'd6372,32'd4211,32'd-956,32'd-4750,32'd9072,32'd1040,32'd2780,32'd4257,32'd152,32'd-407,32'd-2105,32'd1802,32'd418,32'd-907,32'd-2937,32'd1561,32'd1604,32'd-1444,32'd-1525,32'd-6752,32'd75,32'd2663,32'd5678,32'd1202,32'd-4880,32'd6152,32'd4179,32'd9638,32'd171,32'd25,32'd9013,32'd2198,32'd7309,32'd-5864,32'd-11630,32'd-4978,32'd-232,32'd-1545,32'd499,32'd-6860,32'd3911,32'd-5312,32'd2978,32'd-642,32'd-4587,32'd8701,32'd2386,32'd5117,32'd2496,32'd1567,32'd1378,32'd4213,32'd-3027,32'd-691,32'd-1159,32'd-2585,32'd-6967,32'd2514,32'd-5273,32'd-1435,32'd-1499,32'd5317,32'd3254,32'd-5151,32'd-8120,32'd-1468,32'd-7861,32'd4829,32'd-3393,32'd-1986,32'd4755,32'd-2171,32'd-1821,32'd1257,32'd1937,32'd-2050,32'd1821,32'd9296,32'd-4187,32'd11640,32'd119,32'd-6201,32'd3759,32'd-185,32'd-3232,32'd-6806,32'd-5751,32'd-3762,32'd-5078,32'd2440,32'd10703,32'd3098,32'd5346,32'd3291,32'd-3000,32'd3229,32'd-11044,32'd-6513,32'd664,32'd-3381,32'd2697,32'd4655,32'd-4016,32'd2081,32'd3051,32'd2127,32'd7177,32'd1495,32'd4145,32'd-3735,32'd-1983,32'd-5253,32'd-541,32'd-4360,32'd1052,32'd7270,32'd-51,32'd-1233,32'd-3337,32'd-1578,32'd1413,32'd1365,32'd-2553,32'd-2067,32'd-5014};
    Wx[70]='{32'd-1296,32'd8701,32'd1584,32'd-1429,32'd974,32'd786,32'd1901,32'd5195,32'd1984,32'd632,32'd1364,32'd1093,32'd1166,32'd-300,32'd4636,32'd6860,32'd9340,32'd5214,32'd1804,32'd-479,32'd-809,32'd1562,32'd40,32'd-3483,32'd-1157,32'd-372,32'd2375,32'd1258,32'd-20,32'd-1947,32'd673,32'd-3593,32'd-3874,32'd2469,32'd-1033,32'd-126,32'd-1848,32'd-721,32'd-5927,32'd-6186,32'd3344,32'd-795,32'd-2449,32'd-2043,32'd-2260,32'd-1674,32'd-620,32'd4948,32'd-3427,32'd826,32'd3073,32'd247,32'd-345,32'd-1857,32'd2929,32'd6948,32'd-587,32'd1230,32'd-581,32'd353,32'd-329,32'd472,32'd-1448,32'd2014,32'd2890,32'd842,32'd-241,32'd1917,32'd-2048,32'd1645,32'd972,32'd-4631,32'd1866,32'd-4487,32'd1424,32'd3212,32'd-5410,32'd275,32'd-2500,32'd1333,32'd1512,32'd-1853,32'd-563,32'd3190,32'd-5454,32'd3413,32'd-1555,32'd-2008,32'd6801,32'd-3862,32'd422,32'd-3840,32'd1881,32'd29,32'd-6386,32'd-1676,32'd4067,32'd-1734,32'd3439,32'd545,32'd2343,32'd11103,32'd1137,32'd481,32'd-2191,32'd1491,32'd-4501,32'd-4951,32'd-59,32'd141,32'd10351,32'd-3796,32'd3803,32'd11318,32'd-13808,32'd-222,32'd3713,32'd3757,32'd-4360,32'd430,32'd-1733,32'd607,32'd-228,32'd10869,32'd-172,32'd4980,32'd4638,32'd-9511,32'd-13906,32'd-3059,32'd5571,32'd-976,32'd1560,32'd14472,32'd-2396,32'd3525,32'd-1138,32'd-1002,32'd2839,32'd-7587,32'd1054,32'd24433,32'd-8833,32'd8696,32'd1348,32'd-3901,32'd27,32'd-3134,32'd-2476,32'd9018,32'd-6611,32'd2471,32'd7006,32'd1407,32'd-2895,32'd-770,32'd1109,32'd-1202,32'd-5800,32'd799,32'd-2705,32'd548,32'd4780,32'd-3515,32'd2753,32'd2048,32'd-3918,32'd1329,32'd3864,32'd-3559,32'd3498,32'd-17207,32'd-7407,32'd3093,32'd-829,32'd-6293,32'd3618,32'd-6601,32'd-3337,32'd-1459,32'd1417,32'd12939,32'd-8085,32'd2819,32'd-2990,32'd-8056,32'd903,32'd-3691,32'd-7802,32'd-75,32'd-2104,32'd-1706,32'd-3640,32'd461,32'd4880,32'd-2331,32'd-3781,32'd-9873,32'd-145,32'd2717,32'd-445,32'd-4316,32'd3596,32'd-3037,32'd825,32'd1748,32'd-4301,32'd3710,32'd-3076,32'd3452,32'd-1015,32'd1722,32'd-7348,32'd-744,32'd4655,32'd3266,32'd1607,32'd874,32'd-1492,32'd-1446,32'd168,32'd3767,32'd-46,32'd-1268,32'd-7841,32'd-4240,32'd-8315,32'd2486,32'd-2032,32'd-2220,32'd-674,32'd3510,32'd9414,32'd-95,32'd-4602,32'd-6049,32'd-3051,32'd-1346,32'd5981,32'd2851,32'd-5537,32'd-588,32'd2546,32'd6416,32'd-4309,32'd-850,32'd-781,32'd8984,32'd396,32'd4873,32'd-1346,32'd-5083,32'd-263,32'd-1232,32'd813,32'd-63,32'd-6235,32'd2546,32'd-3786,32'd2817,32'd7373,32'd-3562,32'd-7597,32'd2081,32'd3474,32'd-1606,32'd97,32'd-4013,32'd-950,32'd1605,32'd-1914,32'd370,32'd-545,32'd1254,32'd1154,32'd1275,32'd-919,32'd-2717,32'd-2673,32'd-3791,32'd2165,32'd-6191,32'd-3845,32'd-6264,32'd-3105,32'd6425,32'd2871,32'd1203,32'd-11093,32'd-2242,32'd-5581,32'd2592,32'd3210,32'd1462,32'd315,32'd4106,32'd-6918,32'd6718,32'd273,32'd-4931,32'd2778,32'd634,32'd-198,32'd2995,32'd-2333,32'd4013,32'd3315,32'd4172,32'd2524,32'd8740,32'd-3322,32'd2673,32'd-1661,32'd-6625,32'd-1392,32'd3969,32'd3344,32'd4172,32'd-2276,32'd-3815,32'd-4655,32'd3322,32'd-230,32'd-2548,32'd-7358,32'd-1439,32'd-2131,32'd5122,32'd-1549,32'd622,32'd477,32'd-5126,32'd-532,32'd-4147,32'd-13398,32'd-5000,32'd-1881,32'd-297,32'd4467,32'd366,32'd-1206,32'd-3876,32'd4077,32'd4626,32'd3112,32'd-4555,32'd-2578,32'd925,32'd3591,32'd738,32'd10087,32'd2570,32'd208,32'd-3010,32'd-880,32'd4980,32'd-1136,32'd-85,32'd-8417,32'd-2561,32'd1141,32'd-3364,32'd-4851,32'd8671,32'd8935,32'd-9809,32'd-808,32'd-6845,32'd-10332,32'd-1702,32'd-4904,32'd-3937,32'd2502,32'd3957,32'd6254,32'd-5424,32'd-3522,32'd-1737,32'd-3249,32'd-2675,32'd5986,32'd-1398,32'd-2768,32'd-4624,32'd-10976,32'd6264,32'd5092,32'd4365,32'd476,32'd-7192,32'd-2805,32'd-2797,32'd5703,32'd-309,32'd-4094,32'd11406,32'd-3239,32'd-874,32'd-683,32'd-3093};
    Wx[71]='{32'd-2653,32'd35,32'd1745,32'd1099,32'd-666,32'd-1396,32'd1441,32'd4685,32'd-260,32'd-4392,32'd3310,32'd3212,32'd4643,32'd-314,32'd-4768,32'd5107,32'd546,32'd-1110,32'd1529,32'd-518,32'd1224,32'd1694,32'd23,32'd-358,32'd4699,32'd-2504,32'd1036,32'd-1386,32'd4895,32'd-5532,32'd-1875,32'd4492,32'd911,32'd4887,32'd-2590,32'd-4716,32'd2291,32'd-845,32'd-4477,32'd3437,32'd551,32'd-4313,32'd-3557,32'd-2144,32'd-5419,32'd-3225,32'd11953,32'd-1956,32'd4680,32'd2687,32'd4189,32'd-2307,32'd543,32'd3173,32'd-226,32'd3691,32'd2895,32'd-1989,32'd-1894,32'd3850,32'd415,32'd304,32'd510,32'd-4313,32'd5048,32'd1545,32'd-1723,32'd7304,32'd1749,32'd874,32'd4121,32'd-1737,32'd3422,32'd-5444,32'd2714,32'd3710,32'd4223,32'd-5029,32'd-201,32'd2043,32'd3305,32'd5625,32'd-3933,32'd-2736,32'd1542,32'd6508,32'd866,32'd3161,32'd1562,32'd3200,32'd977,32'd-8642,32'd-71,32'd1165,32'd186,32'd1458,32'd3000,32'd-4265,32'd4440,32'd3076,32'd213,32'd-6250,32'd-683,32'd-8740,32'd-6508,32'd-2396,32'd-2507,32'd-3288,32'd-4855,32'd-5141,32'd-12431,32'd8730,32'd10283,32'd7675,32'd8046,32'd992,32'd9624,32'd2322,32'd2949,32'd30,32'd205,32'd9165,32'd-5107,32'd4765,32'd1795,32'd2276,32'd-7529,32'd-575,32'd21250,32'd2636,32'd-5537,32'd-353,32'd-4045,32'd-466,32'd5117,32'd1584,32'd-571,32'd3337,32'd3164,32'd10527,32'd-3127,32'd9794,32'd-3298,32'd3388,32'd12392,32'd-9482,32'd-3857,32'd-14248,32'd5366,32'd-11015,32'd-15703,32'd-13242,32'd-9511,32'd-5693,32'd-4309,32'd8891,32'd-2626,32'd1441,32'd1140,32'd4040,32'd1549,32'd6508,32'd10849,32'd2495,32'd14697,32'd-7729,32'd7944,32'd531,32'd-2890,32'd2120,32'd9604,32'd4445,32'd-1196,32'd2680,32'd-2232,32'd-6381,32'd5595,32'd-1801,32'd-4462,32'd-3825,32'd-6557,32'd-1365,32'd4458,32'd-11132,32'd7495,32'd922,32'd2094,32'd8457,32'd-5800,32'd5073,32'd3054,32'd33281,32'd-7055,32'd1205,32'd-2111,32'd-1649,32'd2258,32'd6933,32'd913,32'd6289,32'd974,32'd-821,32'd2205,32'd4206,32'd-905,32'd-1773,32'd4392,32'd2939,32'd436,32'd-3750,32'd2071,32'd351,32'd-784,32'd1317,32'd-992,32'd-5908,32'd-9042,32'd-4729,32'd3112,32'd-2467,32'd-1059,32'd1928,32'd2995,32'd2961,32'd3146,32'd-3547,32'd4636,32'd-74,32'd-7583,32'd8808,32'd3159,32'd-13085,32'd-4753,32'd-4775,32'd-5463,32'd2238,32'd-1633,32'd-874,32'd-3032,32'd-6313,32'd4062,32'd-9667,32'd3266,32'd-5029,32'd-621,32'd1773,32'd-2951,32'd357,32'd5815,32'd-4365,32'd-6953,32'd-11455,32'd-1689,32'd-481,32'd5688,32'd7954,32'd-742,32'd-1058,32'd2293,32'd-3991,32'd4692,32'd3273,32'd5146,32'd1608,32'd16425,32'd-1536,32'd-4353,32'd2778,32'd-889,32'd-2773,32'd-2396,32'd-9331,32'd-3691,32'd-1663,32'd854,32'd-1456,32'd-11396,32'd-2646,32'd-2573,32'd-4050,32'd5512,32'd-3842,32'd-1267,32'd-13398,32'd4494,32'd1158,32'd2332,32'd-1904,32'd2668,32'd-3032,32'd3950,32'd-4580,32'd-3339,32'd5449,32'd5893,32'd-7534,32'd2375,32'd-3859,32'd3427,32'd-6811,32'd-6972,32'd4194,32'd5742,32'd-9619,32'd217,32'd-3151,32'd2739,32'd1124,32'd-315,32'd-8969,32'd6538,32'd7299,32'd733,32'd-8046,32'd-2980,32'd-4431,32'd-3251,32'd-9370,32'd822,32'd-2875,32'd-3994,32'd-1889,32'd4724,32'd2812,32'd-291,32'd-4995,32'd7397,32'd-4526,32'd4902,32'd3630,32'd-1057,32'd-5039,32'd1340,32'd1030,32'd-1942,32'd1188,32'd-2305,32'd603,32'd-7617,32'd3212,32'd1153,32'd-6542,32'd4057,32'd-5234,32'd14,32'd4001,32'd1223,32'd-7036,32'd346,32'd-4533,32'd-4504,32'd-10908,32'd1944,32'd-1203,32'd9301,32'd7138,32'd-634,32'd2302,32'd-960,32'd-542,32'd1984,32'd3706,32'd8876,32'd2570,32'd5390,32'd-6269,32'd-3986,32'd1216,32'd1475,32'd-5639,32'd-986,32'd-418,32'd-1322,32'd603,32'd7729,32'd11074,32'd-2147,32'd-3771,32'd2817,32'd-8149,32'd3420,32'd-58,32'd-10585,32'd797,32'd7338,32'd-4709,32'd7504,32'd-876,32'd1557,32'd-10078,32'd5649,32'd-3537,32'd5463,32'd10947,32'd-5854,32'd-8139,32'd-268,32'd-1171,32'd2824,32'd-10585};
    Wx[72]='{32'd24,32'd-6411,32'd-2768,32'd-3674,32'd-1595,32'd1599,32'd-6235,32'd-4274,32'd-2519,32'd2233,32'd1074,32'd-3791,32'd-1362,32'd-1372,32'd1982,32'd-6982,32'd-4389,32'd-1723,32'd-3200,32'd446,32'd-1306,32'd1788,32'd-1882,32'd-3366,32'd-2824,32'd835,32'd-1639,32'd-2011,32'd-4084,32'd5117,32'd-4023,32'd-5122,32'd-3730,32'd-4389,32'd1425,32'd3586,32'd178,32'd-3625,32'd-2242,32'd-535,32'd-3718,32'd-6259,32'd-2810,32'd941,32'd-1394,32'd-4794,32'd-1845,32'd1450,32'd-2169,32'd-932,32'd-1356,32'd-7246,32'd-1425,32'd-878,32'd1263,32'd-12031,32'd2119,32'd-2641,32'd3449,32'd-3925,32'd-3256,32'd-2651,32'd-2320,32'd-745,32'd-1723,32'd14,32'd1021,32'd-5517,32'd-2768,32'd779,32'd-3339,32'd2099,32'd-902,32'd-766,32'd-2127,32'd-1950,32'd-4306,32'd1412,32'd-15,32'd695,32'd1992,32'd857,32'd1063,32'd1458,32'd2077,32'd2281,32'd584,32'd1895,32'd-2763,32'd-3796,32'd2121,32'd75,32'd-2264,32'd-1766,32'd-3757,32'd-5761,32'd-2595,32'd-9003,32'd-4531,32'd1121,32'd-949,32'd18046,32'd-1894,32'd-1350,32'd4411,32'd-167,32'd-7221,32'd665,32'd5024,32'd-3754,32'd-4943,32'd-4006,32'd178,32'd-1064,32'd-25449,32'd4709,32'd-742,32'd4211,32'd-1024,32'd-2037,32'd-2443,32'd-8022,32'd-3427,32'd-5825,32'd1391,32'd2423,32'd174,32'd7099,32'd8002,32'd-2687,32'd-1524,32'd-7939,32'd-461,32'd-14345,32'd-2106,32'd2238,32'd-5468,32'd-11748,32'd-3364,32'd-6254,32'd11201,32'd12529,32'd6137,32'd-2340,32'd-5097,32'd-4916,32'd-922,32'd7753,32'd-682,32'd1591,32'd-4587,32'd-13642,32'd-2415,32'd-11259,32'd-1373,32'd-7119,32'd6376,32'd5688,32'd332,32'd-6069,32'd2768,32'd11054,32'd-6533,32'd-6440,32'd-16621,32'd3210,32'd691,32'd-11435,32'd1107,32'd-433,32'd278,32'd3918,32'd-3076,32'd-9746,32'd3759,32'd1713,32'd-15380,32'd4760,32'd2276,32'd-1938,32'd6914,32'd17451,32'd-338,32'd-2722,32'd3342,32'd-15029,32'd-2113,32'd-10,32'd973,32'd-3315,32'd-8500,32'd-7436,32'd11611,32'd114,32'd5649,32'd-5756,32'd4306,32'd-4497,32'd164,32'd-6420,32'd1340,32'd4287,32'd-407,32'd-3173,32'd2028,32'd101,32'd2203,32'd-2644,32'd10273,32'd-653,32'd6381,32'd918,32'd2856,32'd-7729,32'd3266,32'd1364,32'd2293,32'd-5668,32'd600,32'd229,32'd-673,32'd-1342,32'd4235,32'd906,32'd-1914,32'd1058,32'd-4291,32'd-2961,32'd4860,32'd-6210,32'd-270,32'd-2773,32'd5678,32'd5263,32'd-6826,32'd-3049,32'd344,32'd3693,32'd5156,32'd3496,32'd120,32'd2365,32'd-631,32'd81,32'd-2861,32'd-1838,32'd-165,32'd-252,32'd-1750,32'd2863,32'd401,32'd-4135,32'd167,32'd-6870,32'd-3139,32'd13447,32'd-1062,32'd-1876,32'd-9624,32'd3239,32'd-3476,32'd-4201,32'd10917,32'd-447,32'd-6064,32'd1412,32'd2199,32'd-16201,32'd1557,32'd-1520,32'd-5219,32'd2609,32'd-3840,32'd-4313,32'd-167,32'd471,32'd-151,32'd-443,32'd3391,32'd-583,32'd50,32'd-3117,32'd-197,32'd6538,32'd4350,32'd2290,32'd-1170,32'd1212,32'd477,32'd-281,32'd-2492,32'd692,32'd-7578,32'd758,32'd-7001,32'd3369,32'd-187,32'd761,32'd-2683,32'd5190,32'd10849,32'd-4819,32'd-66,32'd-2709,32'd6845,32'd9077,32'd-4694,32'd3769,32'd6899,32'd2790,32'd-4084,32'd-4714,32'd1654,32'd-4365,32'd-1751,32'd3747,32'd5805,32'd-10205,32'd5014,32'd-4689,32'd6738,32'd-2420,32'd2536,32'd-232,32'd-4672,32'd-4218,32'd-2976,32'd5581,32'd-4719,32'd-5781,32'd2200,32'd-2376,32'd2963,32'd-650,32'd4956,32'd49,32'd3996,32'd1654,32'd-1136,32'd2692,32'd-3466,32'd-6044,32'd-4838,32'd-7641,32'd-1749,32'd-646,32'd6865,32'd3852,32'd-1146,32'd-427,32'd36,32'd2778,32'd-6000,32'd-3728,32'd1805,32'd6040,32'd-2739,32'd-4663,32'd-4729,32'd2036,32'd-4758,32'd-3977,32'd-1092,32'd4848,32'd629,32'd5722,32'd1084,32'd-5175,32'd607,32'd7128,32'd2174,32'd-4699,32'd-1723,32'd-5971,32'd1929,32'd-3281,32'd-308,32'd-6079,32'd-946,32'd5332,32'd-1605,32'd1845,32'd27,32'd1485,32'd10185,32'd5371,32'd4606,32'd-508,32'd-324,32'd-1350,32'd-755,32'd-7016,32'd-6269,32'd249,32'd-10498,32'd483,32'd886,32'd397,32'd-4536,32'd1008};
    Wx[73]='{32'd1799,32'd-900,32'd-4531,32'd2817,32'd2966,32'd1423,32'd1738,32'd-2990,32'd1622,32'd744,32'd9580,32'd-4528,32'd4265,32'd406,32'd8417,32'd871,32'd6518,32'd639,32'd2644,32'd1767,32'd-973,32'd-1791,32'd-3374,32'd157,32'd-2687,32'd-1954,32'd-3754,32'd1937,32'd-879,32'd1491,32'd2114,32'd10576,32'd-877,32'd-1779,32'd2362,32'd5957,32'd4812,32'd1700,32'd4365,32'd6250,32'd5781,32'd8911,32'd4160,32'd-1829,32'd1762,32'd3701,32'd-645,32'd4428,32'd2415,32'd-48,32'd-1721,32'd917,32'd-1141,32'd4079,32'd-1994,32'd-107,32'd-1943,32'd5239,32'd-479,32'd3356,32'd40,32'd-583,32'd435,32'd-289,32'd864,32'd55,32'd949,32'd4653,32'd-4099,32'd-3178,32'd1357,32'd3518,32'd-2934,32'd6010,32'd2863,32'd5053,32'd2541,32'd2902,32'd2910,32'd121,32'd1427,32'd4167,32'd1191,32'd4345,32'd-1450,32'd-3034,32'd974,32'd1113,32'd-3427,32'd-798,32'd1842,32'd3229,32'd1470,32'd-5004,32'd-2252,32'd-2030,32'd-203,32'd4853,32'd-4509,32'd3112,32'd1716,32'd-16904,32'd1618,32'd-10849,32'd-153,32'd-525,32'd-9736,32'd-1772,32'd1375,32'd-7495,32'd10019,32'd-1159,32'd-5668,32'd5849,32'd1850,32'd-10185,32'd-4418,32'd-2590,32'd7016,32'd-1760,32'd-2932,32'd-1496,32'd-1520,32'd1290,32'd-3054,32'd-2003,32'd5458,32'd-7290,32'd6831,32'd-11650,32'd3247,32'd-3339,32'd-2687,32'd7880,32'd-1806,32'd495,32'd4331,32'd1066,32'd7133,32'd-5024,32'd-2272,32'd3430,32'd1408,32'd-4482,32'd-13505,32'd6875,32'd15703,32'd-1910,32'd-5195,32'd-3415,32'd11914,32'd-8071,32'd-219,32'd-5195,32'd6152,32'd17441,32'd-812,32'd-2165,32'd14238,32'd200,32'd-7275,32'd-6445,32'd-1054,32'd-4321,32'd9921,32'd1202,32'd1962,32'd-639,32'd2415,32'd-2685,32'd-2153,32'd3515,32'd3811,32'd5927,32'd289,32'd-1160,32'd-8359,32'd2219,32'd4726,32'd-1771,32'd-2268,32'd11835,32'd-1088,32'd-22050,32'd-5463,32'd4274,32'd501,32'd5888,32'd6621,32'd3642,32'd7758,32'd9057,32'd-1206,32'd-1191,32'd-786,32'd3354,32'd-6254,32'd-734,32'd286,32'd-3400,32'd1920,32'd7353,32'd-5380,32'd3149,32'd3090,32'd-606,32'd-1562,32'd-9130,32'd-4060,32'd335,32'd-6933,32'd4270,32'd5107,32'd-4475,32'd-2841,32'd-10244,32'd3967,32'd1176,32'd-2116,32'd-645,32'd-2187,32'd-3059,32'd-380,32'd2150,32'd-5371,32'd1861,32'd995,32'd1607,32'd-327,32'd255,32'd7661,32'd-5244,32'd-5029,32'd-93,32'd-3627,32'd1618,32'd914,32'd-2727,32'd-9770,32'd-4587,32'd-1343,32'd-667,32'd-9165,32'd-4455,32'd-8569,32'd-4094,32'd4853,32'd-6743,32'd3869,32'd-1293,32'd-6708,32'd-1270,32'd-6884,32'd-4091,32'd2780,32'd-6396,32'd-2185,32'd1628,32'd112,32'd-2944,32'd-1594,32'd-2971,32'd-3520,32'd2558,32'd-13710,32'd-3774,32'd-2939,32'd-331,32'd-2148,32'd-5214,32'd-471,32'd-4260,32'd-222,32'd-7080,32'd-770,32'd-3688,32'd1259,32'd-530,32'd5498,32'd-4948,32'd-3195,32'd11396,32'd-9199,32'd601,32'd-4140,32'd-5234,32'd-1246,32'd-3630,32'd2420,32'd2624,32'd1940,32'd-1459,32'd-1033,32'd-6933,32'd-2629,32'd-3991,32'd-4370,32'd-336,32'd-4501,32'd-787,32'd1201,32'd4519,32'd-6552,32'd5546,32'd2963,32'd-2097,32'd-726,32'd-8105,32'd-2929,32'd160,32'd-653,32'd1661,32'd3745,32'd-4782,32'd-1354,32'd-4995,32'd4604,32'd310,32'd-4782,32'd526,32'd2705,32'd-130,32'd1973,32'd256,32'd-3112,32'd1597,32'd-7216,32'd-789,32'd6923,32'd-955,32'd10585,32'd1278,32'd8076,32'd2971,32'd-7475,32'd3933,32'd-692,32'd-3271,32'd1893,32'd7124,32'd-2312,32'd3122,32'd2495,32'd321,32'd3388,32'd-5185,32'd-3193,32'd1823,32'd977,32'd-1619,32'd-670,32'd-1568,32'd216,32'd2437,32'd-10683,32'd5698,32'd-2313,32'd5375,32'd245,32'd5952,32'd9208,32'd-2722,32'd6425,32'd273,32'd-177,32'd917,32'd-10498,32'd-241,32'd-7011,32'd-1696,32'd-1109,32'd12304,32'd-214,32'd107,32'd-3840,32'd1613,32'd4978,32'd-1551,32'd2868,32'd-8808,32'd-7363,32'd564,32'd-1928,32'd5410,32'd-13085,32'd-8564,32'd373,32'd-2440,32'd6665,32'd2687,32'd-6059,32'd3581,32'd-3989,32'd-2788,32'd304,32'd-3464,32'd-8354,32'd1101,32'd-6972,32'd2641};
    Wx[74]='{32'd702,32'd5625,32'd-3049,32'd759,32'd1800,32'd394,32'd61,32'd1231,32'd-4592,32'd-1390,32'd-253,32'd-2419,32'd1702,32'd7060,32'd-1276,32'd-4418,32'd-3146,32'd-1518,32'd1401,32'd-1701,32'd-1296,32'd2038,32'd2326,32'd1481,32'd-2287,32'd798,32'd-2849,32'd-1292,32'd540,32'd-1978,32'd2326,32'd-5336,32'd-883,32'd4226,32'd-5219,32'd-3017,32'd3950,32'd-522,32'd-5156,32'd-5097,32'd1557,32'd-9995,32'd6381,32'd-1119,32'd-3540,32'd-2454,32'd-4160,32'd-6132,32'd-2297,32'd1774,32'd-4682,32'd4577,32'd-3652,32'd-3957,32'd-1473,32'd-3415,32'd-1145,32'd-1682,32'd-2966,32'd-5234,32'd-1223,32'd-4174,32'd-474,32'd-2646,32'd-2595,32'd235,32'd-3271,32'd-8159,32'd2019,32'd1822,32'd-718,32'd-12363,32'd3911,32'd-3454,32'd1335,32'd4941,32'd-8417,32'd-4379,32'd3437,32'd-3723,32'd2739,32'd-8730,32'd-337,32'd-3515,32'd-874,32'd931,32'd-4228,32'd12,32'd3112,32'd1420,32'd-789,32'd-6728,32'd-3935,32'd-3698,32'd1328,32'd1226,32'd1392,32'd-4785,32'd899,32'd620,32'd-1475,32'd812,32'd-2276,32'd-16669,32'd1704,32'd-1274,32'd4870,32'd3632,32'd7084,32'd6088,32'd-13505,32'd-1535,32'd4199,32'd-4807,32'd14658,32'd5346,32'd2066,32'd-9379,32'd-96,32'd2871,32'd1619,32'd4699,32'd-13505,32'd-545,32'd3017,32'd2558,32'd-8110,32'd2783,32'd10097,32'd1477,32'd-10712,32'd-4992,32'd8593,32'd7846,32'd-2802,32'd1170,32'd-1988,32'd-2381,32'd-10517,32'd3339,32'd751,32'd-7089,32'd5112,32'd218,32'd-10566,32'd-9287,32'd6904,32'd294,32'd4665,32'd364,32'd11748,32'd-5869,32'd-6079,32'd3388,32'd-2819,32'd2489,32'd-6713,32'd-1639,32'd-5966,32'd429,32'd-1356,32'd-1154,32'd4929,32'd6791,32'd-8876,32'd-70,32'd-874,32'd9125,32'd2369,32'd-814,32'd1630,32'd5268,32'd-2127,32'd5361,32'd1313,32'd-6855,32'd-7119,32'd1624,32'd22187,32'd-3549,32'd4853,32'd-2219,32'd-9394,32'd-9877,32'd2462,32'd6884,32'd-1229,32'd3828,32'd-753,32'd5996,32'd-1335,32'd8779,32'd-9018,32'd1950,32'd2197,32'd-13300,32'd5922,32'd102,32'd-1845,32'd2512,32'd-4174,32'd-2951,32'd1875,32'd343,32'd-5195,32'd969,32'd-6679,32'd-2548,32'd1024,32'd-1252,32'd5146,32'd-7285,32'd-440,32'd-2069,32'd-3037,32'd-1506,32'd-4787,32'd-2347,32'd944,32'd-2404,32'd-1893,32'd254,32'd445,32'd2641,32'd-852,32'd569,32'd-1694,32'd2010,32'd-4729,32'd1,32'd2685,32'd7158,32'd-5952,32'd945,32'd4887,32'd7070,32'd378,32'd-2415,32'd-8876,32'd2556,32'd1416,32'd-8076,32'd-6308,32'd-9155,32'd-7324,32'd-821,32'd-5488,32'd318,32'd-475,32'd539,32'd2309,32'd3608,32'd-6899,32'd-3100,32'd-527,32'd-3393,32'd2012,32'd2325,32'd-2181,32'd-1499,32'd2011,32'd2897,32'd4204,32'd8574,32'd2203,32'd6459,32'd-2138,32'd7626,32'd2279,32'd1229,32'd-6611,32'd2658,32'd-297,32'd4050,32'd-1489,32'd-3847,32'd-4660,32'd-38,32'd-5292,32'd-2963,32'd-835,32'd-3559,32'd-4675,32'd4355,32'd825,32'd-8862,32'd-4375,32'd-5336,32'd-1564,32'd4050,32'd7373,32'd-5253,32'd5761,32'd2624,32'd9882,32'd4123,32'd1563,32'd-9194,32'd-332,32'd-1131,32'd-8833,32'd-1221,32'd2524,32'd163,32'd-443,32'd2656,32'd-3925,32'd-5390,32'd-6093,32'd-186,32'd-491,32'd-903,32'd-3918,32'd-2034,32'd-6254,32'd-4916,32'd-5576,32'd-10917,32'd2543,32'd1639,32'd2512,32'd-1690,32'd2761,32'd-5507,32'd-6108,32'd6303,32'd-3676,32'd-2902,32'd-9433,32'd-2406,32'd-1345,32'd1618,32'd3518,32'd-772,32'd4719,32'd-1691,32'd6323,32'd-2333,32'd-2590,32'd-2236,32'd-3576,32'd-12138,32'd-1195,32'd-4274,32'd-7133,32'd-2122,32'd-1488,32'd-3012,32'd1752,32'd2175,32'd4953,32'd955,32'd-1911,32'd-1435,32'd693,32'd3913,32'd3403,32'd5390,32'd-658,32'd6230,32'd1221,32'd-2274,32'd-8286,32'd8237,32'd4577,32'd-919,32'd-5625,32'd270,32'd-17988,32'd-3293,32'd-6020,32'd-3864,32'd-6577,32'd-1756,32'd4509,32'd-136,32'd-2175,32'd2343,32'd2719,32'd-4587,32'd-3315,32'd-1233,32'd-4384,32'd-1939,32'd-8735,32'd-6118,32'd-9252,32'd-3715,32'd-2683,32'd893,32'd3332,32'd-10634,32'd1064,32'd1184,32'd714,32'd-3312,32'd991,32'd-9140,32'd-1265,32'd-2583};
    Wx[75]='{32'd1287,32'd1462,32'd-1331,32'd-3156,32'd856,32'd437,32'd4851,32'd-1466,32'd2785,32'd-1788,32'd-6977,32'd-2235,32'd-3457,32'd8579,32'd3178,32'd-2071,32'd-4243,32'd3708,32'd2366,32'd-1923,32'd-983,32'd-838,32'd-3100,32'd377,32'd-2883,32'd-1611,32'd-2973,32'd-2277,32'd3752,32'd2341,32'd108,32'd9199,32'd-9345,32'd-316,32'd-3864,32'd2624,32'd-5166,32'd-389,32'd-2753,32'd-225,32'd-2570,32'd-2165,32'd-1756,32'd1105,32'd-3259,32'd-4409,32'd-5664,32'd-380,32'd-813,32'd2463,32'd2119,32'd6137,32'd-2081,32'd-3376,32'd-2731,32'd-5566,32'd-2741,32'd-6005,32'd-2880,32'd-4458,32'd5112,32'd-2985,32'd789,32'd-1655,32'd-5546,32'd-239,32'd-3952,32'd-2883,32'd-102,32'd-1651,32'd-496,32'd-4682,32'd4980,32'd3911,32'd-5825,32'd-4404,32'd3364,32'd-458,32'd-1643,32'd-2910,32'd2248,32'd2641,32'd-4477,32'd-287,32'd1550,32'd-696,32'd-418,32'd606,32'd-731,32'd-2028,32'd480,32'd-5849,32'd-2059,32'd-1798,32'd-10605,32'd173,32'd-1915,32'd-5996,32'd634,32'd201,32'd-2807,32'd-11953,32'd-1838,32'd1357,32'd1185,32'd805,32'd1008,32'd-9433,32'd5664,32'd4685,32'd2386,32'd-2047,32'd-3271,32'd3166,32'd-4179,32'd-7680,32'd-14853,32'd-6948,32'd-4587,32'd-5410,32'd-969,32'd-214,32'd5322,32'd5249,32'd-2626,32'd-606,32'd-3896,32'd7509,32'd4680,32'd-4291,32'd3422,32'd6840,32'd2059,32'd3242,32'd-2946,32'd7846,32'd-3928,32'd-4455,32'd-1098,32'd-949,32'd-4042,32'd617,32'd8432,32'd3303,32'd-5698,32'd5375,32'd8730,32'd-257,32'd-4101,32'd2230,32'd-5947,32'd23125,32'd-5107,32'd10732,32'd418,32'd941,32'd-5195,32'd-3662,32'd20,32'd-1651,32'd-8666,32'd4077,32'd-6303,32'd-520,32'd7719,32'd2705,32'd5317,32'd-510,32'd75,32'd-3513,32'd1218,32'd-5917,32'd-901,32'd4770,32'd-2666,32'd1092,32'd-3571,32'd2457,32'd-4265,32'd-144,32'd6416,32'd-5478,32'd-826,32'd9833,32'd3652,32'd1685,32'd1531,32'd-3730,32'd-1264,32'd-2304,32'd-4052,32'd5937,32'd4353,32'd2297,32'd4936,32'd3601,32'd12714,32'd-6547,32'd-1574,32'd-3149,32'd-93,32'd-10898,32'd2731,32'd-1236,32'd-2379,32'd902,32'd-3808,32'd-489,32'd-3117,32'd-3188,32'd262,32'd5190,32'd1103,32'd-119,32'd-411,32'd2985,32'd8432,32'd-3107,32'd-874,32'd3161,32'd1210,32'd3103,32'd-3750,32'd1771,32'd1914,32'd-2595,32'd-489,32'd-4143,32'd9189,32'd-2500,32'd3740,32'd10751,32'd1788,32'd3278,32'd3017,32'd-47,32'd2121,32'd2939,32'd6611,32'd-380,32'd3225,32'd-8818,32'd8784,32'd-3522,32'd4558,32'd5581,32'd3669,32'd-6196,32'd-2954,32'd4340,32'd-2641,32'd-8237,32'd-2663,32'd-690,32'd4172,32'd1156,32'd-5971,32'd-881,32'd-4663,32'd1557,32'd-196,32'd-127,32'd-1895,32'd949,32'd6586,32'd2316,32'd2519,32'd9472,32'd-2075,32'd-965,32'd3967,32'd1098,32'd-788,32'd-4982,32'd-4755,32'd643,32'd-469,32'd4816,32'd5634,32'd-2249,32'd2413,32'd-809,32'd-1752,32'd-1223,32'd571,32'd2512,32'd-2412,32'd1510,32'd-7221,32'd-1215,32'd-673,32'd4267,32'd-6948,32'd-2326,32'd-6308,32'd422,32'd373,32'd3315,32'd-3352,32'd3142,32'd-4619,32'd-9794,32'd3146,32'd2731,32'd-3181,32'd-13720,32'd-380,32'd-8515,32'd-2832,32'd-2617,32'd1275,32'd744,32'd-6484,32'd-5620,32'd-4523,32'd-62,32'd4519,32'd3937,32'd650,32'd-6811,32'd-15039,32'd-600,32'd-2563,32'd1198,32'd-1303,32'd2565,32'd-346,32'd-10097,32'd-2597,32'd515,32'd-91,32'd47,32'd-5517,32'd-5747,32'd1724,32'd2573,32'd2844,32'd-9326,32'd173,32'd6430,32'd-2963,32'd-4948,32'd-1547,32'd5478,32'd9018,32'd3786,32'd-6723,32'd2875,32'd-4904,32'd5947,32'd5444,32'd800,32'd-83,32'd-3056,32'd4846,32'd-2019,32'd-9238,32'd-1473,32'd-3662,32'd-4919,32'd4653,32'd-1216,32'd1428,32'd-999,32'd2490,32'd3867,32'd-6450,32'd1282,32'd1448,32'd-11250,32'd4841,32'd-3256,32'd-214,32'd8339,32'd-3962,32'd-5781,32'd-3984,32'd2646,32'd4013,32'd-6464,32'd2452,32'd-2648,32'd2257,32'd-4599,32'd2375,32'd6962,32'd-4035,32'd3903,32'd-2086,32'd-6572,32'd4572,32'd-1483,32'd290,32'd-822,32'd-3815,32'd1275,32'd2626,32'd-3640,32'd-5317,32'd-607};
    Wx[76]='{32'd944,32'd3081,32'd-39,32'd-1276,32'd-4479,32'd-3771,32'd3623,32'd-498,32'd1793,32'd-2543,32'd-225,32'd1026,32'd844,32'd-3015,32'd1488,32'd856,32'd723,32'd6479,32'd3107,32'd-2193,32'd-3750,32'd-4174,32'd3627,32'd-83,32'd2008,32'd1608,32'd58,32'd-226,32'd-7207,32'd-2159,32'd2165,32'd1499,32'd-3825,32'd5268,32'd-5668,32'd-4895,32'd2292,32'd1337,32'd20,32'd-1189,32'd-1070,32'd-1339,32'd-764,32'd2827,32'd2670,32'd1842,32'd-273,32'd2592,32'd1140,32'd-213,32'd-1755,32'd2373,32'd-9,32'd1373,32'd-430,32'd4565,32'd-1284,32'd-819,32'd-1162,32'd1634,32'd1435,32'd-1811,32'd-527,32'd2413,32'd4069,32'd-947,32'd83,32'd3754,32'd-2474,32'd1188,32'd-1284,32'd-448,32'd-4831,32'd-2386,32'd-1104,32'd2286,32'd264,32'd412,32'd-116,32'd-2509,32'd-3300,32'd14677,32'd-1636,32'd6865,32'd895,32'd4077,32'd-5629,32'd-1604,32'd-375,32'd-4626,32'd1060,32'd6430,32'd173,32'd-5166,32'd2585,32'd-2863,32'd-1140,32'd1984,32'd3439,32'd5346,32'd5922,32'd-213,32'd1313,32'd-2110,32'd354,32'd2205,32'd-4699,32'd-7646,32'd-1645,32'd-134,32'd9956,32'd-4746,32'd1682,32'd12402,32'd-14990,32'd-7045,32'd5117,32'd7373,32'd-1599,32'd-387,32'd-3444,32'd-6088,32'd-1915,32'd6152,32'd3732,32'd1835,32'd-3503,32'd-5371,32'd-11093,32'd-5957,32'd-6547,32'd2763,32'd1084,32'd6313,32'd-4692,32'd3889,32'd1069,32'd4089,32'd15468,32'd-16435,32'd-7758,32'd-16240,32'd-9262,32'd-7016,32'd2373,32'd-681,32'd-481,32'd-13789,32'd-5131,32'd289,32'd17265,32'd15117,32'd265,32'd-14208,32'd6044,32'd7739,32'd3901,32'd1335,32'd1412,32'd-1948,32'd-7036,32'd-2242,32'd-1508,32'd6298,32'd4306,32'd4077,32'd-952,32'd-8730,32'd-3684,32'd-433,32'd11044,32'd-10654,32'd-2303,32'd6552,32'd1195,32'd5268,32'd9604,32'd-11630,32'd12070,32'd-5585,32'd-2651,32'd-10390,32'd6586,32'd6577,32'd-426,32'd-5961,32'd9243,32'd11992,32'd-2396,32'd-428,32'd2741,32'd1346,32'd-6518,32'd5039,32'd-8007,32'd3291,32'd4294,32'd-4909,32'd4011,32'd-4838,32'd2198,32'd4370,32'd823,32'd-5009,32'd-102,32'd-128,32'd-780,32'd731,32'd-1271,32'd-1660,32'd-5927,32'd-5141,32'd-774,32'd-4094,32'd8608,32'd997,32'd302,32'd-294,32'd3835,32'd-5473,32'd2770,32'd4333,32'd-2135,32'd2116,32'd-4675,32'd1884,32'd3603,32'd-612,32'd-7207,32'd-1000,32'd-1024,32'd-1220,32'd2812,32'd-7509,32'd2209,32'd-2507,32'd-133,32'd538,32'd-3466,32'd-4660,32'd2390,32'd4592,32'd4306,32'd-5004,32'd-1275,32'd-2456,32'd2249,32'd861,32'd4348,32'd-1156,32'd-720,32'd-5673,32'd2023,32'd442,32'd-371,32'd11259,32'd422,32'd2220,32'd130,32'd-631,32'd4311,32'd3657,32'd-1960,32'd-3881,32'd1926,32'd-6372,32'd-1506,32'd3398,32'd-175,32'd4145,32'd-955,32'd-5024,32'd-186,32'd-3823,32'd-1440,32'd4545,32'd2452,32'd-8242,32'd9125,32'd-2895,32'd333,32'd-4213,32'd-5375,32'd-6562,32'd2204,32'd-3925,32'd24,32'd-3564,32'd1292,32'd-2504,32'd3532,32'd-1139,32'd-141,32'd2666,32'd-7558,32'd-2502,32'd-7446,32'd-6572,32'd3347,32'd-3078,32'd-4089,32'd4689,32'd-1859,32'd579,32'd-2185,32'd-3425,32'd5366,32'd9033,32'd-1540,32'd3146,32'd-7167,32'd-4790,32'd-4675,32'd-357,32'd-488,32'd-3093,32'd-3024,32'd5170,32'd1029,32'd-3642,32'd174,32'd1783,32'd1218,32'd2644,32'd484,32'd4062,32'd4538,32'd-3330,32'd-9272,32'd109,32'd920,32'd1211,32'd-3520,32'd2644,32'd-5224,32'd-2541,32'd-4560,32'd6738,32'd4064,32'd-6938,32'd374,32'd1227,32'd5092,32'd-1328,32'd5732,32'd-82,32'd-7148,32'd-7114,32'd4738,32'd3127,32'd-3598,32'd-7700,32'd5063,32'd4467,32'd10693,32'd-3061,32'd1120,32'd161,32'd2196,32'd-1430,32'd7392,32'd-1639,32'd2453,32'd80,32'd4609,32'd-455,32'd-8554,32'd4621,32'd9799,32'd1550,32'd-859,32'd1232,32'd3022,32'd-4384,32'd-825,32'd7709,32'd-1480,32'd-4775,32'd1195,32'd-4055,32'd-718,32'd-4926,32'd-7998,32'd-908,32'd11435,32'd932,32'd-9643,32'd-2269,32'd-654,32'd477,32'd1414,32'd-7407,32'd3061,32'd2727,32'd-1445,32'd-1611,32'd3574,32'd1945,32'd4758,32'd-756};
    Wx[77]='{32'd-2631,32'd-3928,32'd-2156,32'd-1724,32'd-406,32'd-1066,32'd-1110,32'd-2427,32'd3356,32'd-3173,32'd9072,32'd-225,32'd2479,32'd-4316,32'd-6074,32'd3867,32'd3969,32'd1252,32'd-4560,32'd893,32'd3632,32'd-623,32'd-2912,32'd-479,32'd-2416,32'd-3176,32'd-1271,32'd-1341,32'd3764,32'd1818,32'd2712,32'd-1188,32'd-5346,32'd1734,32'd-3493,32'd-801,32'd2507,32'd-5253,32'd296,32'd-2418,32'd-4101,32'd-5292,32'd1128,32'd-7944,32'd2476,32'd2268,32'd1921,32'd-1444,32'd466,32'd-1617,32'd2770,32'd1762,32'd3032,32'd1007,32'd3164,32'd-2832,32'd-371,32'd3132,32'd-2181,32'd-594,32'd-3244,32'd-7934,32'd743,32'd1464,32'd2976,32'd2326,32'd-3725,32'd4855,32'd-4174,32'd-1403,32'd5146,32'd-3120,32'd-1071,32'd-3405,32'd4479,32'd-3444,32'd1958,32'd-1298,32'd-147,32'd-1828,32'd112,32'd5439,32'd-3549,32'd4609,32'd-1319,32'd1905,32'd-664,32'd2687,32'd-546,32'd5219,32'd-16,32'd-9370,32'd-8662,32'd4333,32'd-3708,32'd-1959,32'd1784,32'd-470,32'd-5043,32'd-5229,32'd1014,32'd2497,32'd936,32'd-6694,32'd-8881,32'd1776,32'd123,32'd-6879,32'd-2121,32'd-2602,32'd17294,32'd-1978,32'd-7724,32'd-8652,32'd7509,32'd-4311,32'd-6611,32'd-318,32'd4682,32'd4946,32'd-291,32'd1273,32'd-550,32'd2495,32'd-4248,32'd-8945,32'd-2401,32'd-2770,32'd7480,32'd-3967,32'd8676,32'd2124,32'd-10634,32'd20273,32'd2086,32'd-1617,32'd-6098,32'd-4289,32'd5371,32'd14804,32'd4863,32'd-1931,32'd-5883,32'd4650,32'd-8681,32'd-9609,32'd-3310,32'd3317,32'd5981,32'd-5908,32'd-19423,32'd-8378,32'd-7993,32'd419,32'd-2929,32'd9926,32'd13183,32'd-927,32'd-534,32'd-5537,32'd-2639,32'd-11806,32'd-822,32'd-4587,32'd4924,32'd-487,32'd-1768,32'd8359,32'd-2099,32'd538,32'd5297,32'd5493,32'd-1143,32'd-9858,32'd3942,32'd-19902,32'd-3879,32'd4624,32'd-1535,32'd3354,32'd-6235,32'd1999,32'd-1613,32'd-10302,32'd111,32'd8608,32'd-6826,32'd6171,32'd-492,32'd1785,32'd9487,32'd24199,32'd2912,32'd-471,32'd-5854,32'd4438,32'd-6362,32'd-16162,32'd-8808,32'd-6367,32'd5395,32'd-988,32'd-2258,32'd264,32'd5048,32'd-657,32'd-955,32'd5053,32'd1391,32'd3793,32'd3796,32'd-341,32'd2749,32'd6274,32'd2440,32'd4309,32'd1331,32'd1380,32'd-2890,32'd7084,32'd-3056,32'd-180,32'd2561,32'd-1491,32'd339,32'd1116,32'd7832,32'd682,32'd11914,32'd3911,32'd-531,32'd-6333,32'd4511,32'd8481,32'd-1884,32'd-153,32'd-3830,32'd-145,32'd-1507,32'd-4543,32'd1949,32'd1123,32'd5747,32'd1155,32'd9184,32'd819,32'd14882,32'd9985,32'd4584,32'd-1336,32'd-4040,32'd2712,32'd-3718,32'd-13632,32'd2802,32'd-1,32'd2053,32'd-1149,32'd3891,32'd-6430,32'd217,32'd2551,32'd-3044,32'd-8403,32'd-3222,32'd677,32'd-376,32'd7026,32'd-322,32'd-309,32'd-7812,32'd2644,32'd419,32'd-435,32'd3559,32'd2136,32'd-2125,32'd2498,32'd-2023,32'd123,32'd1021,32'd-6044,32'd-4089,32'd6367,32'd7241,32'd-3037,32'd4116,32'd2369,32'd184,32'd108,32'd-4304,32'd174,32'd817,32'd3015,32'd13623,32'd1439,32'd-349,32'd19199,32'd-3991,32'd1217,32'd1335,32'd1420,32'd-14980,32'd-3806,32'd2917,32'd-2661,32'd-1015,32'd6982,32'd-7309,32'd-155,32'd7216,32'd-1711,32'd4787,32'd-2773,32'd5937,32'd-3808,32'd1658,32'd-4150,32'd-1386,32'd-6787,32'd5913,32'd3195,32'd-1296,32'd-1064,32'd812,32'd596,32'd1018,32'd-2863,32'd8081,32'd2196,32'd-3027,32'd-5092,32'd2432,32'd-3085,32'd-3154,32'd-1065,32'd-2130,32'd-56,32'd4665,32'd-2529,32'd-6469,32'd-4873,32'd2172,32'd5932,32'd2225,32'd520,32'd1761,32'd31,32'd7094,32'd-1645,32'd-4909,32'd-4550,32'd-16103,32'd-5351,32'd4887,32'd5932,32'd2985,32'd-8193,32'd-7504,32'd-8935,32'd-3286,32'd-1975,32'd2384,32'd-3337,32'd-2692,32'd490,32'd-7910,32'd2824,32'd-10078,32'd-5009,32'd-1947,32'd-2729,32'd-1531,32'd3356,32'd4890,32'd3576,32'd2575,32'd-4047,32'd-403,32'd-3791,32'd-1451,32'd-3022,32'd-4719,32'd7480,32'd6669,32'd-6240,32'd1700,32'd345,32'd-1628,32'd-8369,32'd-514,32'd2282,32'd-3630,32'd-3024,32'd9965,32'd246,32'd-4914,32'd2148,32'd-2412,32'd-4775};
    Wx[78]='{32'd-2902,32'd-3862,32'd-4235,32'd4418,32'd-960,32'd1879,32'd-1754,32'd-624,32'd-2568,32'd893,32'd-3310,32'd-1163,32'd-2014,32'd2470,32'd-295,32'd-1402,32'd-6352,32'd-752,32'd-5791,32'd-760,32'd-2000,32'd-552,32'd-4287,32'd-239,32'd-4863,32'd-3798,32'd1392,32'd-1132,32'd-1882,32'd-2770,32'd-1090,32'd-4611,32'd6337,32'd-561,32'd56,32'd-1932,32'd-4738,32'd1553,32'd-3447,32'd3056,32'd-4018,32'd-5029,32'd-3364,32'd-3847,32'd-10029,32'd-40,32'd2484,32'd574,32'd4399,32'd2885,32'd3596,32'd-2858,32'd1523,32'd-2761,32'd-4978,32'd-4375,32'd-3723,32'd-762,32'd-1497,32'd-1341,32'd-7827,32'd810,32'd-1009,32'd-5234,32'd-3063,32'd6137,32'd-1892,32'd-3859,32'd447,32'd191,32'd-4128,32'd-617,32'd-3933,32'd-953,32'd645,32'd-9301,32'd1125,32'd-213,32'd4746,32'd334,32'd1335,32'd7329,32'd2144,32'd3122,32'd6044,32'd-4421,32'd-287,32'd3554,32'd96,32'd917,32'd-1076,32'd3901,32'd-7470,32'd6533,32'd-3725,32'd-1398,32'd-3708,32'd-3608,32'd-1492,32'd-3344,32'd-4533,32'd-8496,32'd-504,32'd2683,32'd-3789,32'd-2324,32'd-4030,32'd14082,32'd2932,32'd-1060,32'd-9111,32'd-313,32'd8129,32'd-10224,32'd-2071,32'd-6059,32'd7539,32'd1397,32'd5034,32'd572,32'd-908,32'd-2468,32'd4602,32'd-10273,32'd-10605,32'd-6958,32'd4038,32'd-993,32'd-32,32'd127,32'd-1768,32'd-9980,32'd5107,32'd15839,32'd389,32'd-3608,32'd-5595,32'd-3122,32'd5839,32'd2905,32'd2900,32'd-4050,32'd3354,32'd-4611,32'd-14472,32'd12216,32'd3205,32'd4804,32'd-2427,32'd-2440,32'd2399,32'd-4140,32'd-2309,32'd4079,32'd-1201,32'd6040,32'd-7768,32'd-2211,32'd-9223,32'd-1320,32'd-432,32'd6860,32'd457,32'd1130,32'd9252,32'd-2978,32'd-1187,32'd-3937,32'd2075,32'd-2631,32'd-4245,32'd11982,32'd4536,32'd-1279,32'd3364,32'd972,32'd-6743,32'd10234,32'd10947,32'd9165,32'd-127,32'd7968,32'd-4199,32'd-5234,32'd3430,32'd2641,32'd-4584,32'd12568,32'd7563,32'd2100,32'd-4475,32'd8085,32'd5136,32'd817,32'd-15664,32'd877,32'd524,32'd-20332,32'd-6206,32'd-4055,32'd1297,32'd5454,32'd-2391,32'd1044,32'd7080,32'd-95,32'd759,32'd-7485,32'd505,32'd2319,32'd4216,32'd-4584,32'd-8261,32'd2985,32'd1269,32'd-874,32'd3291,32'd5498,32'd-7871,32'd-92,32'd-689,32'd-184,32'd-4077,32'd-914,32'd-2174,32'd-942,32'd1335,32'd75,32'd5815,32'd2152,32'd6508,32'd-5249,32'd2083,32'd8554,32'd4396,32'd-1676,32'd12001,32'd7211,32'd-4060,32'd-3803,32'd10322,32'd665,32'd13750,32'd1634,32'd-1951,32'd5019,32'd-22226,32'd-2392,32'd-2248,32'd6586,32'd-4282,32'd3083,32'd-1778,32'd-2478,32'd2006,32'd13925,32'd-3515,32'd5908,32'd6176,32'd-1816,32'd2890,32'd3459,32'd6503,32'd-2238,32'd8789,32'd3632,32'd-226,32'd-12509,32'd1955,32'd-932,32'd-1918,32'd2346,32'd-1975,32'd-9638,32'd1343,32'd-2246,32'd6669,32'd-618,32'd1436,32'd5195,32'd941,32'd-1827,32'd281,32'd-3840,32'd3378,32'd7827,32'd-930,32'd1591,32'd-32,32'd2309,32'd4702,32'd-2761,32'd276,32'd6430,32'd841,32'd252,32'd952,32'd10400,32'd-3447,32'd10048,32'd6826,32'd5751,32'd4162,32'd2722,32'd8823,32'd1221,32'd-1287,32'd-6899,32'd-4196,32'd-6909,32'd906,32'd-3725,32'd-2631,32'd6005,32'd-502,32'd-5844,32'd1688,32'd-3156,32'd-2836,32'd2917,32'd3081,32'd3029,32'd-645,32'd1922,32'd-2384,32'd-2082,32'd3264,32'd2308,32'd7910,32'd-2512,32'd5874,32'd-4729,32'd1058,32'd5122,32'd-2504,32'd3881,32'd1669,32'd5380,32'd335,32'd3442,32'd235,32'd-771,32'd3569,32'd8774,32'd-2783,32'd2213,32'd-9350,32'd-1513,32'd14873,32'd-4074,32'd-5166,32'd-823,32'd1711,32'd2319,32'd2034,32'd7939,32'd-3483,32'd3764,32'd-492,32'd-3605,32'd-3349,32'd-2199,32'd3310,32'd-1796,32'd-371,32'd3461,32'd-912,32'd761,32'd-7241,32'd-10302,32'd-2410,32'd-5024,32'd-5361,32'd-6303,32'd582,32'd-2517,32'd7021,32'd2187,32'd-199,32'd881,32'd-2873,32'd-3806,32'd-1384,32'd-1641,32'd5058,32'd7822,32'd-696,32'd-3085,32'd-2670,32'd4465,32'd-3366,32'd839,32'd-2369,32'd6801,32'd5683,32'd56,32'd4604,32'd1113,32'd-12001,32'd5307};
    Wx[79]='{32'd1622,32'd-254,32'd-1959,32'd1168,32'd3474,32'd-953,32'd-7631,32'd-462,32'd16,32'd-142,32'd5390,32'd2410,32'd4411,32'd-3315,32'd2592,32'd4172,32'd-2131,32'd4338,32'd3051,32'd-1019,32'd791,32'd2324,32'd376,32'd-2421,32'd2766,32'd1188,32'd1187,32'd-572,32'd2639,32'd-1076,32'd-962,32'd4089,32'd-4228,32'd339,32'd3232,32'd1611,32'd5805,32'd-5151,32'd1141,32'd1087,32'd1833,32'd2321,32'd2626,32'd3735,32'd3488,32'd-757,32'd-1818,32'd3649,32'd4721,32'd1993,32'd1644,32'd-6030,32'd-285,32'd1328,32'd-1721,32'd8901,32'd-1239,32'd-4592,32'd6855,32'd8457,32'd3959,32'd-1630,32'd4758,32'd3959,32'd3564,32'd2447,32'd4504,32'd-4885,32'd4152,32'd3425,32'd5527,32'd7480,32'd1695,32'd-4125,32'd-117,32'd877,32'd2496,32'd-2144,32'd-884,32'd1734,32'd-2244,32'd-1501,32'd-1680,32'd2998,32'd2983,32'd-1470,32'd2668,32'd-2934,32'd6391,32'd819,32'd-2467,32'd-6474,32'd-2041,32'd3576,32'd2534,32'd5361,32'd442,32'd-3791,32'd-2143,32'd3125,32'd-1015,32'd6284,32'd2357,32'd-973,32'd11542,32'd2341,32'd2349,32'd6132,32'd760,32'd3205,32'd-16103,32'd-3066,32'd-5141,32'd-17314,32'd8369,32'd-6708,32'd-17119,32'd-8666,32'd2712,32'd361,32'd-1055,32'd123,32'd-2675,32'd808,32'd419,32'd5766,32'd-6020,32'd-4179,32'd5610,32'd-3430,32'd-11484,32'd-13369,32'd1242,32'd-4257,32'd1433,32'd9326,32'd3291,32'd-3188,32'd-9931,32'd1911,32'd-2413,32'd1654,32'd-5517,32'd4636,32'd-570,32'd1312,32'd-1612,32'd-485,32'd9692,32'd-1778,32'd-3271,32'd5312,32'd2006,32'd9125,32'd-1959,32'd-4956,32'd-750,32'd3706,32'd-4118,32'd-209,32'd-62,32'd-16484,32'd-2397,32'd300,32'd-10488,32'd-1524,32'd-3820,32'd-10585,32'd1020,32'd745,32'd679,32'd-3281,32'd-1262,32'd517,32'd162,32'd4326,32'd-2478,32'd-3669,32'd4868,32'd-1618,32'd-217,32'd836,32'd-2308,32'd17373,32'd-7358,32'd-8471,32'd-1204,32'd-7724,32'd-8886,32'd-1085,32'd-4118,32'd9018,32'd2163,32'd-2880,32'd12431,32'd2507,32'd3532,32'd-6181,32'd-274,32'd6157,32'd-2622,32'd15205,32'd-1568,32'd-2595,32'd262,32'd-1807,32'd3105,32'd2006,32'd2934,32'd-75,32'd-1391,32'd-1754,32'd-112,32'd-270,32'd8310,32'd-457,32'd-2595,32'd-8735,32'd136,32'd826,32'd328,32'd7724,32'd2629,32'd2724,32'd289,32'd-4409,32'd-2081,32'd153,32'd909,32'd-1052,32'd1650,32'd-9194,32'd-3447,32'd-1254,32'd1898,32'd1354,32'd-2985,32'd-2966,32'd-1306,32'd2954,32'd-1271,32'd2949,32'd5224,32'd2248,32'd6440,32'd2398,32'd-404,32'd-3393,32'd983,32'd2150,32'd-1137,32'd-16220,32'd-877,32'd-440,32'd-3330,32'd-4191,32'd2171,32'd-895,32'd-2624,32'd-6435,32'd3100,32'd-677,32'd-2954,32'd-8134,32'd4426,32'd-2314,32'd3415,32'd3117,32'd-2087,32'd-118,32'd922,32'd-704,32'd-608,32'd-3947,32'd861,32'd3488,32'd-7973,32'd-81,32'd1019,32'd-5507,32'd-1357,32'd-13671,32'd-2583,32'd-4296,32'd3503,32'd11865,32'd865,32'd1072,32'd1430,32'd-3591,32'd983,32'd-3676,32'd3532,32'd-4072,32'd-14042,32'd3205,32'd3928,32'd-5087,32'd3625,32'd-6416,32'd149,32'd4426,32'd-10429,32'd-1937,32'd3513,32'd5292,32'd-2197,32'd-1361,32'd3923,32'd1225,32'd-1450,32'd3186,32'd-5249,32'd-9501,32'd-4184,32'd-2683,32'd383,32'd-5424,32'd4816,32'd-999,32'd2617,32'd4157,32'd-1188,32'd-4130,32'd-2670,32'd-3100,32'd2680,32'd1671,32'd-3417,32'd-4667,32'd-4792,32'd-3249,32'd-1121,32'd-708,32'd-4218,32'd2091,32'd5288,32'd580,32'd127,32'd4992,32'd964,32'd-9335,32'd10644,32'd-7377,32'd1528,32'd7509,32'd7114,32'd5766,32'd4951,32'd-3295,32'd-4655,32'd-8051,32'd-4230,32'd3408,32'd6083,32'd4301,32'd5590,32'd1973,32'd1078,32'd5756,32'd5268,32'd2841,32'd-12187,32'd1525,32'd2495,32'd3129,32'd10429,32'd-12792,32'd-5556,32'd2580,32'd2512,32'd-2658,32'd624,32'd1185,32'd7255,32'd-92,32'd4226,32'd-2292,32'd-7871,32'd-1622,32'd-1833,32'd-9091,32'd-3259,32'd-9687,32'd-5327,32'd-299,32'd3273,32'd4157,32'd3920,32'd-2751,32'd5214,32'd-5454,32'd2379,32'd4155,32'd-4760,32'd3576,32'd1351,32'd6176,32'd5893,32'd-6391};
    Wx[80]='{32'd725,32'd4389,32'd-338,32'd-2003,32'd-1462,32'd-491,32'd-631,32'd2861,32'd-423,32'd-1601,32'd-2094,32'd-956,32'd2482,32'd4260,32'd-7973,32'd7436,32'd-1065,32'd-1569,32'd-4497,32'd232,32'd1081,32'd809,32'd-714,32'd-2651,32'd18,32'd434,32'd728,32'd1789,32'd-2287,32'd3447,32'd1683,32'd8813,32'd4812,32'd-1901,32'd-2368,32'd-3186,32'd1405,32'd99,32'd4360,32'd3159,32'd715,32'd1157,32'd-5200,32'd2342,32'd-2457,32'd6865,32'd-3469,32'd3176,32'd1209,32'd-1569,32'd-1690,32'd347,32'd3662,32'd2924,32'd2709,32'd8505,32'd-467,32'd-372,32'd717,32'd3017,32'd453,32'd2871,32'd1219,32'd1260,32'd-7714,32'd864,32'd-1818,32'd1182,32'd1450,32'd1499,32'd121,32'd5205,32'd1099,32'd-3967,32'd597,32'd1174,32'd714,32'd-154,32'd114,32'd-2729,32'd-4118,32'd-2971,32'd-841,32'd4816,32'd2177,32'd1892,32'd2578,32'd-759,32'd2885,32'd1577,32'd-6264,32'd-4372,32'd5639,32'd4902,32'd4162,32'd1881,32'd3603,32'd1005,32'd-3063,32'd7514,32'd1693,32'd-583,32'd5751,32'd632,32'd-4213,32'd1190,32'd391,32'd-1809,32'd-597,32'd11123,32'd-998,32'd-6572,32'd169,32'd-7954,32'd808,32'd-6074,32'd-3757,32'd1328,32'd1745,32'd-852,32'd1408,32'd4936,32'd-1350,32'd-2338,32'd-872,32'd-8500,32'd935,32'd-984,32'd-9184,32'd-2406,32'd3068,32'd-8930,32'd-3386,32'd1258,32'd-3503,32'd-8583,32'd-6821,32'd5742,32'd-2634,32'd8676,32'd-4357,32'd-2827,32'd-21386,32'd-9521,32'd-1336,32'd-3293,32'd-15234,32'd-2773,32'd2221,32'd-492,32'd969,32'd-4379,32'd491,32'd426,32'd-1976,32'd502,32'd1849,32'd-2185,32'd8779,32'd-4384,32'd2426,32'd-10019,32'd7050,32'd-7729,32'd14560,32'd-4479,32'd4077,32'd-1573,32'd-2644,32'd1529,32'd18896,32'd-5937,32'd4187,32'd-28,32'd-4606,32'd-7133,32'd-7636,32'd5512,32'd9453,32'd-4123,32'd-8305,32'd-5854,32'd-221,32'd17646,32'd2391,32'd-2785,32'd-2995,32'd340,32'd-5039,32'd-639,32'd5849,32'd-5117,32'd1588,32'd1748,32'd3000,32'd7758,32'd-5708,32'd4819,32'd-7387,32'd-22050,32'd-4333,32'd-13730,32'd-2639,32'd-4294,32'd-3818,32'd-1231,32'd6435,32'd6513,32'd7875,32'd-3208,32'd-8603,32'd4316,32'd2377,32'd339,32'd9609,32'd5527,32'd9160,32'd1779,32'd-4187,32'd791,32'd2758,32'd427,32'd-2922,32'd-1800,32'd-8027,32'd-539,32'd2430,32'd567,32'd187,32'd-1752,32'd294,32'd-1231,32'd-1807,32'd-1964,32'd3046,32'd-3491,32'd5043,32'd-986,32'd1395,32'd2292,32'd-4274,32'd8437,32'd3161,32'd4287,32'd-5312,32'd-2066,32'd20644,32'd7236,32'd-1357,32'd-11142,32'd-4431,32'd-5625,32'd2286,32'd-3549,32'd3808,32'd-12070,32'd-2966,32'd-114,32'd7578,32'd993,32'd-2397,32'd-583,32'd498,32'd630,32'd3300,32'd-600,32'd-2871,32'd-3991,32'd4284,32'd1279,32'd1855,32'd8510,32'd3210,32'd-148,32'd190,32'd11630,32'd-4611,32'd579,32'd-8149,32'd471,32'd5375,32'd4431,32'd-3884,32'd266,32'd1405,32'd-76,32'd345,32'd3425,32'd4042,32'd-1152,32'd31,32'd1533,32'd4094,32'd5170,32'd1357,32'd2119,32'd-1983,32'd2565,32'd313,32'd-1174,32'd-1496,32'd-5151,32'd955,32'd3933,32'd-6225,32'd1657,32'd7050,32'd8940,32'd2846,32'd-2961,32'd-2678,32'd2829,32'd-2924,32'd-1461,32'd2802,32'd523,32'd8867,32'd-1961,32'd-10683,32'd-1894,32'd3479,32'd2301,32'd-1011,32'd-7333,32'd-2861,32'd-1228,32'd-166,32'd-1923,32'd-2484,32'd5224,32'd-315,32'd-654,32'd7177,32'd2663,32'd-6787,32'd-3918,32'd-6547,32'd410,32'd-2440,32'd-2292,32'd456,32'd828,32'd-2426,32'd2496,32'd3295,32'd-648,32'd-3400,32'd2954,32'd2697,32'd-760,32'd1375,32'd-4567,32'd4338,32'd4604,32'd-2565,32'd-14902,32'd1586,32'd-3989,32'd3671,32'd-1295,32'd-2556,32'd1855,32'd5131,32'd-7524,32'd-4899,32'd-1077,32'd-6372,32'd-6235,32'd-2797,32'd3481,32'd727,32'd774,32'd-4497,32'd-5146,32'd-7382,32'd-1700,32'd-5312,32'd3122,32'd5449,32'd-3249,32'd187,32'd614,32'd-11103,32'd1260,32'd-938,32'd-1610,32'd-6992,32'd6035,32'd3857,32'd-1021,32'd-3588,32'd2651,32'd4487,32'd5820,32'd2071,32'd5922,32'd4592,32'd1419,32'd-3054,32'd2325};
    Wx[81]='{32'd819,32'd-668,32'd-3854,32'd-614,32'd213,32'd1276,32'd-2675,32'd3793,32'd-2186,32'd-1649,32'd-877,32'd-2512,32'd-498,32'd-349,32'd3325,32'd3776,32'd2824,32'd-561,32'd2539,32'd2067,32'd2225,32'd-354,32'd-569,32'd-1164,32'd594,32'd2160,32'd2590,32'd774,32'd1364,32'd428,32'd-507,32'd-1658,32'd-1671,32'd-2814,32'd3439,32'd811,32'd1607,32'd173,32'd3688,32'd-3039,32'd-296,32'd-3500,32'd-858,32'd-8593,32'd4667,32'd-2521,32'd3747,32'd-518,32'd-872,32'd963,32'd-3747,32'd-4138,32'd-1589,32'd4995,32'd-2487,32'd-432,32'd-1372,32'd-1333,32'd-3681,32'd4099,32'd-2822,32'd-5375,32'd3505,32'd1715,32'd-4514,32'd2976,32'd217,32'd-3884,32'd-1187,32'd305,32'd-2604,32'd5083,32'd-1940,32'd2800,32'd-2851,32'd-2292,32'd-900,32'd-757,32'd-2182,32'd-795,32'd-4543,32'd-3259,32'd-2150,32'd459,32'd-3989,32'd-2435,32'd106,32'd-5166,32'd-168,32'd392,32'd-673,32'd-1242,32'd2636,32'd134,32'd-5932,32'd4167,32'd1868,32'd2114,32'd2924,32'd-3813,32'd743,32'd-3503,32'd868,32'd2822,32'd2257,32'd128,32'd-6093,32'd-6665,32'd-1243,32'd-53,32'd-9833,32'd2763,32'd-4372,32'd-4467,32'd7270,32'd561,32'd-9335,32'd2895,32'd646,32'd-5712,32'd1591,32'd-6333,32'd7148,32'd-2817,32'd2958,32'd6909,32'd2534,32'd-1887,32'd-2641,32'd-5195,32'd2563,32'd17949,32'd8437,32'd5791,32'd3361,32'd4082,32'd2529,32'd1594,32'd3559,32'd-9809,32'd1562,32'd5024,32'd-8891,32'd6840,32'd-4682,32'd7539,32'd276,32'd1367,32'd2327,32'd-4345,32'd8334,32'd-16767,32'd-1022,32'd-7192,32'd2712,32'd-2907,32'd-6513,32'd-4006,32'd3757,32'd-1805,32'd-3215,32'd1748,32'd2578,32'd1010,32'd-1405,32'd894,32'd-2934,32'd-14345,32'd3784,32'd-6015,32'd-4470,32'd7622,32'd678,32'd6049,32'd-163,32'd-3801,32'd-6782,32'd4035,32'd3183,32'd6352,32'd3583,32'd2075,32'd-6093,32'd-4802,32'd-874,32'd5312,32'd439,32'd-2403,32'd4914,32'd4631,32'd-3864,32'd4916,32'd6562,32'd-5351,32'd6689,32'd4602,32'd-158,32'd-11689,32'd4580,32'd5483,32'd-989,32'd-8437,32'd-1039,32'd98,32'd-2954,32'd2043,32'd2486,32'd-4445,32'd-1716,32'd787,32'd-4692,32'd1520,32'd3884,32'd-3339,32'd-2386,32'd3190,32'd-7836,32'd-5546,32'd838,32'd927,32'd308,32'd2629,32'd-5043,32'd1242,32'd2073,32'd-3017,32'd2415,32'd1452,32'd-2478,32'd-3430,32'd6264,32'd-5034,32'd5771,32'd-393,32'd-6308,32'd1705,32'd63,32'd2866,32'd-4914,32'd-449,32'd5942,32'd114,32'd4621,32'd7543,32'd-3947,32'd-2753,32'd-11699,32'd6176,32'd-677,32'd2242,32'd-1961,32'd802,32'd-3684,32'd-2496,32'd2484,32'd-4177,32'd-4716,32'd77,32'd-6333,32'd-2438,32'd-1861,32'd-12119,32'd-6538,32'd-2008,32'd2868,32'd-97,32'd1289,32'd283,32'd-578,32'd-2341,32'd2214,32'd-4443,32'd-4343,32'd-4143,32'd-1182,32'd-1028,32'd10068,32'd3806,32'd-97,32'd1069,32'd-4265,32'd-4577,32'd3613,32'd1466,32'd2056,32'd1821,32'd-2988,32'd-854,32'd-4570,32'd-309,32'd-1254,32'd3552,32'd-904,32'd-8662,32'd7094,32'd-6831,32'd830,32'd503,32'd-536,32'd-4545,32'd2174,32'd-4401,32'd1198,32'd2602,32'd-974,32'd3051,32'd7602,32'd-4309,32'd-9418,32'd3063,32'd-7319,32'd-569,32'd160,32'd3994,32'd-1436,32'd-4287,32'd-5019,32'd-3964,32'd1658,32'd-6333,32'd3249,32'd921,32'd-2457,32'd-702,32'd-1016,32'd-2529,32'd1147,32'd803,32'd-5332,32'd-4897,32'd-2871,32'd-9809,32'd2156,32'd-3447,32'd-5151,32'd-1110,32'd-1684,32'd808,32'd4899,32'd1899,32'd-5595,32'd-5112,32'd2424,32'd3974,32'd192,32'd-7412,32'd-10029,32'd5317,32'd8159,32'd-975,32'd602,32'd383,32'd-1386,32'd-4074,32'd7866,32'd-1864,32'd-6489,32'd517,32'd-4284,32'd747,32'd1201,32'd-5532,32'd-1842,32'd-721,32'd-28,32'd4880,32'd-573,32'd-1112,32'd-4511,32'd-2541,32'd-3254,32'd-6899,32'd-1291,32'd-3503,32'd1124,32'd-659,32'd3872,32'd1134,32'd996,32'd-6738,32'd-6113,32'd-1006,32'd2009,32'd5102,32'd413,32'd-3837,32'd-2272,32'd-2194,32'd-132,32'd7026,32'd-2078,32'd2692,32'd-8344,32'd-8745,32'd-5405,32'd2819,32'd4729,32'd1712,32'd1768,32'd-10683};
    Wx[82]='{32'd2091,32'd337,32'd3483,32'd2183,32'd-3671,32'd52,32'd2448,32'd2524,32'd1359,32'd-2469,32'd-7475,32'd5566,32'd1947,32'd5888,32'd5952,32'd1440,32'd4257,32'd-5864,32'd1078,32'd-1600,32'd-328,32'd868,32'd3723,32'd-338,32'd-384,32'd941,32'd-2307,32'd207,32'd1534,32'd-1705,32'd-246,32'd-8657,32'd6044,32'd1732,32'd7944,32'd4594,32'd1986,32'd2119,32'd4248,32'd-579,32'd4465,32'd-263,32'd3967,32'd-3237,32'd4790,32'd-8359,32'd7626,32'd2429,32'd-1870,32'd621,32'd-266,32'd-2301,32'd5576,32'd-465,32'd3847,32'd3195,32'd-1972,32'd-1308,32'd2976,32'd7163,32'd3759,32'd4677,32'd3100,32'd-3078,32'd-5053,32'd-3364,32'd2905,32'd-6416,32'd1561,32'd2807,32'd1065,32'd753,32'd2301,32'd1939,32'd1721,32'd7446,32'd717,32'd-1356,32'd459,32'd-1361,32'd-120,32'd2978,32'd2106,32'd7612,32'd-1990,32'd-2071,32'd-3889,32'd858,32'd3911,32'd655,32'd-5942,32'd80,32'd5766,32'd-1872,32'd-2309,32'd-525,32'd1308,32'd-407,32'd4274,32'd-538,32'd1502,32'd10937,32'd-1864,32'd-6093,32'd-1645,32'd607,32'd12158,32'd-877,32'd2165,32'd2780,32'd-3659,32'd3249,32'd3852,32'd5112,32'd-4060,32'd-817,32'd9667,32'd-8540,32'd-2988,32'd-3627,32'd1110,32'd3613,32'd-6796,32'd7602,32'd5629,32'd6000,32'd570,32'd787,32'd2001,32'd5083,32'd-4846,32'd18085,32'd-693,32'd-1457,32'd3974,32'd-6948,32'd1937,32'd2604,32'd-214,32'd9399,32'd-9428,32'd-6240,32'd7504,32'd2355,32'd6757,32'd8041,32'd-13242,32'd4167,32'd-5263,32'd-2495,32'd-9497,32'd-9418,32'd4963,32'd-493,32'd-6376,32'd1906,32'd-1447,32'd4418,32'd14775,32'd6328,32'd1251,32'd4606,32'd14267,32'd3574,32'd1241,32'd3713,32'd-3178,32'd13125,32'd-905,32'd4028,32'd1607,32'd14990,32'd-2226,32'd3767,32'd-3913,32'd7998,32'd8916,32'd4619,32'd-9423,32'd-11650,32'd1064,32'd-7612,32'd8217,32'd-701,32'd1275,32'd-712,32'd4541,32'd1973,32'd3232,32'd5375,32'd9052,32'd-2839,32'd-2770,32'd514,32'd21269,32'd2683,32'd-3100,32'd-2237,32'd8930,32'd5122,32'd-2036,32'd5800,32'd1689,32'd-967,32'd-6547,32'd-1855,32'd327,32'd2337,32'd-1536,32'd-3789,32'd7368,32'd433,32'd-4804,32'd5024,32'd-2744,32'd-6201,32'd-2196,32'd-1416,32'd5092,32'd585,32'd2583,32'd-89,32'd-1348,32'd-4479,32'd550,32'd-1193,32'd-3989,32'd-1602,32'd-1539,32'd-4057,32'd-1329,32'd422,32'd-6503,32'd-863,32'd-11240,32'd4645,32'd-7280,32'd-2005,32'd-1279,32'd348,32'd-6474,32'd-2169,32'd-1083,32'd-2200,32'd-11357,32'd1306,32'd2019,32'd-2218,32'd-2257,32'd-6401,32'd629,32'd8208,32'd1861,32'd-946,32'd6411,32'd-6020,32'd4533,32'd-2218,32'd-1772,32'd-43,32'd-1405,32'd-3637,32'd-5498,32'd7592,32'd-2390,32'd3679,32'd-2719,32'd-5942,32'd-1932,32'd403,32'd3693,32'd-2985,32'd-2260,32'd9580,32'd520,32'd626,32'd-8427,32'd2912,32'd-4006,32'd-3032,32'd-655,32'd-5166,32'd725,32'd-2432,32'd-2204,32'd3784,32'd3642,32'd1762,32'd-2604,32'd-1309,32'd-3129,32'd-1157,32'd-2807,32'd-4162,32'd9892,32'd6210,32'd-7216,32'd-635,32'd-3325,32'd-2929,32'd-888,32'd7163,32'd9414,32'd-2041,32'd-3664,32'd5986,32'd-522,32'd1590,32'd1678,32'd-3837,32'd3251,32'd6074,32'd3728,32'd-1811,32'd529,32'd763,32'd1864,32'd4165,32'd-955,32'd90,32'd1394,32'd-671,32'd5000,32'd1203,32'd-8911,32'd2565,32'd-850,32'd97,32'd1197,32'd7583,32'd4682,32'd5292,32'd-1575,32'd-941,32'd3137,32'd2211,32'd3198,32'd-2150,32'd-7104,32'd-2149,32'd-3420,32'd-4731,32'd5053,32'd-8212,32'd-1993,32'd1730,32'd4821,32'd3066,32'd-7324,32'd2521,32'd2702,32'd4438,32'd7895,32'd8457,32'd1910,32'd3281,32'd4916,32'd-8232,32'd4516,32'd6708,32'd-9023,32'd1790,32'd5209,32'd-952,32'd2844,32'd-7802,32'd-1243,32'd-1411,32'd-3735,32'd5722,32'd3474,32'd-3916,32'd-8198,32'd10546,32'd-4560,32'd3688,32'd4680,32'd10273,32'd2182,32'd-2756,32'd-656,32'd1950,32'd4328,32'd60,32'd-14609,32'd5771,32'd-3959,32'd4157,32'd2687,32'd-6401,32'd1051,32'd2276,32'd1774,32'd-25976,32'd-7011,32'd3432,32'd-8798,32'd-14257,32'd534,32'd-1916};
    Wx[83]='{32'd-582,32'd-1033,32'd-401,32'd-1933,32'd2026,32'd-577,32'd-912,32'd-972,32'd223,32'd-3911,32'd-905,32'd-5029,32'd2587,32'd-1739,32'd1628,32'd6660,32'd3608,32'd-1771,32'd-1656,32'd347,32'd621,32'd-2966,32'd-1280,32'd-131,32'd2465,32'd-3894,32'd-2232,32'd-1411,32'd-1236,32'd2583,32'd1002,32'd1259,32'd-809,32'd-999,32'd-3876,32'd1892,32'd-3303,32'd-1593,32'd-786,32'd-3964,32'd-1370,32'd-55,32'd574,32'd-5595,32'd-1088,32'd-2471,32'd-4663,32'd-6445,32'd364,32'd-948,32'd-8164,32'd-2512,32'd-1979,32'd4440,32'd2719,32'd-1582,32'd3085,32'd-5478,32'd5122,32'd-6108,32'd861,32'd-3525,32'd-4113,32'd2934,32'd-301,32'd913,32'd-941,32'd-5898,32'd1672,32'd-219,32'd-2973,32'd-1334,32'd5781,32'd-301,32'd-1090,32'd-1550,32'd-4826,32'd-3613,32'd6899,32'd-3422,32'd-1053,32'd-120,32'd-759,32'd6000,32'd642,32'd509,32'd-234,32'd-785,32'd832,32'd-698,32'd1522,32'd-701,32'd-4401,32'd4128,32'd-5546,32'd1606,32'd2263,32'd3854,32'd1580,32'd2517,32'd5053,32'd-2651,32'd827,32'd933,32'd-1412,32'd-1651,32'd5327,32'd-1815,32'd-12812,32'd-209,32'd10634,32'd-981,32'd5473,32'd-9262,32'd-15214,32'd-4467,32'd-14873,32'd-4526,32'd-5034,32'd-4250,32'd-2863,32'd-7963,32'd-6035,32'd-6967,32'd2449,32'd-11777,32'd-2397,32'd3886,32'd3627,32'd-6840,32'd4108,32'd629,32'd-5942,32'd4670,32'd-4916,32'd-3479,32'd219,32'd-533,32'd-15253,32'd6494,32'd5761,32'd12558,32'd-5434,32'd-18310,32'd-14716,32'd2274,32'd-13798,32'd-4846,32'd1132,32'd896,32'd-6816,32'd1259,32'd-3129,32'd-5058,32'd9023,32'd-949,32'd8354,32'd1516,32'd-4382,32'd-6503,32'd887,32'd11992,32'd4243,32'd-9760,32'd-1523,32'd277,32'd-3364,32'd1087,32'd-1124,32'd4985,32'd7763,32'd4606,32'd803,32'd-9042,32'd451,32'd-3732,32'd-6464,32'd15927,32'd4838,32'd5493,32'd3425,32'd-13662,32'd-2303,32'd5966,32'd-3078,32'd-1063,32'd-505,32'd744,32'd173,32'd-233,32'd5766,32'd9970,32'd1649,32'd847,32'd2607,32'd4904,32'd2087,32'd-6826,32'd731,32'd-15039,32'd-2448,32'd-441,32'd-725,32'd-284,32'd-4636,32'd710,32'd2829,32'd-3583,32'd314,32'd-3549,32'd191,32'd-1904,32'd-5395,32'd-5463,32'd-8725,32'd3425,32'd3132,32'd-1496,32'd1596,32'd844,32'd-1851,32'd-3317,32'd-3176,32'd-2185,32'd-2556,32'd-1783,32'd-2519,32'd-5454,32'd5385,32'd-2181,32'd43,32'd1724,32'd9497,32'd-442,32'd-3723,32'd-3054,32'd1413,32'd3166,32'd-3024,32'd9497,32'd-3256,32'd12617,32'd-2482,32'd969,32'd-7558,32'd1682,32'd219,32'd11923,32'd-727,32'd1809,32'd2475,32'd-2259,32'd-2301,32'd497,32'd-2437,32'd4992,32'd5454,32'd-6040,32'd-4313,32'd1252,32'd1994,32'd277,32'd-3151,32'd8168,32'd-3452,32'd330,32'd3698,32'd11953,32'd2147,32'd-554,32'd1959,32'd4086,32'd2176,32'd3742,32'd-890,32'd2812,32'd6928,32'd4465,32'd5292,32'd-794,32'd2873,32'd9755,32'd-4296,32'd8769,32'd997,32'd-1842,32'd-1508,32'd54,32'd545,32'd2517,32'd-7890,32'd780,32'd262,32'd4880,32'd-1484,32'd7666,32'd-791,32'd896,32'd-6625,32'd-8730,32'd1109,32'd-6660,32'd-19511,32'd3811,32'd-3337,32'd-1440,32'd-1100,32'd1915,32'd-6298,32'd-3317,32'd-3957,32'd-3586,32'd7978,32'd-3596,32'd-5932,32'd-4638,32'd-3972,32'd-5522,32'd-3784,32'd-5712,32'd-825,32'd955,32'd-9287,32'd-3222,32'd4270,32'd-572,32'd-1655,32'd-2022,32'd8872,32'd-969,32'd-3254,32'd1726,32'd8417,32'd-2092,32'd9819,32'd334,32'd-4118,32'd4965,32'd-778,32'd10585,32'd-3710,32'd1079,32'd-679,32'd-5620,32'd1148,32'd-3586,32'd7309,32'd3889,32'd409,32'd-336,32'd-2836,32'd1608,32'd44,32'd509,32'd-8354,32'd-1884,32'd8110,32'd-10302,32'd-1156,32'd-3596,32'd-953,32'd-1264,32'd329,32'd-1979,32'd-2624,32'd-8193,32'd8349,32'd7080,32'd-1848,32'd186,32'd6542,32'd-1215,32'd-1683,32'd6660,32'd-6894,32'd1354,32'd3967,32'd44,32'd9365,32'd2392,32'd3210,32'd-5488,32'd-5781,32'd2614,32'd-603,32'd-181,32'd-1414,32'd-448,32'd3928,32'd1954,32'd-5346,32'd733,32'd-5400,32'd2797,32'd1901,32'd2137,32'd3906,32'd-9921,32'd3073,32'd-6938};
    Wx[84]='{32'd2491,32'd1916,32'd-1733,32'd-1373,32'd622,32'd-1369,32'd1494,32'd-1162,32'd1933,32'd-1331,32'd2215,32'd653,32'd33,32'd4189,32'd5297,32'd84,32'd2670,32'd732,32'd-223,32'd969,32'd-1589,32'd-3686,32'd-3789,32'd-1995,32'd3383,32'd-5151,32'd2027,32'd-765,32'd1516,32'd21,32'd-562,32'd-486,32'd3974,32'd2368,32'd802,32'd547,32'd-409,32'd-74,32'd1319,32'd-5957,32'd-662,32'd2810,32'd1601,32'd-3457,32'd265,32'd1568,32'd10830,32'd3442,32'd-1833,32'd-280,32'd-3757,32'd3745,32'd1379,32'd-319,32'd2597,32'd-3798,32'd-153,32'd3815,32'd1405,32'd-6098,32'd-1754,32'd164,32'd2271,32'd-1965,32'd2458,32'd-1821,32'd-2396,32'd-3100,32'd1580,32'd1094,32'd-149,32'd3388,32'd-2348,32'd-1689,32'd-2680,32'd-1674,32'd3112,32'd-125,32'd5688,32'd252,32'd1231,32'd6201,32'd1297,32'd-598,32'd4865,32'd2276,32'd-2354,32'd5659,32'd-4008,32'd-1041,32'd2731,32'd-2578,32'd5854,32'd-3586,32'd-5092,32'd3381,32'd2934,32'd761,32'd1115,32'd4841,32'd3657,32'd9013,32'd1309,32'd-3874,32'd-3613,32'd-269,32'd5122,32'd-6962,32'd-1163,32'd5195,32'd2280,32'd-3164,32'd2768,32'd5341,32'd423,32'd-19980,32'd5590,32'd-5937,32'd-4868,32'd500,32'd-465,32'd-3452,32'd-1844,32'd3811,32'd4768,32'd22,32'd-3745,32'd3364,32'd-5141,32'd-6655,32'd4433,32'd-1300,32'd3754,32'd-2817,32'd-6674,32'd6938,32'd2402,32'd-1134,32'd-4523,32'd-6171,32'd-5297,32'd5615,32'd-1408,32'd-2114,32'd-8417,32'd1429,32'd4104,32'd4826,32'd566,32'd3828,32'd9648,32'd-358,32'd1226,32'd14736,32'd4941,32'd8940,32'd8061,32'd1414,32'd-1296,32'd-3110,32'd-852,32'd-11171,32'd-8046,32'd-6381,32'd-7172,32'd3627,32'd-570,32'd21660,32'd-4106,32'd120,32'd9697,32'd-6840,32'd-98,32'd-7749,32'd-1441,32'd4916,32'd1369,32'd1229,32'd422,32'd-8378,32'd918,32'd-8417,32'd2022,32'd9169,32'd6733,32'd-443,32'd2548,32'd8657,32'd-5888,32'd3034,32'd-1658,32'd3493,32'd-2587,32'd4213,32'd-6464,32'd3647,32'd10136,32'd1182,32'd2707,32'd-17998,32'd-1466,32'd-11074,32'd-2229,32'd806,32'd-6313,32'd894,32'd-4931,32'd-1051,32'd-4672,32'd-4812,32'd612,32'd-21,32'd-5703,32'd-11904,32'd-209,32'd-1313,32'd-7548,32'd-1663,32'd3002,32'd1588,32'd1138,32'd-897,32'd908,32'd-9907,32'd-2924,32'd244,32'd1939,32'd-1052,32'd235,32'd-1235,32'd-6352,32'd-8354,32'd-5639,32'd-6645,32'd-4028,32'd-1066,32'd-4572,32'd-1049,32'd-1582,32'd3872,32'd-5502,32'd7832,32'd4213,32'd-2741,32'd-2082,32'd375,32'd-10361,32'd2919,32'd-1062,32'd-1773,32'd8989,32'd-1320,32'd-907,32'd-894,32'd-2093,32'd7500,32'd320,32'd881,32'd1707,32'd8588,32'd339,32'd-3828,32'd-6406,32'd-2983,32'd-3381,32'd2614,32'd274,32'd12597,32'd-911,32'd3366,32'd-6718,32'd458,32'd2614,32'd-3208,32'd-6523,32'd-1057,32'd5590,32'd-5322,32'd1682,32'd-1922,32'd-3266,32'd-7353,32'd-7119,32'd-3686,32'd-104,32'd-6962,32'd-578,32'd-1429,32'd4782,32'd2768,32'd-874,32'd-2634,32'd-3713,32'd-738,32'd477,32'd-330,32'd1296,32'd-5102,32'd-2834,32'd-9736,32'd-419,32'd-6318,32'd-5375,32'd-1555,32'd-6445,32'd-1383,32'd-3698,32'd31,32'd-1452,32'd-3439,32'd-2028,32'd5654,32'd-1156,32'd-1674,32'd3471,32'd1943,32'd1835,32'd2070,32'd-247,32'd-1728,32'd-1389,32'd-3527,32'd-6269,32'd-1844,32'd-2360,32'd12158,32'd-769,32'd-2639,32'd9809,32'd-6767,32'd92,32'd-1630,32'd-732,32'd-1389,32'd2060,32'd21,32'd-1495,32'd-802,32'd-1776,32'd-2442,32'd355,32'd8364,32'd2215,32'd-1640,32'd-11,32'd1992,32'd-4187,32'd-869,32'd-8417,32'd5825,32'd8339,32'd-2335,32'd-6333,32'd1566,32'd949,32'd51,32'd6777,32'd-4392,32'd-1998,32'd-8037,32'd-881,32'd1168,32'd-9428,32'd-6826,32'd-1990,32'd2104,32'd-5483,32'd1629,32'd6948,32'd-2846,32'd-417,32'd1700,32'd4394,32'd-2456,32'd-4667,32'd-1644,32'd121,32'd-5092,32'd6904,32'd814,32'd-2047,32'd-7045,32'd-4865,32'd-5229,32'd3823,32'd-1549,32'd-2944,32'd3403,32'd5776,32'd-2849,32'd8735,32'd-6259,32'd228,32'd1278,32'd5517,32'd-6079,32'd10751,32'd-7275,32'd-6020,32'd-3190};
    Wx[85]='{32'd1004,32'd131,32'd2238,32'd-1044,32'd1313,32'd289,32'd3151,32'd2631,32'd3447,32'd414,32'd4130,32'd436,32'd4050,32'd3879,32'd2055,32'd4602,32'd-154,32'd2700,32'd3266,32'd-281,32'd-673,32'd-625,32'd3596,32'd-3535,32'd826,32'd3437,32'd-663,32'd4475,32'd-162,32'd1242,32'd-464,32'd-370,32'd-4997,32'd-29,32'd7094,32'd1867,32'd5258,32'd2193,32'd-8496,32'd3178,32'd2366,32'd-1922,32'd1446,32'd-1623,32'd-535,32'd4291,32'd8041,32'd3127,32'd-392,32'd2807,32'd9648,32'd3410,32'd4616,32'd-4565,32'd515,32'd13339,32'd-212,32'd-729,32'd-281,32'd5688,32'd6484,32'd3281,32'd3247,32'd7343,32'd5366,32'd-1716,32'd-26,32'd9375,32'd1818,32'd1109,32'd5068,32'd1668,32'd2788,32'd1101,32'd2111,32'd5883,32'd1055,32'd1768,32'd1522,32'd7231,32'd1846,32'd3149,32'd-719,32'd-2115,32'd6396,32'd1162,32'd745,32'd3208,32'd3649,32'd2404,32'd4543,32'd-6542,32'd1079,32'd4995,32'd-4560,32'd5527,32'd9643,32'd-470,32'd-3286,32'd-858,32'd-1074,32'd-21875,32'd2286,32'd-3601,32'd-23,32'd1358,32'd-7485,32'd153,32'd1774,32'd2741,32'd9458,32'd2917,32'd-1988,32'd-3562,32'd-5517,32'd10429,32'd-2491,32'd-7402,32'd-1594,32'd1403,32'd-729,32'd-5327,32'd-8349,32'd3183,32'd-1326,32'd-3361,32'd574,32'd-3286,32'd-6030,32'd370,32'd-1420,32'd-9951,32'd4309,32'd-14521,32'd-52,32'd841,32'd-1861,32'd7504,32'd-7973,32'd-7739,32'd-7387,32'd7724,32'd2312,32'd5395,32'd-9833,32'd-18945,32'd-12509,32'd-166,32'd2286,32'd-1457,32'd-5786,32'd14951,32'd-3757,32'd8364,32'd-7983,32'd1556,32'd-5341,32'd4,32'd-11123,32'd4296,32'd-8120,32'd-204,32'd7592,32'd4399,32'd3991,32'd-792,32'd-77,32'd10273,32'd-2524,32'd4086,32'd-15410,32'd-461,32'd-59,32'd4975,32'd-1122,32'd-9458,32'd15781,32'd-3623,32'd6347,32'd11044,32'd-7412,32'd-15322,32'd-3632,32'd17304,32'd-445,32'd3737,32'd-5629,32'd2658,32'd-2047,32'd-3398,32'd8115,32'd5825,32'd7622,32'd-675,32'd10546,32'd6401,32'd-2573,32'd-6279,32'd-6923,32'd11103,32'd-494,32'd-703,32'd-319,32'd3515,32'd2600,32'd-420,32'd-4921,32'd8354,32'd5620,32'd3232,32'd6870,32'd4868,32'd-1406,32'd18437,32'd7319,32'd-98,32'd186,32'd3469,32'd1853,32'd3142,32'd1481,32'd6479,32'd-38,32'd-3476,32'd-2434,32'd1702,32'd4794,32'd2252,32'd9965,32'd-1175,32'd2995,32'd12021,32'd-4233,32'd-1672,32'd-5703,32'd794,32'd-4423,32'd1258,32'd2636,32'd3527,32'd941,32'd2435,32'd-3107,32'd-1550,32'd13789,32'd607,32'd-3149,32'd6313,32'd2719,32'd2983,32'd784,32'd1027,32'd759,32'd2276,32'd2408,32'd-4416,32'd-974,32'd-2966,32'd4504,32'd-4252,32'd-2015,32'd4345,32'd-4697,32'd2807,32'd1041,32'd-2041,32'd-4013,32'd-494,32'd1074,32'd417,32'd-438,32'd4328,32'd4731,32'd2309,32'd1018,32'd-1160,32'd-8315,32'd6250,32'd-5292,32'd6181,32'd1175,32'd2126,32'd8164,32'd-6113,32'd-933,32'd-2785,32'd2238,32'd5634,32'd-1815,32'd316,32'd-3430,32'd4282,32'd3740,32'd-4252,32'd7285,32'd-7177,32'd-1634,32'd11044,32'd3969,32'd1141,32'd-3781,32'd8706,32'd-549,32'd6459,32'd3884,32'd7895,32'd13300,32'd-5200,32'd2319,32'd1429,32'd15488,32'd8696,32'd-1247,32'd13837,32'd942,32'd-2795,32'd-2797,32'd12744,32'd1838,32'd-3081,32'd-7641,32'd9145,32'd629,32'd-3159,32'd-7407,32'd621,32'd-2154,32'd90,32'd-1905,32'd606,32'd996,32'd4821,32'd2812,32'd-2775,32'd-1730,32'd1378,32'd-4489,32'd-2006,32'd4833,32'd8720,32'd-3134,32'd7954,32'd2675,32'd4470,32'd4206,32'd-2194,32'd-4472,32'd5410,32'd9663,32'd3317,32'd-4516,32'd7788,32'd11884,32'd14414,32'd4094,32'd-4443,32'd4238,32'd-13691,32'd2100,32'd-7241,32'd-2335,32'd4450,32'd769,32'd3305,32'd-2008,32'd-13691,32'd-2949,32'd433,32'd10781,32'd946,32'd6630,32'd6748,32'd3305,32'd10058,32'd-129,32'd8251,32'd-3454,32'd8271,32'd-1965,32'd-1950,32'd-427,32'd10400,32'd9799,32'd-7758,32'd-12929,32'd3010,32'd3288,32'd9189,32'd-1560,32'd-9545,32'd2614,32'd2617,32'd9423,32'd-13574,32'd12275,32'd2420,32'd-6103,32'd-8735,32'd715,32'd9355};
    Wx[86]='{32'd-1188,32'd3090,32'd4682,32'd125,32'd-1761,32'd2448,32'd1728,32'd2418,32'd920,32'd3261,32'd-6420,32'd-1583,32'd-3864,32'd5483,32'd8383,32'd-1411,32'd7216,32'd-354,32'd-2083,32'd2319,32'd-488,32'd1821,32'd-128,32'd1960,32'd-195,32'd-3500,32'd-2377,32'd-824,32'd2878,32'd1857,32'd675,32'd5249,32'd4550,32'd3596,32'd-3217,32'd1510,32'd4780,32'd-1683,32'd1533,32'd5805,32'd-369,32'd48,32'd-3959,32'd3459,32'd-8334,32'd1635,32'd-3889,32'd-3276,32'd-4204,32'd-337,32'd-259,32'd665,32'd-1740,32'd-466,32'd-1734,32'd-6215,32'd-2731,32'd-2117,32'd-127,32'd-4958,32'd-3747,32'd475,32'd-2963,32'd1387,32'd-622,32'd-1949,32'd-966,32'd-459,32'd-3322,32'd-4111,32'd-1917,32'd-2731,32'd-3361,32'd3271,32'd-588,32'd4226,32'd1328,32'd-483,32'd175,32'd-3803,32'd512,32'd-249,32'd3156,32'd4760,32'd-4162,32'd-3090,32'd-3398,32'd120,32'd238,32'd-213,32'd-134,32'd2391,32'd1972,32'd-3354,32'd10478,32'd-4326,32'd-1048,32'd-814,32'd-1267,32'd-4108,32'd3476,32'd-1425,32'd-4428,32'd-1604,32'd-2785,32'd-3461,32'd-4633,32'd-10029,32'd-4426,32'd-6528,32'd6069,32'd1162,32'd6166,32'd1904,32'd-21757,32'd3952,32'd-4670,32'd-4345,32'd-860,32'd-1293,32'd3911,32'd294,32'd717,32'd-223,32'd1755,32'd-1706,32'd-641,32'd-6640,32'd-5874,32'd1501,32'd-5703,32'd2274,32'd-1474,32'd623,32'd-1502,32'd-5751,32'd2724,32'd1713,32'd-3479,32'd3481,32'd1612,32'd-11708,32'd-4973,32'd2430,32'd-8110,32'd-2291,32'd-679,32'd-843,32'd259,32'd-635,32'd-862,32'd5375,32'd-472,32'd-5639,32'd-8852,32'd3132,32'd-3371,32'd1373,32'd-8432,32'd2062,32'd-518,32'd171,32'd-1379,32'd2519,32'd-17128,32'd1505,32'd3024,32'd3120,32'd1771,32'd-1845,32'd-3637,32'd10429,32'd1734,32'd8437,32'd1060,32'd-6259,32'd10546,32'd-2517,32'd1893,32'd2551,32'd-9306,32'd19003,32'd1566,32'd-2232,32'd-2805,32'd10117,32'd-4416,32'd4111,32'd477,32'd-58,32'd-5610,32'd2687,32'd10292,32'd-5444,32'd-1655,32'd-485,32'd1477,32'd-15302,32'd-9174,32'd299,32'd-4074,32'd3740,32'd1192,32'd2883,32'd3383,32'd527,32'd-5156,32'd-8896,32'd-508,32'd-362,32'd3659,32'd-35,32'd-442,32'd1155,32'd-6367,32'd-3767,32'd-6166,32'd3601,32'd-1746,32'd-4770,32'd1165,32'd-1745,32'd-3715,32'd2386,32'd2409,32'd968,32'd19,32'd-3125,32'd-2902,32'd-49,32'd4135,32'd3427,32'd1431,32'd-491,32'd-1370,32'd3813,32'd-2963,32'd634,32'd7192,32'd-3527,32'd-463,32'd-9536,32'd-1352,32'd-3881,32'd-4111,32'd1860,32'd-4331,32'd4235,32'd4348,32'd4130,32'd-184,32'd1362,32'd-154,32'd-1695,32'd-2054,32'd4086,32'd4282,32'd-5249,32'd214,32'd2888,32'd-1492,32'd-1062,32'd-218,32'd667,32'd3859,32'd127,32'd-3820,32'd5576,32'd-1619,32'd-4206,32'd1236,32'd5312,32'd-2481,32'd6743,32'd-1881,32'd-6621,32'd-11748,32'd-610,32'd-2019,32'd2352,32'd-273,32'd-4682,32'd-1341,32'd9912,32'd3247,32'd-8642,32'd-4,32'd-203,32'd-1782,32'd433,32'd9189,32'd7192,32'd-3713,32'd-811,32'd2626,32'd-831,32'd-1856,32'd-945,32'd-7871,32'd7182,32'd2990,32'd-929,32'd1190,32'd5019,32'd5214,32'd-3081,32'd-2268,32'd3300,32'd2717,32'd5698,32'd-637,32'd-4606,32'd-715,32'd-156,32'd-7402,32'd5415,32'd2565,32'd-3610,32'd4570,32'd-4638,32'd9638,32'd5234,32'd2048,32'd3852,32'd5449,32'd737,32'd-2209,32'd-3315,32'd-10283,32'd889,32'd281,32'd2393,32'd-707,32'd2875,32'd1436,32'd3659,32'd1359,32'd-813,32'd2797,32'd155,32'd-1674,32'd-5878,32'd2209,32'd1904,32'd-3491,32'd2459,32'd2658,32'd3986,32'd4846,32'd-1882,32'd-442,32'd3737,32'd4311,32'd-7944,32'd-3420,32'd4172,32'd1071,32'd-2995,32'd1158,32'd4321,32'd-2517,32'd-2327,32'd7631,32'd-772,32'd-1582,32'd-4475,32'd-12197,32'd1539,32'd-3432,32'd494,32'd-2463,32'd-480,32'd-10458,32'd-3559,32'd545,32'd-1002,32'd-7514,32'd-364,32'd-4975,32'd-4179,32'd4711,32'd773,32'd770,32'd8437,32'd848,32'd1018,32'd230,32'd2393,32'd356,32'd-5131,32'd867,32'd1032,32'd-2568,32'd-15761,32'd10556,32'd-1633,32'd879,32'd-3815,32'd-5766,32'd4960};
    Wx[87]='{32'd3398,32'd1440,32'd1127,32'd-91,32'd650,32'd-1536,32'd-7763,32'd-612,32'd-370,32'd-82,32'd2163,32'd887,32'd4372,32'd-2412,32'd882,32'd6162,32'd-5322,32'd-4355,32'd1099,32'd2712,32'd1966,32'd-3210,32'd-4140,32'd4291,32'd-3220,32'd3669,32'd-568,32'd3793,32'd-2468,32'd-3840,32'd772,32'd-2377,32'd3083,32'd1,32'd7280,32'd1588,32'd243,32'd2810,32'd3959,32'd-2917,32'd-1202,32'd2670,32'd316,32'd3808,32'd3176,32'd-4291,32'd2409,32'd1634,32'd4650,32'd4023,32'd-2398,32'd-531,32'd-3981,32'd3305,32'd420,32'd-2819,32'd-1689,32'd3483,32'd-572,32'd-5361,32'd1206,32'd1572,32'd-1267,32'd-850,32'd851,32'd-1303,32'd-285,32'd11406,32'd3344,32'd-2744,32'd1395,32'd-315,32'd2734,32'd-258,32'd895,32'd-2037,32'd-1992,32'd-4555,32'd3703,32'd358,32'd-2459,32'd3066,32'd1357,32'd5981,32'd-3461,32'd-1984,32'd-747,32'd-1108,32'd-1300,32'd-175,32'd-4702,32'd3991,32'd-1181,32'd170,32'd1295,32'd4926,32'd-3527,32'd496,32'd-897,32'd102,32'd1427,32'd-19052,32'd-153,32'd2453,32'd3068,32'd-249,32'd24687,32'd6508,32'd289,32'd4460,32'd15791,32'd385,32'd1861,32'd-11484,32'd12021,32'd-1557,32'd-6708,32'd-1206,32'd3344,32'd3,32'd-510,32'd2653,32'd3745,32'd5092,32'd2944,32'd-4177,32'd-797,32'd-5434,32'd-6528,32'd-2452,32'd405,32'd1278,32'd-13476,32'd4948,32'd4707,32'd-3964,32'd7553,32'd1462,32'd1441,32'd9643,32'd-1562,32'd-10830,32'd-1588,32'd-4235,32'd115,32'd11884,32'd-7998,32'd-101,32'd-5854,32'd-2585,32'd19599,32'd-867,32'd-9106,32'd4477,32'd9902,32'd1662,32'd-2905,32'd-5346,32'd10175,32'd1671,32'd-5205,32'd6308,32'd-2768,32'd3095,32'd13994,32'd839,32'd312,32'd-8193,32'd-1651,32'd-361,32'd-108,32'd-683,32'd2976,32'd1402,32'd-4338,32'd2680,32'd1887,32'd3972,32'd9697,32'd1956,32'd-10761,32'd-9326,32'd685,32'd-7197,32'd-1491,32'd9130,32'd-687,32'd1380,32'd7475,32'd-2481,32'd12285,32'd-10087,32'd2456,32'd3305,32'd2358,32'd3955,32'd-8437,32'd-8789,32'd-2066,32'd-2517,32'd3740,32'd-972,32'd1181,32'd3190,32'd850,32'd-855,32'd4641,32'd-3867,32'd1966,32'd-2854,32'd-5639,32'd56,32'd-231,32'd-2095,32'd5151,32'd3315,32'd11503,32'd5048,32'd-1643,32'd3613,32'd2731,32'd-2093,32'd-3029,32'd2044,32'd-2230,32'd-3669,32'd-2902,32'd2406,32'd4343,32'd3464,32'd3437,32'd593,32'd9516,32'd-4860,32'd-414,32'd2136,32'd3234,32'd-1535,32'd1329,32'd-873,32'd5043,32'd-646,32'd-10292,32'd-1678,32'd-408,32'd4558,32'd-6289,32'd-1213,32'd-1259,32'd1529,32'd-9213,32'd1704,32'd-1601,32'd539,32'd551,32'd-7578,32'd-1423,32'd614,32'd5332,32'd-632,32'd-3059,32'd556,32'd-6645,32'd4624,32'd-1157,32'd-2839,32'd1791,32'd-6772,32'd4948,32'd-3796,32'd-9057,32'd-3447,32'd1682,32'd2670,32'd338,32'd9135,32'd8237,32'd2844,32'd-4997,32'd6132,32'd1809,32'd-3518,32'd1409,32'd-650,32'd-1485,32'd1222,32'd107,32'd-1645,32'd60,32'd-2646,32'd7387,32'd-939,32'd5756,32'd-1632,32'd3261,32'd3022,32'd7543,32'd-6728,32'd-4272,32'd-3251,32'd3623,32'd-60,32'd5292,32'd-670,32'd2471,32'd4035,32'd5078,32'd-8012,32'd2043,32'd5771,32'd-2565,32'd-4284,32'd12158,32'd-8486,32'd-1383,32'd-3818,32'd-494,32'd-3234,32'd-4638,32'd7187,32'd1849,32'd-1998,32'd-1453,32'd293,32'd1137,32'd-535,32'd-8745,32'd-1150,32'd7329,32'd8056,32'd2551,32'd3649,32'd2817,32'd-5810,32'd-8085,32'd4274,32'd-7656,32'd1696,32'd3022,32'd343,32'd2563,32'd-7153,32'd1849,32'd1150,32'd-4182,32'd-7583,32'd174,32'd-2985,32'd2303,32'd932,32'd7138,32'd-4208,32'd-3813,32'd4709,32'd-11230,32'd-6440,32'd-1719,32'd9414,32'd6977,32'd-7294,32'd3308,32'd955,32'd11240,32'd-3054,32'd-8085,32'd345,32'd-7250,32'd-3752,32'd9477,32'd-1518,32'd2873,32'd-4641,32'd1456,32'd1606,32'd-4245,32'd3518,32'd3906,32'd16,32'd-661,32'd791,32'd-2709,32'd-13593,32'd2083,32'd8754,32'd-4028,32'd239,32'd-5917,32'd-438,32'd3876,32'd12441,32'd-647,32'd-1853,32'd-5024,32'd579,32'd8950,32'd6875,32'd-2680,32'd-4880,32'd791,32'd1501};
    Wx[88]='{32'd2800,32'd-3378,32'd65,32'd-1748,32'd-2604,32'd1669,32'd1877,32'd1329,32'd-856,32'd115,32'd-3159,32'd1519,32'd-1369,32'd-5419,32'd-1586,32'd-6533,32'd2634,32'd-1289,32'd1287,32'd678,32'd-969,32'd-739,32'd3217,32'd1794,32'd-5073,32'd281,32'd-80,32'd-2834,32'd2749,32'd-3383,32'd-901,32'd-8291,32'd6416,32'd1397,32'd-3381,32'd-5019,32'd193,32'd3400,32'd-593,32'd3059,32'd561,32'd-161,32'd-2036,32'd-11708,32'd-3100,32'd1947,32'd2819,32'd-3952,32'd-1093,32'd1956,32'd-1568,32'd4628,32'd333,32'd-654,32'd-2858,32'd-1564,32'd-3610,32'd-492,32'd-723,32'd2565,32'd726,32'd-2421,32'd2073,32'd-1668,32'd-2954,32'd4558,32'd-4162,32'd-7124,32'd-1040,32'd1212,32'd-2243,32'd-5170,32'd1667,32'd-5976,32'd736,32'd2292,32'd-4487,32'd-3505,32'd-963,32'd-1649,32'd-808,32'd4089,32'd-3173,32'd2680,32'd-1660,32'd2003,32'd-1275,32'd-1220,32'd1676,32'd544,32'd-5908,32'd-4099,32'd3679,32'd1982,32'd1793,32'd1130,32'd-6914,32'd6679,32'd1854,32'd-4138,32'd-1292,32'd-7451,32'd-30,32'd-2907,32'd2785,32'd-27,32'd-2067,32'd-11025,32'd4033,32'd6132,32'd-905,32'd-1552,32'd2124,32'd1707,32'd-6699,32'd2817,32'd-9248,32'd189,32'd3937,32'd1781,32'd3940,32'd4204,32'd-2521,32'd3496,32'd654,32'd-1026,32'd2626,32'd-2338,32'd-7285,32'd6411,32'd-9296,32'd-7495,32'd-2524,32'd670,32'd-2624,32'd-4431,32'd-2790,32'd-1744,32'd3146,32'd20546,32'd-12480,32'd-1154,32'd-1853,32'd1324,32'd-10185,32'd8403,32'd-12089,32'd4555,32'd2352,32'd-7939,32'd-611,32'd8496,32'd-1677,32'd1420,32'd-2377,32'd1385,32'd2312,32'd379,32'd2458,32'd-1604,32'd1916,32'd-7290,32'd803,32'd-2927,32'd-2133,32'd170,32'd-1512,32'd2666,32'd2790,32'd-2919,32'd1798,32'd-6450,32'd3413,32'd8100,32'd-119,32'd-8486,32'd-1196,32'd-8007,32'd8300,32'd411,32'd4816,32'd-7016,32'd-2471,32'd-1267,32'd-1485,32'd-1484,32'd1450,32'd655,32'd3366,32'd5541,32'd-1159,32'd-4587,32'd-4267,32'd-2475,32'd-5000,32'd8320,32'd-12314,32'd4296,32'd2441,32'd-9082,32'd378,32'd-3581,32'd-3476,32'd1102,32'd35,32'd-566,32'd2719,32'd-5375,32'd1464,32'd895,32'd-1575,32'd-3581,32'd-431,32'd-610,32'd5527,32'd8911,32'd-4357,32'd-3361,32'd-4555,32'd1051,32'd-569,32'd1229,32'd-3872,32'd-2148,32'd-274,32'd3486,32'd-1236,32'd2770,32'd-1945,32'd-2177,32'd-2988,32'd1330,32'd-12724,32'd4770,32'd5390,32'd4760,32'd-4423,32'd-645,32'd3930,32'd-1456,32'd5458,32'd3005,32'd10058,32'd6494,32'd11875,32'd-5400,32'd-5473,32'd-358,32'd-4008,32'd5288,32'd-6074,32'd-3508,32'd-4406,32'd-7036,32'd-431,32'd-216,32'd-2016,32'd597,32'd579,32'd-2371,32'd6948,32'd-1845,32'd1072,32'd707,32'd4357,32'd-2275,32'd-373,32'd-10927,32'd1530,32'd-2352,32'd-10029,32'd6401,32'd5395,32'd206,32'd-860,32'd1243,32'd8393,32'd1983,32'd3916,32'd-4338,32'd795,32'd-1727,32'd-1044,32'd167,32'd3435,32'd-29,32'd938,32'd-7978,32'd3701,32'd4343,32'd6323,32'd-689,32'd1204,32'd2644,32'd18925,32'd5429,32'd-5468,32'd4482,32'd-2563,32'd1915,32'd-3154,32'd-1085,32'd-15400,32'd-1735,32'd1455,32'd-13886,32'd708,32'd-4562,32'd205,32'd4116,32'd-3286,32'd-1368,32'd1768,32'd-7700,32'd-3222,32'd2539,32'd3581,32'd3542,32'd2160,32'd2792,32'd-5786,32'd1314,32'd1381,32'd-734,32'd995,32'd4558,32'd-4,32'd-434,32'd-1719,32'd-283,32'd-1839,32'd37,32'd-7036,32'd-1158,32'd4147,32'd-720,32'd-245,32'd6811,32'd-1429,32'd-5952,32'd5395,32'd-1172,32'd-571,32'd1324,32'd-156,32'd-4663,32'd-6474,32'd230,32'd-6704,32'd737,32'd-2362,32'd-7944,32'd-11005,32'd-1168,32'd4521,32'd2595,32'd3457,32'd-4555,32'd195,32'd11962,32'd-3762,32'd5107,32'd2160,32'd262,32'd-4411,32'd-8271,32'd0,32'd-10361,32'd-2995,32'd-1353,32'd-3315,32'd-2692,32'd1766,32'd-5014,32'd4167,32'd3972,32'd3159,32'd-1334,32'd-4284,32'd-6992,32'd2592,32'd791,32'd1511,32'd-3176,32'd-9082,32'd1202,32'd-3403,32'd-9516,32'd-2425,32'd-4645,32'd3122,32'd-1207,32'd2229,32'd6875,32'd9799,32'd2709,32'd-4868,32'd2824,32'd1760,32'd-3374};
    Wx[89]='{32'd2014,32'd-2607,32'd-1076,32'd5043,32'd1578,32'd1616,32'd-1625,32'd-6420,32'd2028,32'd1015,32'd177,32'd-2464,32'd112,32'd5214,32'd-717,32'd-4140,32'd364,32'd-3198,32'd581,32'd-845,32'd3823,32'd-2321,32'd-1276,32'd-1093,32'd-916,32'd2069,32'd-1529,32'd476,32'd5976,32'd-5913,32'd2778,32'd-3557,32'd-1324,32'd159,32'd-5756,32'd-2070,32'd2839,32'd-3925,32'd-4719,32'd3134,32'd-2410,32'd-2374,32'd971,32'd-3547,32'd6459,32'd-1722,32'd3339,32'd-5283,32'd2244,32'd1359,32'd-4191,32'd-3530,32'd4746,32'd-1666,32'd-1564,32'd-3520,32'd464,32'd-2015,32'd-2827,32'd-2902,32'd2348,32'd1119,32'd-4873,32'd1331,32'd-274,32'd-839,32'd-313,32'd4926,32'd4050,32'd66,32'd362,32'd1291,32'd65,32'd339,32'd-2927,32'd-1619,32'd-552,32'd-3413,32'd3388,32'd-3696,32'd-1151,32'd-2320,32'd345,32'd-4782,32'd-4255,32'd-811,32'd3146,32'd-1456,32'd-2761,32'd-1998,32'd-355,32'd-2460,32'd442,32'd1182,32'd-1799,32'd3535,32'd-2941,32'd3256,32'd-215,32'd-5654,32'd-7221,32'd-12666,32'd1137,32'd4462,32'd-995,32'd-635,32'd-14121,32'd13408,32'd-2047,32'd2856,32'd-7006,32'd-10146,32'd7465,32'd-2432,32'd-444,32'd834,32'd1546,32'd-4501,32'd1234,32'd-332,32'd850,32'd-6679,32'd-3596,32'd97,32'd-1668,32'd-746,32'd-765,32'd587,32'd-2138,32'd-6264,32'd-1334,32'd-2441,32'd-9711,32'd-9072,32'd-7265,32'd4038,32'd-3747,32'd-41,32'd8559,32'd167,32'd-927,32'd-15371,32'd2922,32'd-7167,32'd15625,32'd-16416,32'd-8608,32'd-666,32'd-4355,32'd14,32'd18994,32'd6508,32'd-2196,32'd-7124,32'd2902,32'd5336,32'd-728,32'd1301,32'd8032,32'd-2949,32'd-498,32'd13554,32'd-14794,32'd12138,32'd1104,32'd-2185,32'd1422,32'd-1566,32'd-1042,32'd-4,32'd1905,32'd-6381,32'd1704,32'd-2277,32'd-289,32'd-688,32'd-14443,32'd9028,32'd-7666,32'd-8862,32'd-10937,32'd3452,32'd5849,32'd-1503,32'd-7651,32'd-3378,32'd82,32'd-1763,32'd6372,32'd-4645,32'd-6738,32'd10888,32'd1406,32'd4111,32'd3862,32'd-817,32'd-3212,32'd3537,32'd9218,32'd-6640,32'd831,32'd3127,32'd-4462,32'd2526,32'd3090,32'd2988,32'd8251,32'd-3867,32'd-7753,32'd1743,32'd-2504,32'd5166,32'd467,32'd-4782,32'd-2573,32'd7348,32'd6235,32'd-2413,32'd1782,32'd-1998,32'd2274,32'd1282,32'd-443,32'd2452,32'd-1307,32'd4450,32'd916,32'd2851,32'd-2580,32'd4436,32'd1667,32'd2839,32'd-8803,32'd-4465,32'd-1333,32'd-5957,32'd2551,32'd-2178,32'd245,32'd-2915,32'd-2636,32'd4416,32'd941,32'd-1628,32'd-516,32'd1669,32'd-5302,32'd-8041,32'd2673,32'd-1002,32'd112,32'd2883,32'd1227,32'd-3024,32'd4042,32'd-197,32'd-2191,32'd-1505,32'd626,32'd1658,32'd-5825,32'd-13437,32'd-4023,32'd775,32'd7343,32'd-4865,32'd-307,32'd-3400,32'd2463,32'd1409,32'd-4628,32'd-2558,32'd227,32'd-2770,32'd-1967,32'd-1857,32'd9033,32'd-6665,32'd-6923,32'd1400,32'd-5058,32'd3437,32'd4497,32'd-2073,32'd1400,32'd187,32'd946,32'd-5991,32'd4135,32'd-2436,32'd-466,32'd7734,32'd-2270,32'd-3686,32'd-18886,32'd-7568,32'd-220,32'd-2260,32'd-4025,32'd-5952,32'd-957,32'd7568,32'd-1067,32'd-810,32'd-1452,32'd1898,32'd5034,32'd-6718,32'd-4672,32'd-2393,32'd4863,32'd4267,32'd42,32'd-429,32'd-8417,32'd-762,32'd5747,32'd3186,32'd-1837,32'd2873,32'd-8002,32'd564,32'd2489,32'd762,32'd-4116,32'd3642,32'd-2470,32'd-1374,32'd-7485,32'd-96,32'd-699,32'd1033,32'd-14130,32'd-5864,32'd1278,32'd-4204,32'd-3024,32'd-7539,32'd-7636,32'd-2775,32'd-1477,32'd-4731,32'd-1343,32'd-233,32'd673,32'd-4528,32'd-16630,32'd-3710,32'd-2084,32'd4230,32'd-4301,32'd-5649,32'd-3105,32'd1232,32'd-321,32'd-5551,32'd-3999,32'd5742,32'd1076,32'd-3444,32'd1120,32'd-2832,32'd-5087,32'd-5810,32'd-4250,32'd-722,32'd-3071,32'd-2182,32'd6054,32'd1395,32'd-212,32'd6215,32'd1189,32'd-5634,32'd-4855,32'd2988,32'd-4882,32'd-4284,32'd366,32'd-1051,32'd-5922,32'd204,32'd458,32'd-4941,32'd-45,32'd-5322,32'd2739,32'd-6152,32'd-3122,32'd319,32'd-3095,32'd7812,32'd-2941,32'd-1096,32'd-8481,32'd-302,32'd1861,32'd-1795,32'd-984,32'd-7988};
    Wx[90]='{32'd-272,32'd-3051,32'd18,32'd-451,32'd-2687,32'd-2575,32'd1196,32'd2626,32'd3366,32'd3132,32'd-1827,32'd603,32'd2492,32'd3571,32'd3669,32'd4409,32'd-8549,32'd863,32'd2548,32'd-672,32'd-2432,32'd1213,32'd-1126,32'd-34,32'd-594,32'd2578,32'd2846,32'd1715,32'd6479,32'd-2536,32'd-2368,32'd-6762,32'd-5366,32'd-1614,32'd2619,32'd-1053,32'd577,32'd1582,32'd-3503,32'd-2469,32'd-112,32'd-5117,32'd5039,32'd-5122,32'd8300,32'd661,32'd-60,32'd4653,32'd2099,32'd-1030,32'd5288,32'd-884,32'd-2973,32'd3793,32'd439,32'd-1871,32'd-2248,32'd-1427,32'd-5312,32'd2534,32'd-500,32'd2507,32'd-834,32'd-247,32'd-3596,32'd-3491,32'd1387,32'd-10615,32'd556,32'd-1060,32'd158,32'd-2448,32'd2529,32'd1531,32'd778,32'd-4272,32'd3569,32'd2388,32'd-1940,32'd-1824,32'd-808,32'd-6401,32'd-115,32'd-1411,32'd-5429,32'd-158,32'd-1058,32'd514,32'd2430,32'd-3989,32'd-5498,32'd-4108,32'd2246,32'd-629,32'd-1770,32'd3666,32'd1501,32'd-710,32'd-2012,32'd-1943,32'd226,32'd3041,32'd1738,32'd6513,32'd5805,32'd-1080,32'd11835,32'd1760,32'd-1639,32'd1361,32'd-4233,32'd-2910,32'd-3005,32'd-5073,32'd-6147,32'd16787,32'd5502,32'd12910,32'd3193,32'd383,32'd-711,32'd-3459,32'd6669,32'd-2792,32'd1824,32'd3896,32'd-1507,32'd-2509,32'd-9599,32'd5991,32'd-3322,32'd15136,32'd5087,32'd4157,32'd1640,32'd-1152,32'd3999,32'd13193,32'd14033,32'd-5576,32'd745,32'd-8120,32'd2016,32'd25664,32'd14199,32'd-14609,32'd11132,32'd-3647,32'd-3972,32'd-3049,32'd12871,32'd12021,32'd-2093,32'd35,32'd-1417,32'd-2049,32'd-1845,32'd935,32'd-12890,32'd5249,32'd1690,32'd4980,32'd19853,32'd-1062,32'd-12802,32'd-565,32'd-5668,32'd608,32'd-870,32'd-1785,32'd321,32'd5175,32'd-126,32'd-3427,32'd5195,32'd-2604,32'd-7709,32'd3068,32'd-321,32'd3916,32'd1660,32'd-2807,32'd2929,32'd270,32'd-3400,32'd-10634,32'd6621,32'd-76,32'd-2349,32'd-4689,32'd3298,32'd329,32'd569,32'd832,32'd6816,32'd3120,32'd-6884,32'd2492,32'd160,32'd-11142,32'd62,32'd8110,32'd501,32'd-682,32'd-797,32'd459,32'd-3530,32'd-7065,32'd3522,32'd1129,32'd-4042,32'd-900,32'd275,32'd-3312,32'd-3737,32'd1890,32'd684,32'd-3955,32'd3222,32'd-3696,32'd103,32'd-2016,32'd-376,32'd-1569,32'd828,32'd431,32'd-4655,32'd2834,32'd-9433,32'd290,32'd663,32'd153,32'd986,32'd1619,32'd-4899,32'd6777,32'd-1302,32'd1190,32'd-6425,32'd2636,32'd-2348,32'd-7104,32'd343,32'd-680,32'd-2687,32'd643,32'd8222,32'd-7597,32'd-2568,32'd-1384,32'd1527,32'd-3566,32'd1625,32'd401,32'd-446,32'd-1071,32'd8925,32'd3601,32'd2435,32'd503,32'd-2924,32'd-698,32'd-4079,32'd6904,32'd-5747,32'd-2980,32'd-1244,32'd-685,32'd-455,32'd-870,32'd258,32'd-1888,32'd3857,32'd4990,32'd2634,32'd-1334,32'd930,32'd-5874,32'd-4670,32'd7797,32'd-1933,32'd4958,32'd-2388,32'd-3466,32'd-6142,32'd1398,32'd1301,32'd3425,32'd1186,32'd-3044,32'd-1429,32'd-2631,32'd-360,32'd1001,32'd6499,32'd1260,32'd-5595,32'd3383,32'd2609,32'd-4645,32'd273,32'd3383,32'd3618,32'd668,32'd-840,32'd2690,32'd-3925,32'd-1251,32'd3088,32'd9819,32'd-5561,32'd1614,32'd8217,32'd2915,32'd-3344,32'd2756,32'd-2398,32'd4694,32'd2404,32'd958,32'd-219,32'd-961,32'd-1876,32'd-2092,32'd-2292,32'd-5908,32'd-5439,32'd4812,32'd1647,32'd-1480,32'd-5449,32'd2880,32'd-5229,32'd924,32'd5053,32'd-514,32'd-1037,32'd4020,32'd-1988,32'd-5854,32'd632,32'd-7885,32'd-236,32'd6625,32'd6645,32'd490,32'd6914,32'd-4455,32'd6025,32'd-1013,32'd573,32'd-1513,32'd5820,32'd-4724,32'd-1528,32'd-5576,32'd-1072,32'd6791,32'd3659,32'd7421,32'd1701,32'd4770,32'd-1759,32'd-416,32'd-1416,32'd-8120,32'd5195,32'd-8359,32'd10253,32'd3317,32'd1287,32'd-3586,32'd5229,32'd3425,32'd8295,32'd-1097,32'd-8027,32'd4584,32'd-4519,32'd2602,32'd3879,32'd2342,32'd260,32'd1695,32'd-11259,32'd5102,32'd-2890,32'd9072,32'd-2290,32'd4221,32'd1336,32'd2976,32'd-145,32'd-1121,32'd-965,32'd3244,32'd-8984,32'd-2156,32'd-223,32'd5390};
    Wx[91]='{32'd-883,32'd-6015,32'd-10468,32'd3513,32'd36,32'd1048,32'd1828,32'd-10185,32'd-2139,32'd1887,32'd4829,32'd4978,32'd4924,32'd-1612,32'd5800,32'd-3664,32'd2128,32'd4609,32'd3520,32'd3984,32'd714,32'd209,32'd-7421,32'd518,32'd2010,32'd1721,32'd1389,32'd1478,32'd5556,32'd1357,32'd1839,32'd1976,32'd7612,32'd-279,32'd-2398,32'd926,32'd-2788,32'd603,32'd-478,32'd3942,32'd26,32'd-1051,32'd-5185,32'd853,32'd3249,32'd914,32'd-1973,32'd1705,32'd5107,32'd-139,32'd1082,32'd-655,32'd266,32'd-200,32'd-5825,32'd-3325,32'd-2868,32'd1745,32'd1063,32'd-2663,32'd2291,32'd4191,32'd-2291,32'd-728,32'd-1870,32'd-957,32'd1168,32'd-3015,32'd-1448,32'd650,32'd405,32'd5346,32'd129,32'd3032,32'd-1081,32'd233,32'd10390,32'd899,32'd165,32'd574,32'd3767,32'd-2822,32'd-3361,32'd-2954,32'd3134,32'd10566,32'd1959,32'd-94,32'd2359,32'd-1782,32'd2604,32'd-3310,32'd5034,32'd-1343,32'd-2397,32'd4038,32'd-1796,32'd3708,32'd-902,32'd2849,32'd-1628,32'd7641,32'd3613,32'd311,32'd-282,32'd-1147,32'd6484,32'd12207,32'd4614,32'd-5214,32'd-498,32'd-2322,32'd4189,32'd-776,32'd-11640,32'd-20000,32'd2890,32'd2597,32'd3139,32'd2731,32'd-5073,32'd-3015,32'd10380,32'd-3786,32'd-690,32'd720,32'd6079,32'd-2934,32'd-463,32'd10439,32'd-2453,32'd884,32'd-365,32'd-2661,32'd-1522,32'd4309,32'd2423,32'd2687,32'd2489,32'd-9726,32'd4626,32'd-6611,32'd-5234,32'd9545,32'd-12021,32'd1944,32'd18906,32'd-2022,32'd6098,32'd-2326,32'd10322,32'd-11103,32'd1512,32'd-9213,32'd3405,32'd-794,32'd5600,32'd-510,32'd1856,32'd-3037,32'd699,32'd-13193,32'd3854,32'd-8251,32'd2636,32'd-2257,32'd-2254,32'd-11611,32'd-1358,32'd-2741,32'd-2441,32'd-4536,32'd-1290,32'd-2546,32'd-3342,32'd3923,32'd3161,32'd1666,32'd5776,32'd-2626,32'd-3217,32'd2954,32'd-8769,32'd-15781,32'd-732,32'd3571,32'd-2885,32'd-12480,32'd240,32'd-8271,32'd-343,32'd6791,32'd-5664,32'd1647,32'd5708,32'd2568,32'd3125,32'd5561,32'd-4401,32'd-1557,32'd6601,32'd-2104,32'd-5361,32'd134,32'd3911,32'd-179,32'd1007,32'd10605,32'd-2087,32'd-477,32'd-3618,32'd-2687,32'd6264,32'd-10947,32'd-1022,32'd2171,32'd-12382,32'd2844,32'd-1907,32'd1976,32'd-3146,32'd-1330,32'd1300,32'd3039,32'd2944,32'd-1472,32'd1856,32'd2479,32'd646,32'd2792,32'd-1101,32'd-5966,32'd875,32'd-3044,32'd4389,32'd-9116,32'd-29,32'd-1967,32'd-3198,32'd-7080,32'd1638,32'd-2231,32'd-3876,32'd-1724,32'd6035,32'd-603,32'd-4421,32'd-6948,32'd-2534,32'd841,32'd-2585,32'd69,32'd-539,32'd5498,32'd1276,32'd-1883,32'd-5654,32'd6538,32'd6269,32'd-1025,32'd-3371,32'd-4719,32'd-3581,32'd-1932,32'd-2409,32'd-1695,32'd1923,32'd-834,32'd-2073,32'd-1053,32'd5190,32'd-8305,32'd-1602,32'd-5400,32'd-1492,32'd304,32'd5786,32'd-1600,32'd72,32'd-4020,32'd2609,32'd680,32'd-5571,32'd6879,32'd661,32'd-3144,32'd638,32'd394,32'd-4497,32'd-1617,32'd4633,32'd-7041,32'd-10917,32'd-102,32'd5107,32'd167,32'd2861,32'd-10048,32'd449,32'd-3361,32'd6206,32'd-2619,32'd-3117,32'd-1207,32'd2210,32'd7021,32'd-5375,32'd-2807,32'd-338,32'd-5986,32'd-6909,32'd288,32'd6440,32'd-8247,32'd-6411,32'd-712,32'd-81,32'd1817,32'd711,32'd7094,32'd4560,32'd-3022,32'd2456,32'd7758,32'd1999,32'd-3708,32'd960,32'd7534,32'd6235,32'd2534,32'd-3156,32'd-4645,32'd-6684,32'd-1790,32'd4331,32'd-6660,32'd3393,32'd6137,32'd-2482,32'd-1597,32'd6298,32'd-3105,32'd-4631,32'd-14375,32'd-4843,32'd-5976,32'd-900,32'd-3449,32'd351,32'd-1192,32'd354,32'd-2393,32'd-9208,32'd-5937,32'd4382,32'd-3735,32'd-8173,32'd6215,32'd-248,32'd-7749,32'd1973,32'd1397,32'd-9169,32'd6093,32'd-3085,32'd9941,32'd5258,32'd-4912,32'd5244,32'd1992,32'd-8310,32'd-8247,32'd12412,32'd-2973,32'd2775,32'd-107,32'd6489,32'd-8051,32'd-1014,32'd385,32'd755,32'd-3889,32'd-3063,32'd-2141,32'd13271,32'd-10322,32'd2661,32'd-3298,32'd2181,32'd8203,32'd4284,32'd-8378,32'd-8774,32'd9243,32'd-3962,32'd-510,32'd9428,32'd1654,32'd-2858,32'd-262};
    Wx[92]='{32'd881,32'd-6499,32'd830,32'd966,32'd-77,32'd-1246,32'd4479,32'd366,32'd4372,32'd1365,32'd3493,32'd424,32'd-3410,32'd-5727,32'd-2403,32'd-1112,32'd4680,32'd2995,32'd-2274,32'd-2279,32'd1512,32'd2795,32'd1439,32'd1036,32'd2198,32'd-295,32'd277,32'd218,32'd2115,32'd-2927,32'd2456,32'd-6508,32'd7563,32'd2224,32'd869,32'd498,32'd-870,32'd3317,32'd-5053,32'd1330,32'd-746,32'd1375,32'd-3391,32'd-204,32'd-1954,32'd1317,32'd-5083,32'd-1918,32'd568,32'd-3894,32'd-6875,32'd-402,32'd-1624,32'd-1590,32'd4211,32'd4233,32'd2026,32'd-6640,32'd-314,32'd10351,32'd-7548,32'd-916,32'd-1491,32'd-1890,32'd-2108,32'd-870,32'd-155,32'd-6835,32'd-5590,32'd-1605,32'd-786,32'd-2453,32'd-450,32'd-1738,32'd1425,32'd-745,32'd-2148,32'd-3779,32'd-1196,32'd97,32'd-1143,32'd-11796,32'd-663,32'd3210,32'd-1011,32'd1390,32'd1083,32'd-247,32'd3017,32'd-3481,32'd-3576,32'd-3691,32'd2416,32'd-323,32'd-717,32'd-2089,32'd-6357,32'd-1205,32'd-2305,32'd-2001,32'd-1073,32'd432,32'd-5693,32'd6977,32'd2878,32'd-731,32'd-8735,32'd-5410,32'd-3156,32'd-4616,32'd-1748,32'd1612,32'd-6420,32'd-2656,32'd-7202,32'd-5874,32'd1225,32'd-540,32'd2467,32'd-5239,32'd385,32'd8872,32'd3408,32'd49,32'd-1336,32'd-5507,32'd-1340,32'd2260,32'd6005,32'd8618,32'd-5253,32'd-10927,32'd-902,32'd-14013,32'd9497,32'd6,32'd5126,32'd-2254,32'd7470,32'd8852,32'd2795,32'd-17675,32'd690,32'd3623,32'd18183,32'd-167,32'd6201,32'd-16894,32'd429,32'd-8779,32'd-5107,32'd9521,32'd9462,32'd-4487,32'd1401,32'd8071,32'd1892,32'd6835,32'd1561,32'd2783,32'd11396,32'd7153,32'd-3444,32'd-5795,32'd541,32'd3122,32'd-2219,32'd4365,32'd4484,32'd-667,32'd-14833,32'd219,32'd436,32'd-12304,32'd-1949,32'd6264,32'd1422,32'd2761,32'd-10087,32'd2370,32'd-3657,32'd21230,32'd-1853,32'd3874,32'd-5673,32'd5942,32'd-2524,32'd4951,32'd-656,32'd-5522,32'd3232,32'd-3920,32'd3500,32'd-3093,32'd-19902,32'd-2507,32'd-4020,32'd-4912,32'd383,32'd7651,32'd4150,32'd7456,32'd4372,32'd536,32'd5781,32'd-351,32'd-1249,32'd7407,32'd1492,32'd654,32'd-642,32'd-2207,32'd2083,32'd2792,32'd-1268,32'd-8173,32'd-9863,32'd-4736,32'd-1555,32'd-3342,32'd879,32'd951,32'd98,32'd-996,32'd4462,32'd3530,32'd-3188,32'd-2851,32'd-3559,32'd5961,32'd-677,32'd2274,32'd996,32'd-2717,32'd-2010,32'd-766,32'd53,32'd618,32'd-674,32'd-514,32'd5268,32'd11376,32'd4331,32'd-1550,32'd10400,32'd-2597,32'd-1507,32'd1759,32'd3989,32'd-310,32'd10722,32'd2048,32'd184,32'd-3847,32'd-5375,32'd841,32'd2666,32'd-4140,32'd-2558,32'd-10673,32'd-3710,32'd4685,32'd3891,32'd-412,32'd5952,32'd-1231,32'd-111,32'd11152,32'd-7299,32'd1150,32'd9936,32'd1378,32'd4924,32'd2680,32'd2963,32'd-300,32'd-4216,32'd1690,32'd12695,32'd2946,32'd-4003,32'd4619,32'd5512,32'd4216,32'd3803,32'd-3222,32'd1126,32'd-891,32'd470,32'd-3320,32'd-2335,32'd-2437,32'd-1472,32'd4489,32'd1878,32'd2471,32'd-3981,32'd-824,32'd4970,32'd5200,32'd6533,32'd5830,32'd-1953,32'd-767,32'd3935,32'd-1804,32'd-7563,32'd3408,32'd43,32'd-9326,32'd-1027,32'd-549,32'd-4980,32'd1622,32'd3061,32'd3149,32'd261,32'd-5761,32'd-4772,32'd-2122,32'd3244,32'd822,32'd-3115,32'd-2239,32'd9355,32'd-6469,32'd851,32'd789,32'd2546,32'd6010,32'd-2639,32'd-32,32'd-6401,32'd-5273,32'd-3015,32'd-1818,32'd-3229,32'd8266,32'd2548,32'd-1486,32'd955,32'd8046,32'd-4165,32'd-6308,32'd-271,32'd-6567,32'd1307,32'd2044,32'd3469,32'd-8056,32'd-3059,32'd-8041,32'd-4921,32'd-8164,32'd-8081,32'd1622,32'd1658,32'd-3149,32'd-4584,32'd1584,32'd-1545,32'd-1947,32'd9370,32'd794,32'd-3505,32'd11220,32'd74,32'd259,32'd2712,32'd7724,32'd-2524,32'd-590,32'd-1304,32'd1832,32'd-2150,32'd-3505,32'd-6928,32'd-4238,32'd-2108,32'd1394,32'd-3547,32'd-1920,32'd-2915,32'd1904,32'd554,32'd2902,32'd-50,32'd1577,32'd1527,32'd-4357,32'd-7773,32'd-13046,32'd6640,32'd-6479,32'd758,32'd-2983,32'd-3103,32'd10917,32'd2773,32'd-6728};
    Wx[93]='{32'd-946,32'd1133,32'd-603,32'd1163,32'd2453,32'd-1799,32'd-270,32'd2880,32'd966,32'd2324,32'd-1215,32'd494,32'd-1297,32'd-2124,32'd-160,32'd-3210,32'd-6826,32'd534,32'd-3994,32'd-4567,32'd1483,32'd2113,32'd4565,32'd4055,32'd-1259,32'd998,32'd111,32'd657,32'd-1463,32'd1912,32'd363,32'd-3405,32'd-717,32'd-3071,32'd2500,32'd1117,32'd-765,32'd874,32'd2344,32'd327,32'd1074,32'd-1430,32'd3403,32'd303,32'd-3359,32'd2216,32'd-6855,32'd4155,32'd-12,32'd-930,32'd12275,32'd1287,32'd842,32'd1741,32'd5571,32'd-2541,32'd418,32'd-1301,32'd-166,32'd-1614,32'd832,32'd-3959,32'd3527,32'd-2194,32'd-3918,32'd2573,32'd1416,32'd186,32'd-3698,32'd870,32'd-360,32'd-4091,32'd-2276,32'd-1588,32'd1629,32'd2548,32'd3962,32'd2734,32'd3935,32'd-3137,32'd2570,32'd1131,32'd3840,32'd3601,32'd3830,32'd2279,32'd-263,32'd-1881,32'd2739,32'd1488,32'd-4028,32'd-464,32'd1785,32'd-4934,32'd5629,32'd-3564,32'd-2221,32'd-6210,32'd1876,32'd757,32'd143,32'd711,32'd1431,32'd4904,32'd-3386,32'd2626,32'd2393,32'd1282,32'd4221,32'd-1689,32'd-6323,32'd-38,32'd-3298,32'd3332,32'd-8310,32'd-1165,32'd1597,32'd3991,32'd4501,32'd-2685,32'd779,32'd8208,32'd-5449,32'd-2445,32'd-3530,32'd-443,32'd-700,32'd773,32'd2236,32'd4997,32'd-1729,32'd-2727,32'd1741,32'd2073,32'd3894,32'd-23,32'd-667,32'd-184,32'd-134,32'd3398,32'd6796,32'd1000,32'd5498,32'd1287,32'd-2966,32'd5463,32'd2976,32'd-6840,32'd-1258,32'd3674,32'd-3999,32'd1359,32'd16416,32'd2907,32'd-6435,32'd5898,32'd261,32'd1694,32'd1748,32'd4052,32'd1282,32'd-7285,32'd-12431,32'd-1345,32'd-5527,32'd-1711,32'd3366,32'd-9604,32'd4655,32'd158,32'd-13828,32'd-5859,32'd-798,32'd676,32'd3798,32'd-2751,32'd-7700,32'd4602,32'd-6577,32'd5136,32'd1490,32'd14296,32'd586,32'd-8647,32'd4636,32'd2580,32'd-2980,32'd-6582,32'd-4418,32'd1815,32'd1834,32'd-5170,32'd1199,32'd-2514,32'd3400,32'd-2406,32'd9916,32'd3876,32'd-3967,32'd-2526,32'd2174,32'd5229,32'd-267,32'd-692,32'd2961,32'd-1092,32'd4721,32'd-3234,32'd1545,32'd-780,32'd-4882,32'd-3159,32'd-1434,32'd-7314,32'd5498,32'd3771,32'd-5712,32'd1837,32'd-1745,32'd-2205,32'd-794,32'd89,32'd-1904,32'd1113,32'd4379,32'd90,32'd-5693,32'd502,32'd-1210,32'd-2878,32'd4006,32'd-6391,32'd505,32'd3671,32'd-6503,32'd-1306,32'd1630,32'd-5097,32'd3435,32'd-2429,32'd-5019,32'd-1278,32'd5288,32'd-1662,32'd1428,32'd-4101,32'd2519,32'd-864,32'd-4519,32'd-1433,32'd-7861,32'd-9794,32'd7250,32'd2331,32'd3374,32'd-4514,32'd602,32'd-3979,32'd349,32'd1000,32'd-2355,32'd-2802,32'd1730,32'd-230,32'd3186,32'd-508,32'd-567,32'd9477,32'd-3764,32'd10,32'd3835,32'd2015,32'd-3903,32'd-40,32'd-36,32'd-1232,32'd-6889,32'd-1468,32'd906,32'd-849,32'd1132,32'd-5795,32'd4895,32'd-3630,32'd-1959,32'd-5219,32'd-26,32'd-772,32'd-3918,32'd-254,32'd-3227,32'd-8818,32'd-518,32'd-1237,32'd8427,32'd1875,32'd-3308,32'd-924,32'd3027,32'd-3181,32'd7797,32'd857,32'd-49,32'd2149,32'd3491,32'd-2617,32'd-534,32'd615,32'd6240,32'd-520,32'd-2032,32'd3803,32'd-473,32'd-9531,32'd2541,32'd4523,32'd1373,32'd-3125,32'd-3847,32'd-3078,32'd-2114,32'd-3569,32'd2412,32'd4653,32'd3847,32'd19,32'd-82,32'd2432,32'd6093,32'd2069,32'd2993,32'd-3847,32'd-545,32'd297,32'd-1839,32'd-2115,32'd7988,32'd-117,32'd5834,32'd-4260,32'd-2551,32'd1785,32'd-4025,32'd-6640,32'd-1207,32'd2464,32'd805,32'd4228,32'd217,32'd-3344,32'd9189,32'd-4670,32'd695,32'd487,32'd5419,32'd3789,32'd-3112,32'd-1313,32'd-1019,32'd-2883,32'd1180,32'd1345,32'd664,32'd-991,32'd-1429,32'd3698,32'd91,32'd1198,32'd-7485,32'd-6118,32'd2949,32'd-6157,32'd614,32'd238,32'd2805,32'd4677,32'd155,32'd3586,32'd2727,32'd-6499,32'd2890,32'd-4536,32'd2290,32'd-3112,32'd3132,32'd-9804,32'd-1006,32'd-1071,32'd1066,32'd532,32'd-6630,32'd-4819,32'd2834,32'd-7314,32'd897,32'd2912,32'd-6542,32'd3266,32'd2937,32'd-3950};
    Wx[94]='{32'd1278,32'd-1942,32'd-554,32'd-3161,32'd2247,32'd-1317,32'd-3459,32'd-257,32'd4523,32'd-1707,32'd53,32'd290,32'd2734,32'd1262,32'd1688,32'd-38,32'd-210,32'd2218,32'd3183,32'd-1376,32'd603,32'd-3034,32'd-1348,32'd20,32'd3537,32'd-789,32'd-402,32'd3537,32'd-47,32'd917,32'd-1695,32'd1552,32'd2556,32'd2216,32'd3493,32'd-2685,32'd-449,32'd-341,32'd1828,32'd98,32'd792,32'd32,32'd4956,32'd3322,32'd3239,32'd2700,32'd-1190,32'd-3005,32'd755,32'd1495,32'd-3547,32'd-6298,32'd-257,32'd3027,32'd-3793,32'd3896,32'd2218,32'd-2358,32'd4189,32'd8681,32'd-214,32'd-3745,32'd-4965,32'd1915,32'd-1173,32'd-2753,32'd2130,32'd1940,32'd3312,32'd-1597,32'd-1844,32'd-5380,32'd-816,32'd1743,32'd-3994,32'd1408,32'd-4055,32'd1503,32'd1008,32'd4018,32'd433,32'd4721,32'd-1651,32'd5737,32'd-1200,32'd2248,32'd2397,32'd2922,32'd-297,32'd-3989,32'd3413,32'd-4980,32'd-3823,32'd1297,32'd1866,32'd1730,32'd1078,32'd736,32'd1713,32'd-2617,32'd4973,32'd453,32'd1364,32'd8989,32'd6445,32'd1612,32'd-969,32'd5092,32'd-5922,32'd-9291,32'd103,32'd-2360,32'd-3569,32'd-6923,32'd13505,32'd-11572,32'd408,32'd-82,32'd-3020,32'd-3884,32'd-4487,32'd-9990,32'd4094,32'd-7744,32'd144,32'd7685,32'd-1816,32'd-4265,32'd-2790,32'd2905,32'd-223,32'd15332,32'd-12841,32'd12353,32'd-692,32'd8701,32'd1850,32'd4011,32'd-1209,32'd-6567,32'd-4802,32'd19033,32'd-662,32'd4726,32'd17626,32'd3452,32'd2395,32'd-2641,32'd11064,32'd-3154,32'd1138,32'd15078,32'd-2189,32'd-10781,32'd5415,32'd-2956,32'd1614,32'd-2770,32'd-12968,32'd-2471,32'd-2812,32'd-1461,32'd-5839,32'd-2237,32'd17255,32'd1453,32'd-1450,32'd1614,32'd-827,32'd-1997,32'd236,32'd709,32'd-1233,32'd8813,32'd-3725,32'd9628,32'd5830,32'd6367,32'd-1514,32'd-816,32'd6186,32'd-5864,32'd5991,32'd6982,32'd-2617,32'd-7524,32'd3007,32'd12080,32'd-578,32'd-2189,32'd2663,32'd16572,32'd1363,32'd-506,32'd6953,32'd4826,32'd-4067,32'd-1607,32'd3447,32'd7700,32'd985,32'd-2744,32'd5078,32'd-3874,32'd3183,32'd423,32'd690,32'd-1779,32'd5000,32'd4111,32'd-7021,32'd280,32'd1402,32'd2707,32'd4316,32'd2800,32'd-2156,32'd-6474,32'd-936,32'd-891,32'd-1857,32'd2624,32'd-1557,32'd-1411,32'd-1977,32'd-4519,32'd4641,32'd44,32'd8,32'd-438,32'd-2385,32'd-5405,32'd-8754,32'd918,32'd-3405,32'd2448,32'd4362,32'd2424,32'd-2922,32'd4165,32'd-3090,32'd1148,32'd-3151,32'd3540,32'd-6850,32'd-3417,32'd8378,32'd-241,32'd-4323,32'd-2318,32'd5336,32'd-3940,32'd-1689,32'd-5800,32'd1884,32'd618,32'd-87,32'd2717,32'd1844,32'd-7587,32'd-7377,32'd-586,32'd-2281,32'd-8422,32'd109,32'd-3581,32'd-2441,32'd1976,32'd-3718,32'd-820,32'd-3295,32'd-3225,32'd1063,32'd-5170,32'd-770,32'd2927,32'd-567,32'd-752,32'd11660,32'd-568,32'd1939,32'd985,32'd3256,32'd-3344,32'd4055,32'd-8,32'd1651,32'd-2509,32'd910,32'd-1806,32'd845,32'd712,32'd-5683,32'd-6611,32'd-440,32'd-426,32'd-2167,32'd-3405,32'd2178,32'd-232,32'd5751,32'd-6254,32'd522,32'd-2495,32'd2077,32'd76,32'd1253,32'd-5117,32'd3264,32'd14023,32'd-3481,32'd-2164,32'd3020,32'd-1354,32'd2658,32'd1301,32'd-3076,32'd4116,32'd-324,32'd-5600,32'd1781,32'd1573,32'd-8471,32'd-1589,32'd4223,32'd-7514,32'd7495,32'd-1718,32'd-12285,32'd-4584,32'd-4162,32'd-7880,32'd-5830,32'd-1463,32'd-1781,32'd1916,32'd5131,32'd3037,32'd-9091,32'd5400,32'd778,32'd-5297,32'd3835,32'd3093,32'd-1342,32'd-3950,32'd341,32'd3691,32'd-1328,32'd3144,32'd-4970,32'd-4313,32'd-5024,32'd-1060,32'd296,32'd328,32'd-623,32'd-5961,32'd3669,32'd-14560,32'd-3767,32'd-1231,32'd-260,32'd-8764,32'd-1912,32'd2331,32'd-2812,32'd-1763,32'd11552,32'd-9233,32'd1008,32'd-8500,32'd-6181,32'd4553,32'd1287,32'd2504,32'd-11914,32'd-4079,32'd5,32'd-896,32'd6542,32'd-6176,32'd-529,32'd-4272,32'd10000,32'd-6098,32'd4975,32'd1499,32'd-60,32'd-9023,32'd1569,32'd-2675,32'd-7221,32'd-5488,32'd-323,32'd893,32'd2364,32'd-3098,32'd4536,32'd573};
    Wx[95]='{32'd1154,32'd456,32'd1268,32'd1986,32'd2487,32'd484,32'd2968,32'd1955,32'd-2700,32'd-1417,32'd5942,32'd1501,32'd2646,32'd4343,32'd4467,32'd4575,32'd2619,32'd-2125,32'd1177,32'd4423,32'd-652,32'd2768,32'd1036,32'd4079,32'd977,32'd-720,32'd557,32'd-546,32'd11582,32'd-5864,32'd-478,32'd11894,32'd5527,32'd2731,32'd3979,32'd2132,32'd-3937,32'd1135,32'd1611,32'd-1981,32'd2193,32'd3090,32'd-1610,32'd4265,32'd-4750,32'd2071,32'd5078,32'd-11,32'd3173,32'd-126,32'd-3273,32'd-2187,32'd-1752,32'd2731,32'd-1800,32'd-3225,32'd1014,32'd76,32'd-1761,32'd222,32'd3991,32'd8037,32'd2934,32'd5991,32'd-4020,32'd620,32'd-4101,32'd4255,32'd1254,32'd-662,32'd-2243,32'd4118,32'd-1354,32'd-223,32'd1119,32'd817,32'd5781,32'd3427,32'd3359,32'd875,32'd1040,32'd14238,32'd7490,32'd-4243,32'd3022,32'd8159,32'd2078,32'd5053,32'd3161,32'd-2062,32'd-793,32'd6816,32'd5131,32'd6201,32'd2573,32'd2270,32'd1687,32'd2875,32'd2388,32'd-1205,32'd-5039,32'd-6816,32'd1176,32'd2352,32'd1768,32'd2443,32'd3720,32'd794,32'd4851,32'd-230,32'd-5898,32'd-2687,32'd2387,32'd8237,32'd7563,32'd-5498,32'd2070,32'd5146,32'd2404,32'd1857,32'd31,32'd834,32'd1510,32'd-1380,32'd-4692,32'd-2795,32'd1093,32'd667,32'd-4152,32'd-5,32'd232,32'd-11923,32'd652,32'd7690,32'd-2181,32'd11123,32'd1075,32'd4028,32'd12089,32'd-11777,32'd-6538,32'd1205,32'd1843,32'd-4987,32'd7812,32'd-6025,32'd-4633,32'd400,32'd4868,32'd5820,32'd11865,32'd7680,32'd-6035,32'd5678,32'd4160,32'd-4052,32'd-3022,32'd-1103,32'd10859,32'd-3542,32'd-321,32'd18486,32'd-4760,32'd6318,32'd8110,32'd-2941,32'd-2093,32'd8486,32'd-3608,32'd2021,32'd-637,32'd5336,32'd-1804,32'd2132,32'd2968,32'd-9047,32'd3339,32'd5073,32'd-3857,32'd-3127,32'd-6035,32'd-15634,32'd4313,32'd1633,32'd1997,32'd-5615,32'd2199,32'd3122,32'd-3286,32'd-1113,32'd-3251,32'd-1630,32'd-2832,32'd553,32'd-873,32'd8642,32'd-3381,32'd1968,32'd6347,32'd-911,32'd-4160,32'd-2836,32'd941,32'd5312,32'd-1170,32'd928,32'd-3735,32'd-2573,32'd-1927,32'd-1431,32'd-322,32'd-3059,32'd-3093,32'd3413,32'd-3962,32'd-3845,32'd-1783,32'd-1801,32'd-1597,32'd744,32'd1585,32'd1356,32'd-2644,32'd-2218,32'd2059,32'd-2283,32'd5151,32'd2958,32'd857,32'd8291,32'd125,32'd820,32'd929,32'd2210,32'd5512,32'd897,32'd-526,32'd2371,32'd2196,32'd1541,32'd-2205,32'd-5117,32'd-472,32'd9150,32'd1571,32'd-1976,32'd3269,32'd257,32'd-1133,32'd4060,32'd-2424,32'd1199,32'd-2283,32'd-4038,32'd-1529,32'd-1455,32'd-6748,32'd2130,32'd5815,32'd-4372,32'd1136,32'd3322,32'd-513,32'd-5629,32'd6093,32'd450,32'd1395,32'd10351,32'd-1005,32'd-263,32'd4277,32'd1734,32'd2076,32'd992,32'd2443,32'd2207,32'd4978,32'd-6430,32'd7915,32'd283,32'd1978,32'd8471,32'd3937,32'd-6538,32'd4296,32'd6547,32'd-1485,32'd657,32'd2419,32'd-5507,32'd-961,32'd681,32'd3107,32'd-504,32'd-4191,32'd-1273,32'd5034,32'd-3715,32'd3405,32'd-1072,32'd-5644,32'd2270,32'd5107,32'd-2993,32'd174,32'd-738,32'd-567,32'd1032,32'd-3737,32'd-3217,32'd11269,32'd1427,32'd2250,32'd10283,32'd3520,32'd-1223,32'd3430,32'd6186,32'd-4709,32'd7387,32'd4960,32'd-3178,32'd-2261,32'd3371,32'd-4677,32'd145,32'd5502,32'd3688,32'd9169,32'd1954,32'd2536,32'd4895,32'd333,32'd3625,32'd1320,32'd546,32'd96,32'd-1307,32'd-3298,32'd3654,32'd-3442,32'd75,32'd596,32'd3076,32'd6230,32'd-1224,32'd-562,32'd-737,32'd-6411,32'd-240,32'd-3820,32'd-1768,32'd1884,32'd-6220,32'd-2277,32'd-6142,32'd-5449,32'd9667,32'd-386,32'd-8999,32'd637,32'd5380,32'd-4160,32'd1087,32'd-2167,32'd4208,32'd3793,32'd5395,32'd-5205,32'd3554,32'd-2301,32'd1928,32'd8789,32'd-5039,32'd6635,32'd5742,32'd1044,32'd-89,32'd-750,32'd997,32'd5634,32'd230,32'd2059,32'd-6259,32'd7695,32'd1888,32'd2207,32'd1911,32'd-2583,32'd3122,32'd260,32'd1068,32'd1282,32'd13134,32'd1628,32'd93,32'd6806,32'd3405,32'd2143,32'd-907};
    Wx[96]='{32'd-952,32'd-673,32'd2875,32'd2812,32'd1784,32'd-1928,32'd-3164,32'd3093,32'd2541,32'd-178,32'd-919,32'd1201,32'd237,32'd-1749,32'd100,32'd7221,32'd-299,32'd1190,32'd-5742,32'd3669,32'd-3493,32'd1835,32'd-2167,32'd7651,32'd2117,32'd2215,32'd3325,32'd-940,32'd980,32'd-6914,32'd95,32'd274,32'd-5454,32'd2282,32'd-88,32'd1452,32'd-3901,32'd-2368,32'd440,32'd4672,32'd-1342,32'd1021,32'd3740,32'd-1611,32'd-2064,32'd-5385,32'd-7294,32'd2145,32'd-4094,32'd2227,32'd-2800,32'd-1674,32'd-34,32'd4602,32'd-2026,32'd-2143,32'd1354,32'd1133,32'd-1345,32'd-5600,32'd2468,32'd-3723,32'd-2352,32'd3112,32'd5732,32'd3400,32'd543,32'd4516,32'd3481,32'd-160,32'd3125,32'd-3127,32'd-3134,32'd-2122,32'd877,32'd7675,32'd-1157,32'd-2116,32'd5078,32'd-4199,32'd1954,32'd-7426,32'd-672,32'd-585,32'd-6040,32'd-6284,32'd-1169,32'd699,32'd2109,32'd-232,32'd-3303,32'd1785,32'd-2675,32'd-3132,32'd-258,32'd-1823,32'd239,32'd-708,32'd-150,32'd-2612,32'd-4855,32'd-2783,32'd-4025,32'd4802,32'd-1381,32'd-2149,32'd6997,32'd4462,32'd-1533,32'd-259,32'd13955,32'd6342,32'd4863,32'd2006,32'd4658,32'd3955,32'd1677,32'd5083,32'd-2072,32'd4768,32'd-3916,32'd7065,32'd-7358,32'd1079,32'd-1782,32'd11503,32'd-2236,32'd-2197,32'd-2106,32'd-2432,32'd-4462,32'd-2646,32'd-15517,32'd8378,32'd-1400,32'd5917,32'd2863,32'd-2919,32'd-7211,32'd-2724,32'd-6083,32'd-10605,32'd-1018,32'd-1524,32'd-2380,32'd2435,32'd14140,32'd6015,32'd4301,32'd4343,32'd-5014,32'd20761,32'd7431,32'd-4077,32'd428,32'd9838,32'd-5493,32'd-1475,32'd-12158,32'd1650,32'd-4213,32'd-610,32'd-1582,32'd4599,32'd8310,32'd-4287,32'd1434,32'd-4582,32'd1127,32'd-2526,32'd1486,32'd5893,32'd-2014,32'd3500,32'd-7148,32'd-255,32'd-2430,32'd-5664,32'd15029,32'd-1563,32'd2354,32'd29726,32'd646,32'd-8750,32'd1502,32'd-12910,32'd-3974,32'd1347,32'd-4355,32'd5551,32'd-1859,32'd13818,32'd-3593,32'd1463,32'd3005,32'd7446,32'd5849,32'd-9863,32'd-1431,32'd7734,32'd3881,32'd232,32'd2746,32'd93,32'd5966,32'd-1007,32'd-465,32'd-8115,32'd-7026,32'd-3742,32'd-6308,32'd-4558,32'd-845,32'd-950,32'd1215,32'd3647,32'd-4536,32'd-2519,32'd-2133,32'd-125,32'd571,32'd1535,32'd-3483,32'd1815,32'd-1265,32'd-5004,32'd-4277,32'd-1613,32'd-3056,32'd7016,32'd2413,32'd2263,32'd1875,32'd-4799,32'd2423,32'd-665,32'd-2990,32'd1916,32'd-440,32'd2846,32'd997,32'd-1549,32'd-8330,32'd-8315,32'd-2644,32'd1375,32'd-5532,32'd-1928,32'd9067,32'd-418,32'd-762,32'd4252,32'd177,32'd-4025,32'd-2283,32'd4267,32'd-3449,32'd-1171,32'd-2437,32'd-996,32'd5751,32'd-8935,32'd-967,32'd2661,32'd6674,32'd-1524,32'd155,32'd1079,32'd1365,32'd-3073,32'd-1422,32'd-994,32'd-919,32'd-1149,32'd-4653,32'd-8588,32'd648,32'd-6425,32'd-6791,32'd-386,32'd669,32'd-4560,32'd-4453,32'd-897,32'd21,32'd-7851,32'd-1566,32'd-4067,32'd-2919,32'd-1182,32'd5205,32'd-1682,32'd-364,32'd-664,32'd823,32'd-2858,32'd5317,32'd1901,32'd-3815,32'd-4597,32'd3166,32'd-9028,32'd-563,32'd-6704,32'd6074,32'd-6694,32'd-725,32'd3642,32'd-2968,32'd-2939,32'd1733,32'd-3186,32'd3706,32'd-8134,32'd-3566,32'd925,32'd-8476,32'd-1583,32'd1102,32'd671,32'd-6230,32'd95,32'd4250,32'd6240,32'd-355,32'd6186,32'd-1440,32'd-692,32'd-1921,32'd95,32'd-106,32'd-5791,32'd-4548,32'd-10781,32'd-1888,32'd-2675,32'd-3056,32'd-4313,32'd-4799,32'd4987,32'd2646,32'd914,32'd5688,32'd-15644,32'd-8886,32'd1531,32'd-1452,32'd1166,32'd-1073,32'd-930,32'd-3337,32'd-11572,32'd-2255,32'd-880,32'd1967,32'd7646,32'd-1192,32'd4311,32'd-2160,32'd1766,32'd5449,32'd-7714,32'd-3320,32'd-3735,32'd2177,32'd-7182,32'd2666,32'd-5312,32'd-4904,32'd-1866,32'd-2307,32'd-192,32'd-839,32'd-3225,32'd-3041,32'd-1793,32'd-3732,32'd-9995,32'd-3684,32'd2292,32'd1303,32'd-7265,32'd6914,32'd-3090,32'd-2624,32'd-1568,32'd966,32'd-3237,32'd-625,32'd1511,32'd-2307,32'd-7680,32'd-4990,32'd5429,32'd2614,32'd-8686,32'd-2619,32'd5493,32'd1429,32'd-5161};
    Wx[97]='{32'd3718,32'd5190,32'd1887,32'd-1628,32'd-1796,32'd-2110,32'd1901,32'd1026,32'd-2890,32'd841,32'd4128,32'd-605,32'd1130,32'd1325,32'd2277,32'd-1851,32'd7124,32'd136,32'd-78,32'd3039,32'd-1431,32'd-3261,32'd-657,32'd-370,32'd2326,32'd-1536,32'd4650,32'd1239,32'd2276,32'd-1745,32'd87,32'd7631,32'd-1069,32'd960,32'd4973,32'd1124,32'd2709,32'd4272,32'd2814,32'd2467,32'd1699,32'd-1773,32'd-266,32'd6386,32'd-9995,32'd-4685,32'd-1133,32'd-321,32'd-3061,32'd-605,32'd-292,32'd-4450,32'd-4868,32'd-2277,32'd3103,32'd3947,32'd-1860,32'd75,32'd-1248,32'd-1978,32'd1095,32'd2575,32'd151,32'd-3911,32'd-5058,32'd-3376,32'd1370,32'd1005,32'd-2619,32'd-2634,32'd692,32'd2805,32'd5463,32'd-3452,32'd-1910,32'd2736,32'd3,32'd-1606,32'd-2066,32'd1501,32'd-1497,32'd6894,32'd-1549,32'd-3320,32'd-957,32'd-6357,32'd-2949,32'd-674,32'd-3339,32'd524,32'd-393,32'd2822,32'd-5952,32'd-3671,32'd-538,32'd2150,32'd1195,32'd-2634,32'd-2995,32'd3208,32'd4140,32'd9384,32'd-1408,32'd-637,32'd1227,32'd2041,32'd192,32'd-4924,32'd623,32'd-5249,32'd-6323,32'd422,32'd-2746,32'd-3049,32'd4414,32'd-7568,32'd5009,32'd10400,32'd-1330,32'd1833,32'd-4221,32'd-879,32'd4091,32'd1870,32'd199,32'd3676,32'd-745,32'd1197,32'd-16318,32'd4521,32'd5947,32'd6630,32'd21601,32'd495,32'd3103,32'd2387,32'd2749,32'd11582,32'd3247,32'd-9091,32'd-9936,32'd65,32'd3657,32'd5434,32'd9663,32'd9604,32'd3769,32'd-11621,32'd-8183,32'd8305,32'd11669,32'd3093,32'd-7021,32'd10205,32'd933,32'd-8701,32'd554,32'd2624,32'd6132,32'd3916,32'd-5122,32'd-3374,32'd1021,32'd2180,32'd-1942,32'd3630,32'd3027,32'd6831,32'd-2194,32'd-877,32'd12832,32'd-4401,32'd-1375,32'd-7592,32'd-961,32'd7783,32'd15859,32'd-2819,32'd5039,32'd-3635,32'd-7299,32'd729,32'd10078,32'd5717,32'd4741,32'd-5917,32'd5551,32'd332,32'd2318,32'd-563,32'd855,32'd-1958,32'd19619,32'd-1345,32'd-9091,32'd7133,32'd-6845,32'd-15527,32'd3125,32'd-7021,32'd-950,32'd-1113,32'd1445,32'd3381,32'd-2174,32'd-2120,32'd4340,32'd-1114,32'd1658,32'd-3496,32'd1674,32'd4775,32'd-5678,32'd592,32'd-4709,32'd-3015,32'd2817,32'd4667,32'd7709,32'd1660,32'd1403,32'd2741,32'd1303,32'd428,32'd-1092,32'd-675,32'd2066,32'd-2077,32'd5141,32'd-3527,32'd656,32'd-733,32'd4802,32'd-10429,32'd3483,32'd2998,32'd-1190,32'd3010,32'd-223,32'd2695,32'd-1231,32'd-7148,32'd-2347,32'd-1947,32'd2125,32'd-1547,32'd10410,32'd1469,32'd-2797,32'd3894,32'd7329,32'd4919,32'd-298,32'd7631,32'd-1363,32'd-5737,32'd4216,32'd4853,32'd-6801,32'd-2360,32'd479,32'd3659,32'd-3735,32'd-3547,32'd-473,32'd-4770,32'd-2976,32'd-5478,32'd-4111,32'd-597,32'd-1881,32'd-1501,32'd-277,32'd-943,32'd-843,32'd4328,32'd2200,32'd1820,32'd7329,32'd4047,32'd-1179,32'd3017,32'd1194,32'd3530,32'd-3352,32'd-312,32'd-847,32'd3356,32'd1629,32'd903,32'd-6679,32'd6030,32'd2319,32'd2919,32'd-3930,32'd881,32'd-9462,32'd2204,32'd-2988,32'd314,32'd-2127,32'd1761,32'd10478,32'd4187,32'd-1043,32'd-8066,32'd4238,32'd917,32'd-476,32'd-1884,32'd5502,32'd-691,32'd2639,32'd5175,32'd-3916,32'd-1914,32'd4807,32'd7988,32'd-5810,32'd-574,32'd2274,32'd3569,32'd-6098,32'd-2021,32'd-471,32'd2841,32'd5844,32'd-1499,32'd6157,32'd-4196,32'd617,32'd-2213,32'd1602,32'd-7460,32'd7529,32'd2290,32'd6835,32'd844,32'd1522,32'd-1663,32'd-644,32'd-919,32'd-4816,32'd6992,32'd3195,32'd-4550,32'd-2033,32'd-6069,32'd-500,32'd-908,32'd4108,32'd6630,32'd-279,32'd3991,32'd11552,32'd516,32'd2110,32'd-5795,32'd-2166,32'd4230,32'd4797,32'd678,32'd-4914,32'd2198,32'd2016,32'd365,32'd-5864,32'd6069,32'd-897,32'd-8061,32'd-7680,32'd484,32'd-3771,32'd404,32'd392,32'd8896,32'd-210,32'd-974,32'd-863,32'd5131,32'd-5136,32'd-2198,32'd2587,32'd5527,32'd5600,32'd6494,32'd-1436,32'd4694,32'd501,32'd663,32'd1492,32'd599,32'd-3112,32'd2863,32'd-57,32'd4719,32'd-7211,32'd2556,32'd-3859,32'd3713};
    Wx[98]='{32'd87,32'd-5517,32'd-1716,32'd991,32'd2712,32'd2304,32'd-54,32'd-6552,32'd-1965,32'd334,32'd1790,32'd-1761,32'd-1981,32'd-1112,32'd-4191,32'd-6542,32'd403,32'd-3342,32'd-1156,32'd6225,32'd1351,32'd828,32'd-242,32'd3237,32'd-2814,32'd476,32'd2322,32'd-405,32'd-718,32'd-3129,32'd-3833,32'd-3212,32'd-1466,32'd-2536,32'd-2027,32'd-1280,32'd-1595,32'd1851,32'd-1979,32'd-2631,32'd-1455,32'd-2519,32'd-2077,32'd-6171,32'd-5322,32'd-6235,32'd-1065,32'd-5981,32'd1170,32'd-1447,32'd-4301,32'd481,32'd1678,32'd830,32'd3159,32'd-10576,32'd656,32'd4814,32'd-809,32'd-4069,32'd1711,32'd-662,32'd-1097,32'd-7905,32'd-1110,32'd4428,32'd-1973,32'd-2707,32'd3654,32'd2381,32'd4482,32'd-5751,32'd-2524,32'd2125,32'd762,32'd-902,32'd-3874,32'd-10996,32'd2609,32'd-1534,32'd-5419,32'd-3088,32'd7133,32'd-225,32'd-7001,32'd-6333,32'd-1179,32'd-1866,32'd68,32'd3728,32'd-4130,32'd212,32'd-1236,32'd21,32'd1679,32'd4707,32'd-8662,32'd-7377,32'd-3708,32'd-3693,32'd-1976,32'd5639,32'd3339,32'd2561,32'd2470,32'd-2546,32'd2990,32'd19121,32'd-3598,32'd3649,32'd4804,32'd-1625,32'd1462,32'd-6074,32'd3376,32'd-2678,32'd883,32'd800,32'd6542,32'd8056,32'd-1604,32'd656,32'd-1689,32'd4570,32'd-9448,32'd4304,32'd-4638,32'd817,32'd70,32'd6840,32'd-4589,32'd8334,32'd-24941,32'd326,32'd-1522,32'd4421,32'd188,32'd6708,32'd-1127,32'd23632,32'd3388,32'd4011,32'd-2208,32'd7895,32'd6508,32'd-914,32'd9121,32'd11953,32'd3730,32'd1381,32'd10458,32'd12949,32'd2543,32'd8876,32'd-1719,32'd10722,32'd-2459,32'd2020,32'd-3071,32'd-501,32'd4296,32'd-4409,32'd-10224,32'd10791,32'd2668,32'd-1726,32'd-1244,32'd-23261,32'd-3439,32'd2207,32'd-9956,32'd-3786,32'd-1922,32'd-902,32'd1654,32'd-12519,32'd1743,32'd-1026,32'd3276,32'd8369,32'd79,32'd4382,32'd-4572,32'd-15810,32'd271,32'd7827,32'd-8427,32'd661,32'd-7421,32'd2573,32'd9833,32'd22480,32'd-9433,32'd2093,32'd-9501,32'd-1096,32'd-6210,32'd-10166,32'd-910,32'd-17060,32'd2294,32'd112,32'd-4633,32'd2077,32'd2384,32'd-358,32'd5424,32'd2922,32'd-2166,32'd-4897,32'd-5234,32'd1822,32'd3413,32'd792,32'd182,32'd8510,32'd-6171,32'd-1605,32'd276,32'd2583,32'd-2152,32'd-218,32'd1273,32'd-2093,32'd1536,32'd5473,32'd-3242,32'd3483,32'd-4763,32'd-1567,32'd3041,32'd-5649,32'd-2683,32'd-10039,32'd1751,32'd9560,32'd6811,32'd-1248,32'd4409,32'd4238,32'd-768,32'd6328,32'd3923,32'd-6997,32'd2683,32'd3354,32'd7148,32'd-2338,32'd3757,32'd3940,32'd-4733,32'd1000,32'd696,32'd1850,32'd-564,32'd3996,32'd-4807,32'd3959,32'd-709,32'd3950,32'd-1244,32'd-6630,32'd-404,32'd-8125,32'd-2291,32'd-1904,32'd1198,32'd6069,32'd4165,32'd1901,32'd6127,32'd-3427,32'd-4301,32'd-2186,32'd407,32'd580,32'd3432,32'd532,32'd3823,32'd34,32'd-614,32'd-4208,32'd1979,32'd3740,32'd-1876,32'd-1634,32'd-592,32'd505,32'd-1409,32'd-1909,32'd653,32'd-2366,32'd-1860,32'd-2519,32'd-8491,32'd-7836,32'd3432,32'd-4887,32'd5083,32'd-10048,32'd-4941,32'd-12333,32'd-950,32'd-7036,32'd2081,32'd6772,32'd2973,32'd4147,32'd-4123,32'd-9873,32'd-6762,32'd-3330,32'd8808,32'd-1561,32'd927,32'd-1035,32'd-3928,32'd-9116,32'd-2863,32'd-1157,32'd-1508,32'd-3518,32'd-5737,32'd1082,32'd102,32'd-2993,32'd2749,32'd7412,32'd-5561,32'd-2414,32'd-7373,32'd-6020,32'd-3925,32'd-17978,32'd1225,32'd-75,32'd-5566,32'd4704,32'd396,32'd-3918,32'd1835,32'd19,32'd-2985,32'd-9267,32'd-6879,32'd56,32'd3027,32'd650,32'd3208,32'd-3254,32'd-13212,32'd-1862,32'd-5312,32'd-2668,32'd8320,32'd-2192,32'd-7890,32'd525,32'd-2663,32'd6206,32'd8193,32'd-7187,32'd-1832,32'd-9462,32'd-6137,32'd770,32'd5673,32'd-3840,32'd21210,32'd-1370,32'd13,32'd-5341,32'd3552,32'd-11289,32'd8544,32'd-2382,32'd-1158,32'd-10273,32'd-5610,32'd8300,32'd-2915,32'd-5717,32'd7314,32'd-11376,32'd-2600,32'd-6987,32'd2485,32'd-6445,32'd-662,32'd2088,32'd567,32'd-260,32'd-6220,32'd12910,32'd-7202,32'd-4785,32'd-14873,32'd7817,32'd4604,32'd-6708};
    Wx[99]='{32'd0,32'd-7602,32'd-2697,32'd-443,32'd1141,32'd1296,32'd-1783,32'd-1112,32'd400,32'd415,32'd-2327,32'd153,32'd-563,32'd1846,32'd-5488,32'd-5634,32'd-360,32'd14,32'd-5288,32'd-829,32'd-4489,32'd1727,32'd125,32'd1754,32'd-3996,32'd-1535,32'd-1577,32'd-1745,32'd-149,32'd290,32'd-5390,32'd-2209,32'd-1810,32'd-378,32'd724,32'd-507,32'd1100,32'd1977,32'd-68,32'd-388,32'd-2863,32'd-1740,32'd586,32'd-3640,32'd-2493,32'd-1866,32'd-1348,32'd-295,32'd-3247,32'd-264,32'd-1042,32'd491,32'd-828,32'd-3513,32'd2568,32'd-6806,32'd-3579,32'd1732,32'd-603,32'd-2067,32'd-3486,32'd-2042,32'd126,32'd-1699,32'd1423,32'd2056,32'd-2634,32'd-4362,32'd2320,32'd463,32'd-1973,32'd-8056,32'd-6606,32'd-2125,32'd-747,32'd-1213,32'd-992,32'd-591,32'd251,32'd1864,32'd1700,32'd4829,32'd457,32'd744,32'd-277,32'd-897,32'd-3154,32'd121,32'd-2998,32'd-1557,32'd-43,32'd2521,32'd-366,32'd57,32'd-3884,32'd-1716,32'd-123,32'd-1049,32'd-1767,32'd141,32'd1118,32'd5976,32'd1807,32'd-3088,32'd-10214,32'd-1951,32'd-1481,32'd-1502,32'd2905,32'd-853,32'd-456,32'd-341,32'd4580,32'd6254,32'd-10507,32'd4501,32'd4860,32'd-3969,32'd1982,32'd3044,32'd-2575,32'd-2949,32'd-1315,32'd-1212,32'd-950,32'd-5810,32'd1614,32'd4150,32'd3237,32'd-5200,32'd1518,32'd190,32'd4799,32'd-7358,32'd-4174,32'd-2883,32'd1636,32'd-5537,32'd15019,32'd-4580,32'd195,32'd2744,32'd-3576,32'd12802,32'd-3481,32'd3037,32'd3337,32'd3632,32'd-3820,32'd2687,32'd8784,32'd10517,32'd2358,32'd6650,32'd-5273,32'd-2252,32'd-3146,32'd-1790,32'd2449,32'd-5834,32'd6606,32'd-10595,32'd-13613,32'd1555,32'd10302,32'd-5322,32'd8774,32'd-6010,32'd-5234,32'd-1428,32'd-3239,32'd995,32'd-6250,32'd77,32'd3566,32'd-8178,32'd-2827,32'd-2778,32'd4047,32'd1341,32'd5996,32'd3017,32'd4306,32'd-13515,32'd3991,32'd-2734,32'd-8481,32'd-1158,32'd1275,32'd19,32'd307,32'd-808,32'd-5356,32'd7011,32'd11845,32'd-10185,32'd-2497,32'd1068,32'd5053,32'd2355,32'd-3066,32'd-10517,32'd-876,32'd986,32'd-2038,32'd2141,32'd2956,32'd835,32'd3498,32'd-779,32'd-612,32'd1542,32'd6894,32'd3828,32'd-152,32'd-5883,32'd4260,32'd-114,32'd2690,32'd842,32'd-2568,32'd-3811,32'd2186,32'd-1673,32'd-1174,32'd1539,32'd2622,32'd2656,32'd2812,32'd-710,32'd-1730,32'd-5629,32'd-10605,32'd11191,32'd222,32'd-6035,32'd-10078,32'd-8413,32'd4143,32'd4604,32'd-329,32'd6767,32'd982,32'd11025,32'd527,32'd-6005,32'd17119,32'd3742,32'd3508,32'd3149,32'd2080,32'd11279,32'd1481,32'd7041,32'd2805,32'd8227,32'd-7939,32'd4233,32'd1612,32'd9833,32'd-3659,32'd-1578,32'd7182,32'd-145,32'd8867,32'd-2746,32'd-359,32'd6616,32'd5439,32'd2563,32'd-2414,32'd1064,32'd-7250,32'd-577,32'd-2252,32'd722,32'd2108,32'd123,32'd-1982,32'd-1748,32'd2237,32'd-5493,32'd-2810,32'd3066,32'd-7382,32'd1713,32'd3076,32'd2722,32'd784,32'd802,32'd-7412,32'd-962,32'd-3925,32'd3596,32'd419,32'd1516,32'd-756,32'd6835,32'd3281,32'd3122,32'd-8378,32'd318,32'd2261,32'd-2646,32'd-9848,32'd-274,32'd-2636,32'd-1668,32'd-1524,32'd-2031,32'd-7104,32'd3527,32'd1087,32'd-1710,32'd-661,32'd1892,32'd-1572,32'd-6396,32'd-6606,32'd-958,32'd-12998,32'd-4206,32'd-200,32'd-1390,32'd-4760,32'd-81,32'd1096,32'd-100,32'd8037,32'd-3078,32'd-4267,32'd-1982,32'd-12685,32'd7553,32'd-7758,32'd-6738,32'd-3234,32'd-3127,32'd3056,32'd2286,32'd3625,32'd8627,32'd5556,32'd7514,32'd126,32'd-1710,32'd8159,32'd-2044,32'd-45,32'd-802,32'd-2476,32'd7124,32'd-1854,32'd-1022,32'd7348,32'd534,32'd-8432,32'd1979,32'd4108,32'd3161,32'd999,32'd695,32'd8178,32'd-570,32'd6088,32'd-847,32'd2005,32'd-2585,32'd15849,32'd4685,32'd-6787,32'd-2561,32'd-1418,32'd-2314,32'd-3957,32'd5546,32'd2941,32'd416,32'd-6567,32'd2266,32'd2626,32'd3610,32'd7016,32'd2968,32'd-2287,32'd4069,32'd5957,32'd1622,32'd-2919,32'd5771,32'd-3891,32'd5976,32'd-4685,32'd17724,32'd-7036,32'd4570,32'd2709,32'd3901,32'd2949,32'd4821};
Wh[0]='{32'd-639,32'd1331,32'd3195,32'd1979,32'd-1818,32'd-1262,32'd-5014,32'd-3674,32'd-2246,32'd218,32'd110,32'd-212,32'd1027,32'd939,32'd9321,32'd730,32'd-2362,32'd-1622,32'd771,32'd-3691,32'd2604,32'd1707,32'd-1196,32'd37,32'd1533,32'd-171,32'd-3359,32'd1143,32'd-4443,32'd-1948,32'd-1206,32'd582,32'd-327,32'd3024,32'd-325,32'd-653,32'd4538,32'd1918,32'd146,32'd1809,32'd-4106,32'd1563,32'd-10683,32'd2702,32'd2073,32'd1412,32'd3740,32'd6674,32'd728,32'd-625,32'd-6787,32'd948,32'd3337,32'd-2044,32'd1254,32'd4880,32'd700,32'd2514,32'd-371,32'd-1955,32'd-5087,32'd-2167,32'd-2509,32'd54,32'd-125,32'd-653,32'd-1619,32'd3762,32'd1617,32'd-1341,32'd344,32'd-66,32'd886,32'd1839,32'd4003,32'd-1707,32'd-461,32'd751,32'd-1530,32'd-1618,32'd1468,32'd5327,32'd-2990,32'd2753,32'd-3623,32'd1536,32'd733,32'd1706,32'd-2362,32'd-4777,32'd-2553,32'd-1270,32'd-571,32'd-2322,32'd-2839,32'd-2497,32'd374,32'd4614,32'd-1005,32'd2006,32'd-1992,32'd2205,32'd-2565,32'd3779,32'd-372,32'd1890,32'd-2480,32'd-2985,32'd-557,32'd628,32'd3605,32'd-329,32'd3540,32'd22,32'd3305,32'd-934,32'd-2113,32'd-9125,32'd-1254,32'd-4633,32'd-3681,32'd-1566,32'd1905,32'd1395,32'd52,32'd4841,32'd2489,32'd606,32'd-4311,32'd-3842,32'd-1079,32'd-1669,32'd-3510,32'd-150,32'd-751,32'd-2707,32'd-1834,32'd2174,32'd2673,32'd1483,32'd-6191,32'd965,32'd-4064,32'd-1433,32'd-438,32'd-1629,32'd-1484,32'd3874,32'd-3515,32'd2900,32'd-590,32'd2866,32'd3879,32'd2678,32'd-5136,32'd-4658,32'd-1062,32'd-397,32'd-2015,32'd183,32'd-4951,32'd-1062,32'd3095,32'd4150,32'd-815,32'd3662,32'd4252,32'd-13,32'd-954,32'd-2337,32'd3945,32'd3710,32'd1706,32'd1744,32'd-4914,32'd4248,32'd593,32'd-423,32'd-1060,32'd-219,32'd-1979,32'd-5371,32'd3764,32'd649,32'd2342,32'd660,32'd2841,32'd-1496,32'd-7802,32'd-4592,32'd1066,32'd-680,32'd1334,32'd-3076,32'd-704,32'd-2702,32'd-72,32'd329,32'd-1895,32'd-830,32'd3037,32'd1015,32'd2607,32'd-5849,32'd2590,32'd-666,32'd-1535,32'd5126,32'd2030,32'd990,32'd7050,32'd307,32'd2261,32'd-4904,32'd-3491,32'd-1177,32'd-1842,32'd2449,32'd4504,32'd-1452,32'd2481,32'd-1495,32'd-2473,32'd3972,32'd-339,32'd3876,32'd3344,32'd1536,32'd-1584,32'd3173,32'd2061,32'd-6132,32'd1099,32'd-938,32'd2819,32'd171,32'd-1054,32'd446,32'd-1343,32'd-2900,32'd4309,32'd-3391,32'd1835,32'd-3588,32'd-1284,32'd-4704,32'd-1397,32'd769,32'd-806,32'd5776,32'd-2347,32'd784,32'd2941,32'd-314,32'd-1849,32'd3149,32'd4396,32'd1118,32'd-1662,32'd-662,32'd2832,32'd-2054,32'd563,32'd3115,32'd-2115,32'd-942,32'd1730,32'd3576,32'd2937,32'd-990,32'd1046,32'd878,32'd3962,32'd-1666,32'd549,32'd3356,32'd664,32'd-470,32'd527,32'd-3188,32'd1059,32'd-3964,32'd1763,32'd-3452,32'd-573,32'd-1571,32'd-2939,32'd614,32'd401,32'd-3063,32'd5126,32'd-557,32'd473,32'd2362,32'd-1123,32'd3576,32'd-245,32'd9,32'd4736,32'd-3210,32'd4929,32'd1600,32'd949,32'd552,32'd1483,32'd3535,32'd2949,32'd-2902,32'd-609,32'd2790,32'd2003,32'd-261,32'd-2287,32'd2414,32'd376,32'd2091,32'd-3349,32'd-699,32'd6455,32'd299,32'd5502,32'd304,32'd-3913,32'd-907,32'd5126,32'd368,32'd443,32'd536,32'd1265,32'd-648,32'd2347,32'd-1766,32'd-6059,32'd230,32'd-1511,32'd6147,32'd4980,32'd4731,32'd1163,32'd-1485,32'd2639,32'd1617,32'd-5385,32'd-4829,32'd-6738,32'd-3688,32'd-7099,32'd159,32'd-1740,32'd-250,32'd1582,32'd1871,32'd393,32'd1245,32'd1171,32'd-3242,32'd2595,32'd4182,32'd-251,32'd-158,32'd-3398,32'd-2226,32'd-1765,32'd4042,32'd-1365,32'd-960,32'd3183,32'd4433,32'd-855,32'd2849,32'd-1947,32'd-2033,32'd1954,32'd5541,32'd6259,32'd132,32'd-726,32'd-2105,32'd-1928,32'd-2321,32'd-1396,32'd-1018,32'd1026,32'd-1156,32'd-2254,32'd1234,32'd1253,32'd1365,32'd-817,32'd2915,32'd-1474,32'd4438,32'd906,32'd-2489,32'd-2368,32'd2054,32'd-2452,32'd-1568,32'd2687,32'd223};
    Wh[1]='{32'd-41,32'd-439,32'd-3120,32'd-6069,32'd139,32'd5219,32'd-13271,32'd-5351,32'd-320,32'd581,32'd-5214,32'd6064,32'd3962,32'd-8251,32'd-4792,32'd-1395,32'd-3481,32'd-2030,32'd3308,32'd-2108,32'd-94,32'd1506,32'd2390,32'd-6733,32'd275,32'd-9199,32'd-5810,32'd859,32'd672,32'd-4895,32'd1300,32'd2141,32'd-3911,32'd-4631,32'd922,32'd3476,32'd1683,32'd-985,32'd-1101,32'd2496,32'd-3486,32'd-4750,32'd1383,32'd-9448,32'd-2536,32'd3354,32'd-10781,32'd-564,32'd4035,32'd-3315,32'd1959,32'd227,32'd544,32'd-2512,32'd-7763,32'd-14179,32'd2646,32'd-4597,32'd-3898,32'd8574,32'd94,32'd-3156,32'd-5839,32'd-25,32'd1602,32'd-3144,32'd-3139,32'd2465,32'd-7128,32'd-596,32'd-3349,32'd-5712,32'd1331,32'd6723,32'd676,32'd-1914,32'd-1097,32'd-6928,32'd-4348,32'd726,32'd3425,32'd-6191,32'd-4062,32'd5468,32'd2978,32'd4841,32'd642,32'd-2248,32'd-7534,32'd1535,32'd-5146,32'd385,32'd2839,32'd-3525,32'd-720,32'd3303,32'd-3625,32'd87,32'd-1174,32'd864,32'd-671,32'd-4992,32'd-679,32'd2670,32'd5258,32'd-526,32'd-5380,32'd1005,32'd15136,32'd-5473,32'd-3076,32'd4702,32'd-2414,32'd-3666,32'd-2902,32'd-839,32'd-718,32'd2142,32'd1301,32'd-4057,32'd51,32'd-2956,32'd-876,32'd147,32'd-1152,32'd-5205,32'd-9106,32'd3339,32'd-741,32'd4394,32'd4035,32'd-1785,32'd-4167,32'd1596,32'd211,32'd-11132,32'd6235,32'd-645,32'd-4230,32'd3049,32'd19248,32'd3752,32'd5336,32'd-4379,32'd261,32'd-9243,32'd5009,32'd-15976,32'd-5292,32'd-12,32'd-7124,32'd1700,32'd-708,32'd-1461,32'd-1464,32'd-6342,32'd6630,32'd3188,32'd-1793,32'd-17646,32'd16953,32'd-9169,32'd-2661,32'd-1024,32'd-4172,32'd736,32'd3874,32'd3789,32'd2265,32'd-5415,32'd-271,32'd52,32'd10996,32'd-1489,32'd6118,32'd-4487,32'd4187,32'd-886,32'd-8105,32'd880,32'd-531,32'd5234,32'd695,32'd2819,32'd5205,32'd2985,32'd-2436,32'd3837,32'd16220,32'd6787,32'd6557,32'd3264,32'd-962,32'd4799,32'd-177,32'd12,32'd1116,32'd-1546,32'd-1894,32'd-7167,32'd5092,32'd3232,32'd-1683,32'd5917,32'd975,32'd2919,32'd7324,32'd8745,32'd-8940,32'd5253,32'd6430,32'd-1875,32'd2321,32'd-2082,32'd491,32'd-2385,32'd-4221,32'd-6293,32'd3957,32'd1241,32'd-3129,32'd3393,32'd538,32'd-7656,32'd2917,32'd-636,32'd3525,32'd-2941,32'd6313,32'd7822,32'd-806,32'd4296,32'd2534,32'd2978,32'd2188,32'd-4189,32'd6616,32'd1001,32'd3781,32'd1379,32'd4782,32'd5986,32'd1779,32'd-2927,32'd954,32'd4528,32'd6533,32'd2661,32'd2856,32'd-657,32'd-3632,32'd-1510,32'd-1618,32'd6127,32'd2900,32'd6821,32'd-19,32'd2739,32'd3,32'd-4084,32'd1043,32'd40,32'd23457,32'd-2800,32'd83,32'd5874,32'd4602,32'd-2352,32'd-3881,32'd661,32'd-1842,32'd7954,32'd2624,32'd2744,32'd-5268,32'd125,32'd135,32'd-3308,32'd2590,32'd-2218,32'd3708,32'd2792,32'd4802,32'd7719,32'd1507,32'd2565,32'd-6557,32'd-2487,32'd8183,32'd6508,32'd-1577,32'd-3942,32'd2597,32'd-8164,32'd7216,32'd167,32'd-299,32'd-2875,32'd-1396,32'd5307,32'd4458,32'd2495,32'd-6108,32'd-3286,32'd3435,32'd-5141,32'd-4389,32'd-2539,32'd323,32'd6586,32'd-2951,32'd-1318,32'd-518,32'd-3952,32'd152,32'd-4870,32'd-1253,32'd-5556,32'd4589,32'd-5839,32'd-1931,32'd1701,32'd1732,32'd-4653,32'd993,32'd-4409,32'd-7192,32'd263,32'd-2727,32'd-215,32'd-5766,32'd-2032,32'd-1238,32'd-1876,32'd3859,32'd4970,32'd-1845,32'd-9047,32'd-2763,32'd3735,32'd1286,32'd-5483,32'd-2143,32'd-4978,32'd-6669,32'd4738,32'd6259,32'd4321,32'd1745,32'd3132,32'd4431,32'd-3256,32'd2980,32'd-1467,32'd8808,32'd3442,32'd1693,32'd9169,32'd-14570,32'd91,32'd-5097,32'd-227,32'd7275,32'd-1188,32'd9135,32'd-3168,32'd-9291,32'd3183,32'd-1964,32'd-1502,32'd1194,32'd5615,32'd-210,32'd-6723,32'd-9790,32'd4326,32'd3071,32'd-4775,32'd-3547,32'd-292,32'd3447,32'd7485,32'd-3188,32'd-5708,32'd6333,32'd-1362,32'd-1214,32'd939,32'd3037,32'd8046,32'd-5073,32'd-2226,32'd8393,32'd10068,32'd-3522,32'd4121,32'd-4123,32'd957,32'd-3132,32'd544};
    Wh[2]='{32'd2076,32'd-4062,32'd574,32'd400,32'd-1826,32'd-2153,32'd-3430,32'd3229,32'd-3078,32'd2000,32'd-301,32'd-2570,32'd1149,32'd-2069,32'd-1693,32'd-75,32'd-2034,32'd-3789,32'd-3593,32'd2054,32'd780,32'd230,32'd1251,32'd1750,32'd-349,32'd180,32'd1948,32'd2442,32'd-1199,32'd-327,32'd286,32'd-2749,32'd583,32'd916,32'd-1315,32'd1612,32'd-4606,32'd-3361,32'd5244,32'd3347,32'd-958,32'd-183,32'd-3996,32'd-523,32'd-8886,32'd7250,32'd2122,32'd-1889,32'd-255,32'd-5732,32'd-1914,32'd-814,32'd-1252,32'd-6938,32'd-824,32'd-3913,32'd4694,32'd1429,32'd1293,32'd-6748,32'd3857,32'd-4360,32'd-1030,32'd-5146,32'd909,32'd-971,32'd-2858,32'd3576,32'd-2084,32'd2993,32'd-5605,32'd-3002,32'd-1196,32'd2912,32'd-1491,32'd-2110,32'd4294,32'd-2106,32'd-6835,32'd-1128,32'd1926,32'd4265,32'd-2122,32'd4931,32'd2587,32'd3303,32'd1518,32'd-217,32'd-2148,32'd-3767,32'd1611,32'd2120,32'd-2866,32'd3210,32'd2507,32'd4069,32'd-1414,32'd-289,32'd1771,32'd-857,32'd839,32'd-5561,32'd1128,32'd447,32'd-2194,32'd-318,32'd-4699,32'd-3237,32'd-15947,32'd14072,32'd-10771,32'd4978,32'd-10146,32'd-1737,32'd724,32'd2775,32'd-2751,32'd-12998,32'd7451,32'd-2407,32'd-3676,32'd-2792,32'd2958,32'd410,32'd-10195,32'd670,32'd-6977,32'd331,32'd8139,32'd-2502,32'd1380,32'd-6552,32'd4250,32'd3225,32'd-3413,32'd-5288,32'd-549,32'd-3027,32'd-2690,32'd-111,32'd5112,32'd-1602,32'd7119,32'd4921,32'd364,32'd-2524,32'd-12109,32'd767,32'd552,32'd-2070,32'd-3576,32'd-6547,32'd-2211,32'd-7070,32'd3571,32'd1822,32'd-2773,32'd1423,32'd1464,32'd-1113,32'd4265,32'd-4721,32'd2224,32'd-9404,32'd-1528,32'd-693,32'd2216,32'd-95,32'd6357,32'd-5087,32'd1243,32'd-1619,32'd-5405,32'd2922,32'd-4653,32'd-3229,32'd-3220,32'd7734,32'd-3020,32'd1101,32'd902,32'd5937,32'd3906,32'd8461,32'd5454,32'd1088,32'd-285,32'd1107,32'd9726,32'd-4746,32'd7514,32'd12324,32'd2087,32'd3239,32'd2344,32'd-11220,32'd-3640,32'd-4648,32'd-3347,32'd-3081,32'd870,32'd6025,32'd2318,32'd2531,32'd-1179,32'd1473,32'd2081,32'd1776,32'd-1034,32'd-1654,32'd5634,32'd-116,32'd259,32'd2193,32'd4267,32'd-390,32'd-5917,32'd-4565,32'd-207,32'd2529,32'd-2496,32'd171,32'd-3137,32'd-1282,32'd-2893,32'd276,32'd-1708,32'd-1356,32'd-1566,32'd3278,32'd2238,32'd-1890,32'd2932,32'd2912,32'd13623,32'd-1008,32'd1571,32'd1143,32'd4084,32'd-2897,32'd700,32'd1455,32'd-245,32'd-4340,32'd2504,32'd-5615,32'd-1632,32'd5678,32'd5229,32'd1663,32'd3422,32'd-11,32'd352,32'd783,32'd3110,32'd809,32'd2193,32'd3000,32'd-6015,32'd12490,32'd2200,32'd-5595,32'd1169,32'd4660,32'd-269,32'd3725,32'd638,32'd-3120,32'd1185,32'd127,32'd1519,32'd-2194,32'd371,32'd-473,32'd-107,32'd-1036,32'd1452,32'd4123,32'd2355,32'd5678,32'd-2929,32'd-6528,32'd3420,32'd-2988,32'd-1435,32'd4411,32'd3481,32'd2810,32'd-4611,32'd-1964,32'd-2839,32'd-217,32'd-526,32'd-1396,32'd-6313,32'd3666,32'd-1905,32'd-1966,32'd5205,32'd-629,32'd4143,32'd-4628,32'd-384,32'd-326,32'd2866,32'd3996,32'd827,32'd-2907,32'd-1705,32'd4099,32'd-1900,32'd-85,32'd3120,32'd-3007,32'd791,32'd-5874,32'd-4416,32'd-246,32'd-1850,32'd4694,32'd3618,32'd2392,32'd-2927,32'd163,32'd-1045,32'd-3498,32'd-3439,32'd4504,32'd2792,32'd3457,32'd432,32'd-1372,32'd1015,32'd509,32'd-2534,32'd2119,32'd-1789,32'd-3806,32'd-4213,32'd6967,32'd-185,32'd1243,32'd4226,32'd6264,32'd-391,32'd3237,32'd2384,32'd1629,32'd-339,32'd-3801,32'd-3576,32'd-1269,32'd7148,32'd2054,32'd-1111,32'd-957,32'd5375,32'd9335,32'd-5776,32'd-1561,32'd2673,32'd-452,32'd-1356,32'd191,32'd-1953,32'd5273,32'd-3400,32'd-5458,32'd-9116,32'd5449,32'd-303,32'd-6323,32'd-8808,32'd-2103,32'd-4726,32'd-2429,32'd-6635,32'd-1296,32'd-1213,32'd-78,32'd-2089,32'd-10156,32'd-937,32'd2519,32'd-1785,32'd6210,32'd7753,32'd-2800,32'd-1646,32'd4680,32'd-3210,32'd2249,32'd-550,32'd-4150,32'd3947,32'd-1578,32'd-5302,32'd-3251,32'd3100,32'd479};
    Wh[3]='{32'd-2863,32'd4489,32'd-1463,32'd-1452,32'd2243,32'd1173,32'd2413,32'd2163,32'd-5385,32'd585,32'd-919,32'd1712,32'd1478,32'd3156,32'd614,32'd726,32'd-1215,32'd-935,32'd3339,32'd2264,32'd729,32'd371,32'd-1062,32'd-5429,32'd-1192,32'd-2210,32'd-1134,32'd1176,32'd1079,32'd-1776,32'd2149,32'd-4062,32'd-5375,32'd-960,32'd3774,32'd906,32'd7285,32'd-60,32'd-3061,32'd6054,32'd249,32'd3125,32'd-3203,32'd-3789,32'd714,32'd2492,32'd2156,32'd-20,32'd-1174,32'd-3066,32'd-3591,32'd4257,32'd50,32'd-2008,32'd808,32'd-3415,32'd-315,32'd-5488,32'd2324,32'd-274,32'd-1921,32'd-4309,32'd1931,32'd-1641,32'd-10,32'd-528,32'd90,32'd3686,32'd2595,32'd540,32'd-1083,32'd1810,32'd1856,32'd-6093,32'd-3955,32'd6025,32'd-6010,32'd2143,32'd-466,32'd1474,32'd550,32'd1217,32'd-933,32'd-3486,32'd-3525,32'd-5312,32'd819,32'd-2224,32'd-6933,32'd-197,32'd-1782,32'd-2641,32'd1264,32'd-1551,32'd5200,32'd2415,32'd-3188,32'd4074,32'd3745,32'd2489,32'd1101,32'd496,32'd719,32'd-7426,32'd3837,32'd-463,32'd-1477,32'd-2475,32'd-3630,32'd179,32'd2526,32'd-1182,32'd-1809,32'd172,32'd660,32'd-295,32'd-657,32'd6230,32'd4934,32'd-2697,32'd-87,32'd4833,32'd-6894,32'd-2060,32'd-562,32'd704,32'd618,32'd5585,32'd501,32'd-451,32'd3208,32'd-4138,32'd302,32'd2863,32'd-6347,32'd-4045,32'd-1861,32'd-2462,32'd149,32'd964,32'd-5493,32'd3374,32'd4187,32'd3950,32'd-477,32'd-3159,32'd1309,32'd-6967,32'd4868,32'd-4953,32'd-306,32'd1200,32'd1843,32'd-5444,32'd-971,32'd-2641,32'd6064,32'd4025,32'd-1298,32'd-3237,32'd3327,32'd-1413,32'd-339,32'd-9423,32'd2753,32'd1872,32'd-755,32'd2044,32'd172,32'd610,32'd-1857,32'd5766,32'd4919,32'd-5522,32'd-1585,32'd-3518,32'd-5156,32'd172,32'd555,32'd-3305,32'd2602,32'd-1820,32'd3642,32'd43,32'd-6313,32'd-4392,32'd3908,32'd-2685,32'd-403,32'd-494,32'd1013,32'd-5610,32'd202,32'd7231,32'd1990,32'd1262,32'd2629,32'd3227,32'd-692,32'd5864,32'd2912,32'd437,32'd-3784,32'd-5073,32'd-315,32'd1662,32'd1982,32'd997,32'd1625,32'd431,32'd1120,32'd-2509,32'd1551,32'd-2126,32'd5263,32'd1296,32'd1029,32'd11982,32'd-913,32'd-3388,32'd2917,32'd-3181,32'd-3574,32'd7709,32'd-2893,32'd-3725,32'd3483,32'd2473,32'd-4133,32'd4321,32'd4243,32'd2758,32'd-455,32'd3916,32'd-2805,32'd2768,32'd-1027,32'd-449,32'd1864,32'd393,32'd-2409,32'd-447,32'd-985,32'd-4550,32'd-650,32'd1583,32'd3879,32'd2415,32'd-3891,32'd2717,32'd1172,32'd2093,32'd899,32'd3137,32'd-528,32'd3601,32'd511,32'd-3750,32'd-1177,32'd-416,32'd-2436,32'd389,32'd-753,32'd-5937,32'd1018,32'd-1385,32'd4658,32'd39,32'd-1734,32'd-1122,32'd2858,32'd3796,32'd-4626,32'd5937,32'd-4018,32'd-1396,32'd4594,32'd-925,32'd1752,32'd-1870,32'd-1494,32'd-2841,32'd-5991,32'd2646,32'd-1195,32'd-777,32'd-2780,32'd-3586,32'd6269,32'd2022,32'd2607,32'd-102,32'd-408,32'd1806,32'd1491,32'd-558,32'd5937,32'd1042,32'd3940,32'd1462,32'd1879,32'd-4226,32'd-3320,32'd-4157,32'd-1894,32'd3161,32'd814,32'd3503,32'd-4321,32'd-1168,32'd-3901,32'd-2961,32'd960,32'd-3183,32'd799,32'd4343,32'd-4645,32'd2690,32'd-1110,32'd1885,32'd2604,32'd-2700,32'd-2536,32'd-3977,32'd-7285,32'd-2147,32'd-805,32'd1851,32'd-2878,32'd1910,32'd-2583,32'd-1851,32'd1205,32'd-1995,32'd680,32'd-2746,32'd-1552,32'd6040,32'd-167,32'd-1,32'd-1101,32'd2380,32'd684,32'd565,32'd1539,32'd3723,32'd1718,32'd3203,32'd3779,32'd-944,32'd859,32'd4316,32'd-150,32'd-2897,32'd2435,32'd913,32'd-3552,32'd-6660,32'd2122,32'd41,32'd2065,32'd-5805,32'd451,32'd-3188,32'd981,32'd-2108,32'd2756,32'd631,32'd4787,32'd-2731,32'd-1066,32'd1779,32'd2878,32'd2956,32'd1614,32'd-255,32'd-2663,32'd-628,32'd1490,32'd-618,32'd-530,32'd-1520,32'd-3569,32'd-6357,32'd1520,32'd-5585,32'd2156,32'd-469,32'd-3886,32'd-4216,32'd5185,32'd-2329,32'd-5190,32'd6298,32'd1268,32'd-1325,32'd6601,32'd2758,32'd-2780,32'd-509};
    Wh[4]='{32'd-845,32'd2348,32'd-3120,32'd-3098,32'd-796,32'd-265,32'd1809,32'd1276,32'd32,32'd-2117,32'd-1944,32'd1028,32'd-1264,32'd2109,32'd-5312,32'd-2032,32'd-6132,32'd-3283,32'd-1325,32'd410,32'd1817,32'd-1213,32'd2203,32'd989,32'd-1770,32'd299,32'd1112,32'd1821,32'd158,32'd-2263,32'd-436,32'd2177,32'd-92,32'd1652,32'd3085,32'd-1467,32'd3349,32'd-1282,32'd2871,32'd-1693,32'd-2437,32'd-2597,32'd2199,32'd-2751,32'd1372,32'd-2673,32'd-2274,32'd-1606,32'd-2475,32'd-202,32'd1110,32'd-2188,32'd3227,32'd2761,32'd-152,32'd-7446,32'd80,32'd-1469,32'd2321,32'd-3012,32'd1362,32'd-428,32'd1070,32'd-3327,32'd-2990,32'd508,32'd2253,32'd-1264,32'd-301,32'd-873,32'd1805,32'd-587,32'd-148,32'd1467,32'd-1380,32'd-2186,32'd-1351,32'd-33,32'd2521,32'd-277,32'd-2264,32'd4233,32'd-1239,32'd-1861,32'd-1063,32'd-1347,32'd-1108,32'd486,32'd668,32'd-1835,32'd-2480,32'd-5263,32'd-1512,32'd-2646,32'd-931,32'd-402,32'd-503,32'd270,32'd1330,32'd-1054,32'd-2062,32'd-853,32'd-1899,32'd5249,32'd-1600,32'd-1047,32'd-91,32'd25,32'd-1984,32'd2590,32'd-564,32'd-6337,32'd-6459,32'd1206,32'd-3039,32'd-2495,32'd181,32'd-693,32'd-21,32'd3161,32'd169,32'd-2878,32'd-3220,32'd-6440,32'd881,32'd2049,32'd422,32'd-1213,32'd2418,32'd5244,32'd-4941,32'd-2156,32'd-390,32'd-3598,32'd957,32'd1026,32'd-1781,32'd2006,32'd-859,32'd3071,32'd4938,32'd-2700,32'd4851,32'd1289,32'd986,32'd4711,32'd1951,32'd2437,32'd-306,32'd-1984,32'd653,32'd5556,32'd197,32'd472,32'd-84,32'd8959,32'd-2534,32'd-2731,32'd-680,32'd-3420,32'd-3234,32'd2368,32'd1732,32'd-3254,32'd1086,32'd-722,32'd-560,32'd-5024,32'd-2161,32'd-1401,32'd-3186,32'd-6718,32'd845,32'd2420,32'd2347,32'd564,32'd-2209,32'd3054,32'd-1064,32'd-873,32'd2092,32'd-1391,32'd-3378,32'd521,32'd513,32'd1663,32'd1719,32'd-569,32'd-207,32'd522,32'd761,32'd-3579,32'd3420,32'd4169,32'd-1833,32'd-5034,32'd1523,32'd-2094,32'd3161,32'd-2221,32'd1920,32'd5708,32'd-25,32'd5146,32'd-1652,32'd2851,32'd856,32'd1518,32'd-3020,32'd709,32'd-2235,32'd1893,32'd-842,32'd83,32'd2868,32'd-6245,32'd-985,32'd-1685,32'd206,32'd2043,32'd-1682,32'd-6030,32'd-2122,32'd-1823,32'd-3481,32'd-502,32'd-4006,32'd1047,32'd2393,32'd3225,32'd-115,32'd8789,32'd-350,32'd1033,32'd-4069,32'd2561,32'd-897,32'd2133,32'd79,32'd6118,32'd-3698,32'd3410,32'd933,32'd4748,32'd-874,32'd2027,32'd-2556,32'd544,32'd-2237,32'd487,32'd1545,32'd142,32'd-191,32'd-3081,32'd-969,32'd422,32'd2004,32'd-314,32'd-168,32'd-834,32'd-533,32'd-2213,32'd-1940,32'd1071,32'd1452,32'd-2121,32'd-750,32'd-1348,32'd-1232,32'd50,32'd727,32'd2578,32'd-443,32'd-1979,32'd-128,32'd-2027,32'd676,32'd593,32'd-3493,32'd-578,32'd-1726,32'd-221,32'd-3186,32'd4475,32'd-1446,32'd147,32'd1227,32'd126,32'd-1480,32'd-1556,32'd-3657,32'd-611,32'd1278,32'd-1196,32'd-1282,32'd2144,32'd-1068,32'd-5048,32'd-2423,32'd-1052,32'd351,32'd-65,32'd161,32'd3024,32'd-578,32'd-2519,32'd-4182,32'd3669,32'd-567,32'd-604,32'd-1417,32'd-1120,32'd-4382,32'd-2379,32'd-1093,32'd-783,32'd-15,32'd-1790,32'd-2685,32'd-1582,32'd-4272,32'd-6181,32'd-962,32'd2954,32'd-1596,32'd2022,32'd-1578,32'd280,32'd-1006,32'd1278,32'd-4499,32'd-823,32'd4365,32'd1953,32'd-680,32'd-1997,32'd1378,32'd-2941,32'd665,32'd-163,32'd-3940,32'd-1064,32'd-223,32'd1146,32'd3068,32'd2980,32'd1453,32'd-4685,32'd-2188,32'd1284,32'd-2702,32'd541,32'd1656,32'd-2556,32'd379,32'd-1463,32'd-2231,32'd-2186,32'd-2377,32'd-3161,32'd-943,32'd-2266,32'd3811,32'd356,32'd2504,32'd-5571,32'd-2409,32'd6459,32'd-4858,32'd-8115,32'd2155,32'd1982,32'd-4650,32'd-2307,32'd-2160,32'd-1146,32'd-1757,32'd-1091,32'd1441,32'd1867,32'd-937,32'd-34,32'd-2836,32'd1843,32'd-2592,32'd-2371,32'd1280,32'd272,32'd-2437,32'd-4091,32'd-1890,32'd1322,32'd-1446,32'd3029,32'd1613,32'd-333,32'd1865,32'd3823,32'd-3237,32'd-3271};
    Wh[5]='{32'd-1496,32'd6523,32'd3295,32'd-1099,32'd-497,32'd-552,32'd-7524,32'd-4521,32'd-1317,32'd671,32'd-3007,32'd-98,32'd-4887,32'd-3542,32'd2086,32'd-1333,32'd1965,32'd-511,32'd-1333,32'd-1536,32'd629,32'd79,32'd-1770,32'd-2854,32'd-1033,32'd-1541,32'd-1412,32'd-1400,32'd-2486,32'd1240,32'd-1680,32'd-5732,32'd2287,32'd1066,32'd-506,32'd762,32'd517,32'd2135,32'd-2117,32'd4611,32'd-34,32'd-426,32'd-2205,32'd-2685,32'd-6367,32'd458,32'd-5869,32'd-1269,32'd2819,32'd-2500,32'd-2409,32'd5122,32'd-483,32'd-1711,32'd-3364,32'd-3833,32'd2312,32'd-2189,32'd2995,32'd722,32'd-2968,32'd424,32'd-3098,32'd3181,32'd585,32'd-1759,32'd-1159,32'd-2661,32'd-747,32'd-2595,32'd-3784,32'd-2235,32'd2807,32'd-792,32'd3723,32'd-3471,32'd-1575,32'd-3789,32'd-2238,32'd547,32'd2270,32'd1563,32'd-5175,32'd6484,32'd328,32'd613,32'd1616,32'd3581,32'd-1192,32'd-3466,32'd-7,32'd-133,32'd-322,32'd-356,32'd-5781,32'd-2141,32'd-530,32'd3273,32'd-2049,32'd2570,32'd-833,32'd-557,32'd363,32'd-7373,32'd-897,32'd1776,32'd-3041,32'd-3908,32'd-4865,32'd2423,32'd1387,32'd384,32'd-236,32'd-1203,32'd5014,32'd3835,32'd733,32'd-2260,32'd751,32'd-122,32'd-1301,32'd-5302,32'd6049,32'd9233,32'd-1252,32'd-4294,32'd2224,32'd1323,32'd-4956,32'd-14326,32'd3034,32'd1016,32'd436,32'd-3383,32'd-3212,32'd1824,32'd-1143,32'd-396,32'd2421,32'd-968,32'd1563,32'd2612,32'd3369,32'd-1801,32'd-225,32'd2252,32'd-5747,32'd-5590,32'd-3220,32'd-3137,32'd-5380,32'd-6191,32'd-3713,32'd3627,32'd231,32'd-1185,32'd-1701,32'd2531,32'd2213,32'd8129,32'd411,32'd-5546,32'd-1335,32'd5268,32'd-414,32'd-1440,32'd2207,32'd2807,32'd367,32'd-3903,32'd2279,32'd13906,32'd-361,32'd4653,32'd2880,32'd-185,32'd5639,32'd-2744,32'd1417,32'd1033,32'd-3378,32'd-8159,32'd499,32'd-2215,32'd-2988,32'd3957,32'd-1358,32'd4829,32'd7768,32'd-346,32'd2022,32'd658,32'd8613,32'd-931,32'd-3198,32'd-9189,32'd879,32'd2103,32'd-4885,32'd-3247,32'd-1286,32'd-2067,32'd-885,32'd-1895,32'd-4763,32'd-258,32'd-995,32'd1149,32'd3598,32'd2121,32'd3286,32'd906,32'd3752,32'd5087,32'd-1171,32'd2661,32'd-3085,32'd294,32'd2374,32'd-6357,32'd983,32'd-411,32'd2124,32'd3198,32'd1174,32'd1928,32'd3161,32'd-3947,32'd440,32'd329,32'd3051,32'd-877,32'd1337,32'd2371,32'd1975,32'd643,32'd3913,32'd1394,32'd9033,32'd-480,32'd4755,32'd-7548,32'd550,32'd878,32'd2648,32'd991,32'd3010,32'd-300,32'd1353,32'd3225,32'd6123,32'd1262,32'd-3400,32'd1334,32'd2517,32'd-4531,32'd892,32'd592,32'd38,32'd50,32'd2502,32'd486,32'd3464,32'd1341,32'd1708,32'd-419,32'd-877,32'd2247,32'd-736,32'd1276,32'd5571,32'd-2780,32'd4760,32'd590,32'd1748,32'd-1916,32'd4560,32'd-2403,32'd2575,32'd1538,32'd3901,32'd-1569,32'd-1845,32'd1398,32'd-2203,32'd-796,32'd-1944,32'd697,32'd770,32'd3752,32'd-369,32'd7548,32'd-199,32'd-3679,32'd559,32'd2038,32'd1604,32'd-4272,32'd6621,32'd-2442,32'd-1770,32'd-366,32'd1364,32'd5102,32'd-293,32'd2783,32'd1007,32'd-4870,32'd-567,32'd2900,32'd587,32'd46,32'd-1467,32'd6640,32'd1479,32'd-6528,32'd-2985,32'd1148,32'd3239,32'd-2399,32'd4797,32'd1937,32'd2797,32'd-1700,32'd-2059,32'd1129,32'd4582,32'd-1779,32'd-1627,32'd-223,32'd5068,32'd1835,32'd-361,32'd713,32'd-3828,32'd5869,32'd-1240,32'd4448,32'd-278,32'd1262,32'd5922,32'd-4775,32'd-808,32'd-1004,32'd-2147,32'd-755,32'd-6259,32'd3864,32'd9843,32'd-1995,32'd-4201,32'd1453,32'd2795,32'd582,32'd1201,32'd-6372,32'd3891,32'd11113,32'd3544,32'd-2875,32'd-3027,32'd664,32'd2227,32'd4997,32'd-2578,32'd1035,32'd-1115,32'd-6596,32'd-1480,32'd2092,32'd-1391,32'd-3305,32'd4985,32'd3098,32'd3320,32'd-3154,32'd-812,32'd-1943,32'd-592,32'd671,32'd-664,32'd-1098,32'd-4482,32'd-1182,32'd2271,32'd916,32'd-1605,32'd360,32'd2318,32'd2454,32'd-8388,32'd-6059,32'd4174,32'd-6289,32'd144,32'd-481,32'd-10595,32'd-4045,32'd1076,32'd181};
    Wh[6]='{32'd-2973,32'd526,32'd1638,32'd1927,32'd-1418,32'd-1130,32'd-357,32'd-3164,32'd511,32'd-684,32'd-1735,32'd-3750,32'd-610,32'd-4489,32'd-1026,32'd-7114,32'd657,32'd9306,32'd694,32'd704,32'd-1702,32'd-433,32'd2352,32'd-2407,32'd-1657,32'd1783,32'd5292,32'd-159,32'd643,32'd6015,32'd3244,32'd6699,32'd-6552,32'd-1015,32'd-9833,32'd883,32'd-7226,32'd-3088,32'd-4406,32'd4794,32'd-2744,32'd-1961,32'd1739,32'd1693,32'd-2985,32'd-1250,32'd3083,32'd-2227,32'd-2512,32'd1108,32'd-2573,32'd1838,32'd8715,32'd366,32'd5317,32'd-5297,32'd2464,32'd-4855,32'd-1472,32'd-2622,32'd-1916,32'd2919,32'd-1750,32'd-2568,32'd-1666,32'd783,32'd1088,32'd1409,32'd1278,32'd2937,32'd-3869,32'd-320,32'd4233,32'd1367,32'd-6904,32'd993,32'd822,32'd1363,32'd-7246,32'd1126,32'd-1406,32'd-7500,32'd-1363,32'd10283,32'd322,32'd-3608,32'd-558,32'd3022,32'd10,32'd-5708,32'd-1883,32'd-1676,32'd8232,32'd3813,32'd5092,32'd-428,32'd1054,32'd2998,32'd4438,32'd-1947,32'd-2341,32'd2093,32'd1610,32'd15673,32'd3349,32'd828,32'd2360,32'd13623,32'd2335,32'd7294,32'd4111,32'd-6000,32'd12080,32'd-3637,32'd-581,32'd-5249,32'd-2695,32'd4973,32'd2851,32'd886,32'd-3078,32'd-11044,32'd751,32'd3146,32'd3984,32'd-2534,32'd3071,32'd6289,32'd2844,32'd-6665,32'd269,32'd467,32'd-1798,32'd-4865,32'd-6049,32'd5712,32'd-2106,32'd-7255,32'd-2396,32'd-1308,32'd-429,32'd9399,32'd6215,32'd-2351,32'd-1004,32'd-2493,32'd-2131,32'd-1787,32'd1043,32'd-1245,32'd2399,32'd-2495,32'd2265,32'd3715,32'd-1148,32'd-3249,32'd-10507,32'd2968,32'd2365,32'd-3266,32'd-1622,32'd3967,32'd-4533,32'd401,32'd-1711,32'd-3376,32'd2915,32'd-502,32'd576,32'd1019,32'd-8828,32'd-1192,32'd353,32'd3510,32'd-11103,32'd1051,32'd-358,32'd-2958,32'd718,32'd-2990,32'd2937,32'd-820,32'd17031,32'd2673,32'd1748,32'd2788,32'd4213,32'd4753,32'd1604,32'd-3264,32'd4724,32'd-1973,32'd-789,32'd-3605,32'd3647,32'd1557,32'd-5332,32'd-4892,32'd9238,32'd-3969,32'd-1579,32'd-1239,32'd1425,32'd2988,32'd-1210,32'd-220,32'd55,32'd5869,32'd4689,32'd-4047,32'd1105,32'd8378,32'd1535,32'd-516,32'd-1845,32'd7304,32'd3847,32'd-1804,32'd1564,32'd-1728,32'd-2487,32'd8950,32'd8662,32'd-3125,32'd-426,32'd3642,32'd4836,32'd-1107,32'd-5366,32'd-1650,32'd-2137,32'd2053,32'd1602,32'd214,32'd6479,32'd2358,32'd1851,32'd2014,32'd8989,32'd-3674,32'd448,32'd-4509,32'd2651,32'd4094,32'd5947,32'd-4138,32'd-3342,32'd-2949,32'd10498,32'd1827,32'd2854,32'd-2846,32'd-1004,32'd-1564,32'd361,32'd5498,32'd2788,32'd-4262,32'd-3002,32'd-3200,32'd-3115,32'd5009,32'd-4240,32'd7714,32'd6284,32'd1292,32'd-3815,32'd2017,32'd-1571,32'd-3098,32'd724,32'd2995,32'd-100,32'd-2849,32'd-3808,32'd-1231,32'd5903,32'd2561,32'd-24,32'd4423,32'd4006,32'd316,32'd-6054,32'd-1428,32'd4738,32'd22,32'd1425,32'd49,32'd-584,32'd2082,32'd-4855,32'd-4912,32'd480,32'd4799,32'd5107,32'd7856,32'd4182,32'd-696,32'd5439,32'd1032,32'd1363,32'd-8930,32'd767,32'd-341,32'd-1790,32'd5947,32'd6738,32'd4826,32'd-953,32'd-4108,32'd2565,32'd-453,32'd10791,32'd1965,32'd-10371,32'd-3371,32'd6098,32'd-5478,32'd3339,32'd2198,32'd1385,32'd8798,32'd2396,32'd-433,32'd-905,32'd6958,32'd9311,32'd3400,32'd4843,32'd3605,32'd-2054,32'd2106,32'd756,32'd-3608,32'd3010,32'd13593,32'd1700,32'd-1156,32'd-6757,32'd3359,32'd-1246,32'd6274,32'd960,32'd3100,32'd-6069,32'd-385,32'd-616,32'd-967,32'd-1741,32'd2946,32'd2365,32'd3789,32'd-1735,32'd4638,32'd952,32'd-4729,32'd4497,32'd-12167,32'd-14443,32'd1034,32'd445,32'd2432,32'd-777,32'd-3872,32'd-7309,32'd196,32'd4252,32'd1616,32'd-3144,32'd989,32'd3940,32'd3525,32'd5444,32'd-8442,32'd3168,32'd-272,32'd903,32'd-2595,32'd-466,32'd445,32'd3435,32'd-1287,32'd6049,32'd3532,32'd-443,32'd-2966,32'd736,32'd-2148,32'd782,32'd-5273,32'd-8681,32'd4619,32'd-588,32'd574,32'd2622,32'd-720,32'd739,32'd-1091,32'd5747,32'd-49};
    Wh[7]='{32'd-858,32'd49,32'd-1000,32'd2321,32'd-608,32'd2902,32'd-1904,32'd7509,32'd-1369,32'd3471,32'd6845,32'd-1602,32'd-5854,32'd4899,32'd-8461,32'd-5800,32'd3203,32'd-1925,32'd-4484,32'd-147,32'd-831,32'd4541,32'd-242,32'd-2177,32'd-1552,32'd2222,32'd-1190,32'd1053,32'd1226,32'd-1650,32'd-3840,32'd6313,32'd-1467,32'd-3017,32'd-4306,32'd2556,32'd-7397,32'd-4199,32'd-233,32'd8774,32'd-2390,32'd-3874,32'd-2580,32'd3845,32'd-6181,32'd-9399,32'd-5590,32'd744,32'd2946,32'd-4814,32'd6347,32'd-1979,32'd3220,32'd-4460,32'd-4804,32'd-835,32'd-1627,32'd7695,32'd-1036,32'd3786,32'd3527,32'd2434,32'd-1862,32'd-5512,32'd-8881,32'd2462,32'd-2673,32'd5825,32'd563,32'd2073,32'd1407,32'd7143,32'd-2565,32'd-1152,32'd-8969,32'd-2143,32'd8833,32'd-1593,32'd-1644,32'd-2302,32'd-1076,32'd2260,32'd-6860,32'd2995,32'd2269,32'd1507,32'd-3002,32'd1545,32'd1840,32'd2283,32'd-3291,32'd-4777,32'd-578,32'd9125,32'd4277,32'd-617,32'd-6879,32'd-1574,32'd5434,32'd1397,32'd3916,32'd-1004,32'd3535,32'd3974,32'd-2467,32'd-1879,32'd-6743,32'd-4826,32'd5737,32'd-2454,32'd5800,32'd774,32'd9658,32'd-2944,32'd-3361,32'd-473,32'd-3898,32'd20488,32'd3137,32'd-4655,32'd-1315,32'd-7602,32'd-4245,32'd2568,32'd6088,32'd-8525,32'd3491,32'd2009,32'd2258,32'd3459,32'd13535,32'd-2749,32'd1303,32'd1199,32'd-8847,32'd-2352,32'd-1835,32'd-720,32'd1145,32'd-1712,32'd11777,32'd5942,32'd12353,32'd-9863,32'd2758,32'd-3913,32'd-6352,32'd-2431,32'd-2661,32'd1188,32'd2814,32'd2636,32'd-3786,32'd-1710,32'd8920,32'd-585,32'd-17412,32'd1365,32'd2324,32'd-8852,32'd21425,32'd4692,32'd2680,32'd6469,32'd-1462,32'd-12636,32'd3295,32'd2014,32'd2695,32'd-3520,32'd1721,32'd-1667,32'd-572,32'd-2410,32'd-5107,32'd-3674,32'd-3481,32'd-4274,32'd2800,32'd3117,32'd2185,32'd2271,32'd2714,32'd-1556,32'd5844,32'd192,32'd777,32'd8266,32'd4992,32'd-5434,32'd7182,32'd1022,32'd1162,32'd1534,32'd1195,32'd386,32'd835,32'd3181,32'd479,32'd-1579,32'd3046,32'd8208,32'd-1738,32'd13281,32'd4572,32'd640,32'd2225,32'd12177,32'd5058,32'd-366,32'd2888,32'd3537,32'd8779,32'd9184,32'd4997,32'd8251,32'd-473,32'd-8251,32'd-1154,32'd8173,32'd1237,32'd-2687,32'd7207,32'd862,32'd3366,32'd3269,32'd1441,32'd1926,32'd-2039,32'd6235,32'd2763,32'd7675,32'd-972,32'd4104,32'd1639,32'd-1127,32'd6582,32'd-2639,32'd6293,32'd-591,32'd344,32'd202,32'd-2478,32'd5185,32'd4042,32'd-1361,32'd-2443,32'd1575,32'd2460,32'd-631,32'd-2095,32'd-2539,32'd1866,32'd778,32'd382,32'd4460,32'd-2445,32'd1403,32'd-674,32'd2641,32'd3627,32'd2895,32'd240,32'd-1741,32'd6538,32'd1367,32'd2016,32'd1062,32'd-2277,32'd1802,32'd2915,32'd10312,32'd-2758,32'd3195,32'd1297,32'd6606,32'd3908,32'd1688,32'd1932,32'd-1483,32'd6054,32'd-702,32'd-2320,32'd-2259,32'd-2744,32'd1292,32'd519,32'd3220,32'd-1855,32'd2758,32'd-910,32'd-1933,32'd6049,32'd93,32'd-2153,32'd-2072,32'd-3723,32'd2412,32'd-348,32'd-1139,32'd-521,32'd-1397,32'd-3715,32'd1314,32'd-2612,32'd4414,32'd2139,32'd3088,32'd1478,32'd-3911,32'd671,32'd4802,32'd11601,32'd-5942,32'd-5917,32'd-1514,32'd1738,32'd1412,32'd-3283,32'd-2924,32'd-1406,32'd3483,32'd4375,32'd2695,32'd-982,32'd3615,32'd-3520,32'd3798,32'd2790,32'd2968,32'd-2756,32'd2493,32'd6782,32'd7470,32'd587,32'd4055,32'd587,32'd-2707,32'd-1901,32'd10263,32'd-4028,32'd2380,32'd-1851,32'd-631,32'd-1826,32'd1843,32'd-5664,32'd3496,32'd7680,32'd7514,32'd-114,32'd-2042,32'd2790,32'd4206,32'd-4223,32'd-6123,32'd482,32'd2990,32'd-5312,32'd3168,32'd4455,32'd358,32'd-1918,32'd1784,32'd1727,32'd4,32'd170,32'd4384,32'd2302,32'd3276,32'd-31,32'd6645,32'd1183,32'd-469,32'd-7524,32'd20,32'd-3535,32'd-1358,32'd-3352,32'd7080,32'd4736,32'd-1160,32'd-292,32'd3530,32'd2080,32'd-2722,32'd-1006,32'd6591,32'd-2636,32'd-4243,32'd-1617,32'd2479,32'd-1433,32'd3308,32'd-2553,32'd-4763,32'd-6372,32'd-3696,32'd-429,32'd5722};
    Wh[8]='{32'd-1418,32'd-455,32'd-2354,32'd-2661,32'd-2048,32'd2297,32'd-7587,32'd-2739,32'd2299,32'd2812,32'd2232,32'd-1697,32'd-3894,32'd984,32'd-852,32'd3415,32'd36,32'd1875,32'd-921,32'd-218,32'd-32,32'd1889,32'd4614,32'd2407,32'd-1918,32'd2873,32'd-3898,32'd-1702,32'd-2221,32'd706,32'd159,32'd1336,32'd-1063,32'd527,32'd-247,32'd-2312,32'd610,32'd-397,32'd3364,32'd2590,32'd625,32'd-2861,32'd-2692,32'd501,32'd-3676,32'd530,32'd156,32'd-507,32'd-919,32'd3837,32'd-2235,32'd-6567,32'd-3615,32'd-4089,32'd-1954,32'd-4472,32'd87,32'd-1148,32'd2971,32'd-1502,32'd-2744,32'd269,32'd-1849,32'd-3337,32'd-6108,32'd-6098,32'd-333,32'd-1183,32'd4577,32'd-550,32'd121,32'd2756,32'd759,32'd-4428,32'd-1925,32'd4079,32'd-4262,32'd1348,32'd-2197,32'd-1614,32'd160,32'd962,32'd-2663,32'd1140,32'd-1130,32'd270,32'd1188,32'd-5063,32'd-5830,32'd-2829,32'd-1012,32'd5449,32'd-939,32'd216,32'd616,32'd-3222,32'd1431,32'd-2261,32'd2474,32'd-1829,32'd2932,32'd-2939,32'd1682,32'd-1541,32'd5454,32'd24,32'd-1652,32'd-2457,32'd125,32'd939,32'd2321,32'd-3979,32'd-2395,32'd-2644,32'd-1494,32'd204,32'd3449,32'd3896,32'd2028,32'd-2358,32'd408,32'd2084,32'd-1252,32'd-2578,32'd-8676,32'd-7744,32'd1861,32'd3203,32'd-1717,32'd1800,32'd-4206,32'd2910,32'd-2192,32'd-2675,32'd481,32'd1744,32'd3513,32'd-1403,32'd2008,32'd331,32'd3925,32'd-1203,32'd4433,32'd-2509,32'd-5341,32'd2083,32'd914,32'd246,32'd1494,32'd-3125,32'd-1047,32'd2661,32'd-984,32'd6938,32'd-6113,32'd7968,32'd924,32'd4162,32'd-7011,32'd-2695,32'd-4624,32'd-1268,32'd-4733,32'd1124,32'd3198,32'd-1394,32'd-1771,32'd3620,32'd1450,32'd547,32'd-6127,32'd-1146,32'd-2084,32'd169,32'd-1094,32'd-611,32'd259,32'd2678,32'd1413,32'd110,32'd623,32'd-2471,32'd2303,32'd-1123,32'd90,32'd1193,32'd63,32'd-1290,32'd2227,32'd-3244,32'd-6967,32'd1133,32'd2585,32'd2420,32'd-6625,32'd6484,32'd2076,32'd-3337,32'd2246,32'd4836,32'd-615,32'd-718,32'd-2178,32'd1768,32'd-317,32'd1038,32'd-1315,32'd1227,32'd96,32'd-578,32'd-4516,32'd120,32'd3935,32'd197,32'd-1660,32'd-3134,32'd-3330,32'd466,32'd-5009,32'd-6040,32'd-1893,32'd3842,32'd-4726,32'd-1776,32'd-1246,32'd-4516,32'd706,32'd-3461,32'd2111,32'd1358,32'd-1959,32'd139,32'd-4768,32'd4631,32'd-329,32'd-1732,32'd852,32'd-1418,32'd3469,32'd-4785,32'd-3215,32'd2089,32'd2678,32'd-3024,32'd-1181,32'd418,32'd850,32'd-1765,32'd-2198,32'd597,32'd-3830,32'd-2785,32'd193,32'd-3063,32'd-4062,32'd-1401,32'd-2320,32'd-3193,32'd1546,32'd653,32'd-2729,32'd-7705,32'd-3554,32'd-5180,32'd-2917,32'd-5307,32'd1185,32'd389,32'd-414,32'd800,32'd-5698,32'd5273,32'd-4355,32'd-248,32'd1657,32'd-523,32'd3601,32'd-1218,32'd2268,32'd267,32'd-4514,32'd2205,32'd-2197,32'd189,32'd-520,32'd2797,32'd349,32'd808,32'd-356,32'd5,32'd3056,32'd6020,32'd691,32'd3171,32'd1207,32'd-1745,32'd2091,32'd-3730,32'd-4875,32'd2685,32'd-293,32'd-3432,32'd-2541,32'd231,32'd-2197,32'd694,32'd-4541,32'd-1865,32'd-427,32'd-6689,32'd6928,32'd-1730,32'd-3842,32'd-4125,32'd418,32'd803,32'd-708,32'd2194,32'd-4245,32'd-5581,32'd-1138,32'd-3261,32'd-967,32'd640,32'd-1174,32'd-1397,32'd-1428,32'd-3330,32'd-6630,32'd1708,32'd-1613,32'd3342,32'd4440,32'd-1669,32'd7485,32'd186,32'd-267,32'd-3803,32'd2187,32'd3283,32'd-3598,32'd2116,32'd2133,32'd-1743,32'd-2391,32'd4716,32'd3654,32'd327,32'd5170,32'd200,32'd3264,32'd-1102,32'd5102,32'd968,32'd2744,32'd1723,32'd-105,32'd-6469,32'd-3327,32'd-3310,32'd-4907,32'd-1917,32'd1789,32'd-3342,32'd-4362,32'd3916,32'd-3107,32'd4060,32'd-1208,32'd701,32'd-5590,32'd5278,32'd-5932,32'd-4992,32'd-5175,32'd-228,32'd-562,32'd-2242,32'd-2641,32'd-2115,32'd-5327,32'd-4841,32'd-4885,32'd-2169,32'd-117,32'd-2457,32'd2244,32'd-913,32'd-6542,32'd655,32'd-740,32'd2241,32'd-6010,32'd-2727,32'd-2687,32'd-2233,32'd-323,32'd-2248,32'd-1750,32'd1829};
    Wh[9]='{32'd-3085,32'd4235,32'd1091,32'd-458,32'd3920,32'd-1107,32'd249,32'd-1989,32'd3657,32'd-1075,32'd4736,32'd216,32'd710,32'd2006,32'd6938,32'd1749,32'd4296,32'd3842,32'd-834,32'd-308,32'd1551,32'd864,32'd-2213,32'd2208,32'd873,32'd-1679,32'd997,32'd-379,32'd3415,32'd3054,32'd1896,32'd1511,32'd2335,32'd2174,32'd1072,32'd2631,32'd-226,32'd2447,32'd1368,32'd-3098,32'd-68,32'd-3161,32'd-4321,32'd3457,32'd-2019,32'd4218,32'd3979,32'd4753,32'd-87,32'd199,32'd-761,32'd-403,32'd2612,32'd3513,32'd1284,32'd5395,32'd186,32'd-108,32'd1798,32'd1026,32'd-1724,32'd4172,32'd3925,32'd-1024,32'd1729,32'd-1144,32'd-1192,32'd6826,32'd1873,32'd-2294,32'd1861,32'd1561,32'd1015,32'd705,32'd2469,32'd4033,32'd3569,32'd2749,32'd-3059,32'd-1238,32'd-105,32'd5966,32'd-764,32'd1397,32'd-3725,32'd888,32'd524,32'd3510,32'd5937,32'd-1826,32'd-387,32'd4733,32'd3825,32'd842,32'd-1220,32'd-447,32'd3464,32'd-1064,32'd3432,32'd5551,32'd1110,32'd-2346,32'd-193,32'd1661,32'd4694,32'd198,32'd5449,32'd3193,32'd-5454,32'd1342,32'd273,32'd-2885,32'd2241,32'd5351,32'd1253,32'd-370,32'd4218,32'd-5917,32'd3469,32'd1340,32'd-1677,32'd991,32'd-3796,32'd4204,32'd-1062,32'd-439,32'd3093,32'd290,32'd-4855,32'd-6367,32'd4028,32'd430,32'd2416,32'd2115,32'd2054,32'd-1190,32'd-3666,32'd2648,32'd-396,32'd-2629,32'd-7495,32'd-3781,32'd640,32'd-2851,32'd-4846,32'd3745,32'd-2575,32'd1594,32'd2770,32'd-1014,32'd-4382,32'd-665,32'd-1280,32'd296,32'd-3112,32'd-3940,32'd469,32'd627,32'd-1510,32'd5175,32'd-670,32'd3117,32'd229,32'd1192,32'd4057,32'd2778,32'd4089,32'd-4,32'd-741,32'd-1155,32'd8203,32'd5966,32'd-2279,32'd-2788,32'd-3620,32'd-1518,32'd1267,32'd137,32'd4912,32'd742,32'd-463,32'd1906,32'd6391,32'd-3596,32'd-39,32'd-2052,32'd-339,32'd-393,32'd-7827,32'd-2456,32'd789,32'd-560,32'd413,32'd3198,32'd4357,32'd91,32'd1289,32'd880,32'd-1362,32'd-3823,32'd2342,32'd-328,32'd-3757,32'd3127,32'd1745,32'd-772,32'd-796,32'd401,32'd5771,32'd4743,32'd20,32'd-1733,32'd-6171,32'd-4067,32'd-4313,32'd-3605,32'd-1267,32'd3176,32'd-63,32'd-659,32'd-189,32'd4675,32'd1844,32'd-233,32'd81,32'd1759,32'd4599,32'd-381,32'd-2734,32'd4140,32'd828,32'd786,32'd4182,32'd-336,32'd5585,32'd1223,32'd3872,32'd725,32'd-1185,32'd940,32'd-1295,32'd-6435,32'd158,32'd-508,32'd-1398,32'd-4663,32'd-1495,32'd-1684,32'd-1997,32'd4816,32'd-1141,32'd-968,32'd1212,32'd-2861,32'd1938,32'd2293,32'd-5278,32'd-3312,32'd-925,32'd-3894,32'd-885,32'd758,32'd-5000,32'd3332,32'd-774,32'd-1723,32'd-1632,32'd-5063,32'd877,32'd-2722,32'd1712,32'd-3110,32'd4130,32'd-4880,32'd-722,32'd-3476,32'd-812,32'd3410,32'd1213,32'd2917,32'd1992,32'd2893,32'd-2839,32'd-5107,32'd-14,32'd2019,32'd-1273,32'd-1041,32'd-3383,32'd-1407,32'd7973,32'd834,32'd-235,32'd56,32'd-892,32'd-1386,32'd1062,32'd-286,32'd-58,32'd2963,32'd210,32'd1228,32'd-4672,32'd406,32'd451,32'd5820,32'd4392,32'd-3632,32'd1942,32'd1082,32'd2202,32'd-2056,32'd-1072,32'd5664,32'd-3034,32'd-249,32'd4609,32'd1605,32'd1545,32'd910,32'd7734,32'd3503,32'd956,32'd-1256,32'd3701,32'd-721,32'd2614,32'd334,32'd-2330,32'd1397,32'd6298,32'd-2897,32'd-4562,32'd905,32'd-3574,32'd4111,32'd2008,32'd6684,32'd3371,32'd-5004,32'd296,32'd-1167,32'd-491,32'd620,32'd-1914,32'd3891,32'd944,32'd1993,32'd10000,32'd-1166,32'd275,32'd794,32'd147,32'd2587,32'd3337,32'd-5771,32'd2788,32'd1948,32'd-2561,32'd4775,32'd-1273,32'd2296,32'd-346,32'd11,32'd1296,32'd-4833,32'd-2597,32'd-5991,32'd-1215,32'd1889,32'd917,32'd-2451,32'd6245,32'd1204,32'd5478,32'd-162,32'd-2215,32'd127,32'd1900,32'd2003,32'd5600,32'd-1983,32'd-1256,32'd-3122,32'd-1643,32'd2142,32'd495,32'd564,32'd-1824,32'd2298,32'd3161,32'd-2000,32'd914,32'd3039,32'd-1900,32'd3974,32'd7998,32'd839,32'd908,32'd4624};
    Wh[10]='{32'd-725,32'd6064,32'd1993,32'd2310,32'd1364,32'd3750,32'd-2352,32'd3896,32'd-299,32'd-1916,32'd-2211,32'd2294,32'd7377,32'd-128,32'd-1846,32'd4465,32'd3981,32'd-236,32'd2770,32'd-3522,32'd739,32'd-4216,32'd-5429,32'd-1472,32'd-181,32'd-1613,32'd-1315,32'd-392,32'd1546,32'd3012,32'd1533,32'd-707,32'd3205,32'd1074,32'd5693,32'd463,32'd-3845,32'd829,32'd-1055,32'd7250,32'd1285,32'd-3427,32'd-2490,32'd4729,32'd-2775,32'd1599,32'd3835,32'd-493,32'd-3166,32'd30,32'd-462,32'd1308,32'd-1807,32'd-734,32'd-5898,32'd6904,32'd3376,32'd2985,32'd-914,32'd-2958,32'd-1915,32'd311,32'd4594,32'd-143,32'd-2218,32'd-3374,32'd558,32'd7236,32'd5175,32'd-3911,32'd3803,32'd6210,32'd-831,32'd105,32'd-214,32'd558,32'd4704,32'd8232,32'd58,32'd-3395,32'd-972,32'd10166,32'd-906,32'd-3208,32'd-2539,32'd4494,32'd-1040,32'd87,32'd-3901,32'd1123,32'd5742,32'd-2242,32'd10937,32'd-2666,32'd7944,32'd888,32'd-3193,32'd1903,32'd3459,32'd-2108,32'd-855,32'd4438,32'd1207,32'd8505,32'd-382,32'd1335,32'd-1678,32'd-6230,32'd5366,32'd-1188,32'd5869,32'd5029,32'd4548,32'd1568,32'd4707,32'd1011,32'd-1480,32'd6801,32'd-2493,32'd-12724,32'd172,32'd384,32'd-4777,32'd7500,32'd3071,32'd-8740,32'd11591,32'd-4082,32'd-8793,32'd-1104,32'd-3854,32'd-2246,32'd-6064,32'd5141,32'd-2734,32'd-2072,32'd-3212,32'd679,32'd-5942,32'd-2132,32'd3945,32'd2226,32'd-4455,32'd4733,32'd-1513,32'd706,32'd4143,32'd-2902,32'd-1416,32'd-2849,32'd-448,32'd3559,32'd-4829,32'd-2873,32'd-686,32'd620,32'd-9726,32'd2692,32'd2502,32'd-162,32'd-13935,32'd4353,32'd1569,32'd-7685,32'd8120,32'd6723,32'd3273,32'd3188,32'd468,32'd-1958,32'd-2435,32'd203,32'd-1762,32'd4401,32'd1439,32'd-6972,32'd5854,32'd-2072,32'd3603,32'd-3811,32'd-1585,32'd-10117,32'd6933,32'd491,32'd-634,32'd2131,32'd1317,32'd3681,32'd-1539,32'd5805,32'd-10214,32'd-4868,32'd-864,32'd4453,32'd2204,32'd1790,32'd2220,32'd-3579,32'd7460,32'd1613,32'd-1021,32'd1993,32'd-2078,32'd-7070,32'd-1307,32'd432,32'd-1124,32'd1035,32'd7739,32'd-2719,32'd-3076,32'd-456,32'd-8784,32'd2536,32'd3720,32'd-2095,32'd2690,32'd8388,32'd-2834,32'd-1832,32'd-1223,32'd354,32'd-1522,32'd-91,32'd-2817,32'd-11220,32'd2915,32'd-187,32'd-4057,32'd-4819,32'd-4914,32'd7856,32'd-3486,32'd-1235,32'd554,32'd-1265,32'd-2751,32'd2301,32'd3737,32'd447,32'd-1064,32'd2658,32'd-1413,32'd8867,32'd2988,32'd-919,32'd-1263,32'd-1026,32'd-3967,32'd-4599,32'd-4370,32'd539,32'd-1801,32'd-94,32'd-5048,32'd-5732,32'd-4323,32'd-1795,32'd-282,32'd-1767,32'd2946,32'd477,32'd3840,32'd-903,32'd2644,32'd-7397,32'd44,32'd-130,32'd1823,32'd-2470,32'd1610,32'd2016,32'd346,32'd-2294,32'd-844,32'd2340,32'd5263,32'd-6582,32'd-785,32'd2468,32'd10849,32'd-1717,32'd-1986,32'd-2629,32'd37,32'd6997,32'd-1542,32'd5224,32'd3886,32'd-116,32'd10615,32'd3535,32'd-4584,32'd2919,32'd2080,32'd-2279,32'd570,32'd-1715,32'd2127,32'd-1877,32'd1132,32'd2807,32'd6879,32'd1243,32'd1928,32'd12080,32'd1833,32'd4257,32'd-1481,32'd-2770,32'd-811,32'd5405,32'd-1041,32'd-3889,32'd-2944,32'd516,32'd4816,32'd1494,32'd7368,32'd-625,32'd-304,32'd-2236,32'd3911,32'd-1896,32'd-1746,32'd1630,32'd2790,32'd3493,32'd5844,32'd3005,32'd-171,32'd-147,32'd3103,32'd-1533,32'd-980,32'd-1867,32'd-621,32'd-94,32'd5971,32'd-3066,32'd363,32'd-279,32'd2412,32'd2915,32'd3908,32'd-2015,32'd2438,32'd-891,32'd-3378,32'd1121,32'd6015,32'd78,32'd3310,32'd-6005,32'd-3369,32'd3374,32'd853,32'd812,32'd1185,32'd-58,32'd-3085,32'd-3879,32'd4670,32'd-2148,32'd6347,32'd-7006,32'd3439,32'd6367,32'd862,32'd-3784,32'd4184,32'd7846,32'd4047,32'd-3312,32'd5351,32'd-159,32'd1395,32'd331,32'd5908,32'd236,32'd4230,32'd-1583,32'd507,32'd291,32'd-2702,32'd3530,32'd-1915,32'd7563,32'd924,32'd-3005,32'd6748,32'd-3876,32'd4931,32'd2883,32'd2800,32'd5180,32'd1701,32'd827,32'd-5043,32'd-5112};
    Wh[11]='{32'd1755,32'd3503,32'd730,32'd511,32'd-2644,32'd-1209,32'd880,32'd617,32'd3742,32'd1267,32'd-1257,32'd-1746,32'd-1163,32'd3225,32'd-856,32'd2250,32'd3120,32'd1384,32'd-3686,32'd-1940,32'd-705,32'd-502,32'd429,32'd-437,32'd-1583,32'd-35,32'd614,32'd-27,32'd-297,32'd-544,32'd-2493,32'd-122,32'd3125,32'd-569,32'd-11,32'd-2509,32'd-2470,32'd-2827,32'd-1436,32'd-597,32'd6035,32'd1373,32'd-942,32'd2009,32'd-3688,32'd-1165,32'd-1093,32'd266,32'd-5288,32'd-591,32'd-177,32'd3068,32'd-3298,32'd-3044,32'd3754,32'd-225,32'd2788,32'd-4020,32'd-302,32'd-247,32'd-734,32'd-75,32'd-128,32'd-167,32'd6015,32'd-2362,32'd2976,32'd-560,32'd-2893,32'd3149,32'd-1944,32'd-117,32'd2687,32'd1679,32'd-1424,32'd-2231,32'd-152,32'd-1820,32'd1545,32'd-3933,32'd455,32'd2563,32'd820,32'd2685,32'd-797,32'd2026,32'd-1345,32'd-1160,32'd4509,32'd-319,32'd-4436,32'd-1220,32'd-196,32'd-1268,32'd769,32'd-1069,32'd182,32'd-2741,32'd-2257,32'd1428,32'd-2004,32'd2171,32'd1933,32'd1510,32'd3564,32'd2482,32'd2563,32'd3747,32'd6181,32'd-3437,32'd2247,32'd-7978,32'd4697,32'd1604,32'd-339,32'd1572,32'd-5390,32'd-1044,32'd-5185,32'd-5146,32'd-501,32'd1796,32'd-1368,32'd-1683,32'd742,32'd-3239,32'd-2374,32'd2358,32'd-410,32'd-1953,32'd-7988,32'd-517,32'd3215,32'd-1468,32'd-3071,32'd-2274,32'd-933,32'd518,32'd-1553,32'd-1774,32'd-1210,32'd321,32'd1956,32'd2484,32'd-3598,32'd-4758,32'd-4843,32'd-252,32'd-1956,32'd748,32'd-608,32'd-1867,32'd299,32'd-6298,32'd1970,32'd5361,32'd-2194,32'd-2298,32'd-464,32'd4426,32'd2062,32'd2548,32'd4118,32'd883,32'd-480,32'd4846,32'd4475,32'd4514,32'd2807,32'd-1580,32'd823,32'd-331,32'd558,32'd-540,32'd-1254,32'd361,32'd-3627,32'd1276,32'd1850,32'd-434,32'd-1740,32'd4941,32'd3159,32'd-2966,32'd6669,32'd-2132,32'd-3610,32'd-6108,32'd1790,32'd2770,32'd-5053,32'd1370,32'd-6660,32'd-1224,32'd-1600,32'd-961,32'd-913,32'd2863,32'd1474,32'd-1478,32'd-862,32'd-616,32'd1558,32'd344,32'd1092,32'd-656,32'd1904,32'd-429,32'd-640,32'd3793,32'd-4331,32'd1546,32'd-2164,32'd-3930,32'd995,32'd-9501,32'd-2348,32'd-2438,32'd-4201,32'd-4758,32'd-419,32'd-3142,32'd1312,32'd-4274,32'd-36,32'd1126,32'd132,32'd-624,32'd-3232,32'd-44,32'd3579,32'd-1343,32'd1331,32'd-5717,32'd-5449,32'd-317,32'd2729,32'd545,32'd-4543,32'd48,32'd1422,32'd-2022,32'd963,32'd-1495,32'd-2707,32'd1549,32'd-1220,32'd594,32'd-2871,32'd-3486,32'd1082,32'd-1811,32'd814,32'd4248,32'd4597,32'd-710,32'd-974,32'd569,32'd2420,32'd-4125,32'd3120,32'd1948,32'd-2468,32'd-3034,32'd-308,32'd-2473,32'd-222,32'd2070,32'd-1486,32'd2080,32'd-53,32'd513,32'd993,32'd844,32'd912,32'd2150,32'd-6333,32'd-2727,32'd1174,32'd3168,32'd8198,32'd5585,32'd2683,32'd1995,32'd-485,32'd-793,32'd-3742,32'd2683,32'd13,32'd-1778,32'd-1049,32'd2556,32'd1186,32'd-736,32'd-638,32'd-238,32'd-147,32'd-5498,32'd169,32'd-1582,32'd1560,32'd1812,32'd979,32'd2690,32'd-98,32'd1632,32'd76,32'd820,32'd-4921,32'd2731,32'd-94,32'd971,32'd-1978,32'd1385,32'd-1184,32'd2380,32'd-949,32'd-1159,32'd2491,32'd4768,32'd2331,32'd4335,32'd3117,32'd938,32'd-4367,32'd-799,32'd3786,32'd823,32'd-3491,32'd2985,32'd71,32'd-76,32'd1481,32'd-2036,32'd-4577,32'd-1418,32'd-4121,32'd656,32'd825,32'd-7,32'd3095,32'd-4936,32'd-455,32'd-3298,32'd-2137,32'd-2739,32'd-3671,32'd-2980,32'd7382,32'd-1192,32'd-2154,32'd173,32'd-957,32'd-2436,32'd1545,32'd-3728,32'd-2873,32'd2231,32'd-809,32'd-48,32'd3823,32'd1728,32'd-78,32'd-837,32'd1569,32'd-2387,32'd3457,32'd4345,32'd-217,32'd484,32'd-5581,32'd-3120,32'd-606,32'd-4064,32'd-852,32'd-1448,32'd2595,32'd-3669,32'd-4938,32'd4311,32'd5468,32'd3698,32'd1756,32'd257,32'd-3918,32'd-4306,32'd-4809,32'd843,32'd775,32'd5356,32'd-4882,32'd-124,32'd292,32'd-1060,32'd1258,32'd-1601,32'd3256,32'd-313,32'd-3723,32'd-4531};
    Wh[12]='{32'd4030,32'd-146,32'd189,32'd2648,32'd929,32'd-1872,32'd-4299,32'd3754,32'd4252,32'd2736,32'd-444,32'd-1186,32'd-3483,32'd-88,32'd-3034,32'd853,32'd-1051,32'd8750,32'd-4589,32'd-3713,32'd870,32'd1102,32'd-3000,32'd2148,32'd4985,32'd-3779,32'd-331,32'd-1032,32'd-14716,32'd791,32'd2797,32'd-7294,32'd3488,32'd980,32'd-3759,32'd-2203,32'd-597,32'd-2336,32'd-1284,32'd3791,32'd3188,32'd3439,32'd3764,32'd2012,32'd-9365,32'd629,32'd-928,32'd203,32'd-1458,32'd3151,32'd-6904,32'd-745,32'd-1650,32'd2807,32'd652,32'd4729,32'd2912,32'd546,32'd1452,32'd5610,32'd3603,32'd1257,32'd3405,32'd-17,32'd1688,32'd-3347,32'd3378,32'd-605,32'd-2435,32'd-814,32'd-8759,32'd-9975,32'd-3579,32'd6293,32'd2105,32'd5205,32'd-690,32'd-384,32'd-3366,32'd1258,32'd-871,32'd-1500,32'd6225,32'd371,32'd3837,32'd1065,32'd2220,32'd-2697,32'd-2023,32'd-4221,32'd822,32'd-1352,32'd7788,32'd921,32'd-2437,32'd-1177,32'd5781,32'd2954,32'd-6093,32'd452,32'd-2880,32'd-814,32'd1816,32'd-8056,32'd-1442,32'd2824,32'd-3220,32'd4750,32'd4829,32'd-5771,32'd3879,32'd11943,32'd-1008,32'd-674,32'd1264,32'd3085,32'd-840,32'd2370,32'd-741,32'd-2646,32'd-2116,32'd2932,32'd-8369,32'd-2949,32'd2629,32'd4511,32'd-3439,32'd-1721,32'd-311,32'd1824,32'd-12343,32'd4208,32'd1878,32'd-373,32'd-112,32'd1707,32'd5039,32'd582,32'd5380,32'd-6362,32'd-396,32'd-3312,32'd-92,32'd488,32'd-2990,32'd372,32'd-4238,32'd-7055,32'd-468,32'd332,32'd-3518,32'd-729,32'd-2678,32'd4372,32'd-4125,32'd2861,32'd-5864,32'd-819,32'd1982,32'd-2521,32'd10537,32'd-2075,32'd-3449,32'd5927,32'd-2500,32'd2127,32'd-1752,32'd2917,32'd643,32'd-1101,32'd4125,32'd3041,32'd10605,32'd-132,32'd-3410,32'd-4768,32'd-874,32'd1503,32'd4558,32'd1105,32'd-4035,32'd-622,32'd4113,32'd-2963,32'd6220,32'd-3022,32'd-3010,32'd-826,32'd-5327,32'd656,32'd-1640,32'd1373,32'd-3735,32'd-913,32'd2376,32'd-1594,32'd-880,32'd1146,32'd220,32'd1014,32'd7,32'd-6489,32'd-2,32'd-38,32'd1168,32'd-1489,32'd-5683,32'd27,32'd-1655,32'd-1871,32'd3046,32'd-1546,32'd887,32'd2314,32'd-2800,32'd-2344,32'd-3984,32'd1235,32'd-4179,32'd-1446,32'd1027,32'd-3088,32'd-8354,32'd3039,32'd3613,32'd3459,32'd-2868,32'd-4479,32'd4572,32'd3847,32'd-3642,32'd-2631,32'd-13857,32'd-494,32'd998,32'd4575,32'd-4787,32'd-5664,32'd524,32'd1002,32'd-245,32'd1787,32'd-459,32'd-419,32'd-509,32'd427,32'd3308,32'd-1623,32'd-7324,32'd-2105,32'd70,32'd2580,32'd11,32'd341,32'd-1165,32'd-1101,32'd-2333,32'd6113,32'd1539,32'd-6347,32'd-2133,32'd6118,32'd4763,32'd-2235,32'd-921,32'd-771,32'd1799,32'd-3288,32'd-142,32'd297,32'd3269,32'd-3967,32'd4509,32'd-2368,32'd3918,32'd-180,32'd5117,32'd-3134,32'd-2536,32'd-2056,32'd6767,32'd-6542,32'd-5483,32'd3327,32'd161,32'd844,32'd547,32'd-12763,32'd2481,32'd499,32'd223,32'd1021,32'd-3457,32'd5043,32'd-1962,32'd-8559,32'd-767,32'd-105,32'd1467,32'd1029,32'd-850,32'd26,32'd6005,32'd3950,32'd56,32'd-1436,32'd-6806,32'd-507,32'd1883,32'd-1832,32'd4433,32'd-5126,32'd-247,32'd624,32'd-3549,32'd7548,32'd-3283,32'd5966,32'd-2127,32'd-2473,32'd7299,32'd-2529,32'd-510,32'd321,32'd3808,32'd1667,32'd-2421,32'd-1209,32'd-4235,32'd-115,32'd628,32'd-4252,32'd3996,32'd5361,32'd-3854,32'd1997,32'd-4663,32'd-3630,32'd4804,32'd709,32'd-2319,32'd-4672,32'd6318,32'd1182,32'd925,32'd1278,32'd-5810,32'd-535,32'd-2250,32'd3676,32'd-4323,32'd744,32'd5014,32'd5732,32'd-3483,32'd-413,32'd-298,32'd278,32'd4648,32'd156,32'd-2498,32'd2644,32'd4204,32'd-817,32'd-5029,32'd5468,32'd5659,32'd-2352,32'd1127,32'd2900,32'd-742,32'd-5117,32'd810,32'd3576,32'd-546,32'd-1407,32'd-2836,32'd5097,32'd-2834,32'd-3945,32'd4975,32'd-6093,32'd-3107,32'd-1766,32'd4514,32'd-2406,32'd2312,32'd-8496,32'd-7075,32'd5883,32'd4223,32'd451,32'd6049,32'd698,32'd-4382,32'd-7646,32'd4011,32'd-1723,32'd-6547,32'd-137};
    Wh[13]='{32'd1318,32'd-2736,32'd2849,32'd3657,32'd798,32'd1824,32'd1989,32'd-4602,32'd-1994,32'd978,32'd-247,32'd-5498,32'd1223,32'd1021,32'd-3222,32'd-7114,32'd4125,32'd1633,32'd-1746,32'd2127,32'd129,32'd5488,32'd-2197,32'd1645,32'd-884,32'd-2239,32'd-3540,32'd-502,32'd-2414,32'd1193,32'd-853,32'd4821,32'd5092,32'd583,32'd1475,32'd1105,32'd-1662,32'd-6459,32'd-2354,32'd6025,32'd6430,32'd6562,32'd-3720,32'd1341,32'd2088,32'd5966,32'd-7036,32'd4489,32'd-288,32'd-1296,32'd3356,32'd1312,32'd3083,32'd-3356,32'd-4018,32'd2266,32'd2822,32'd2519,32'd3388,32'd1905,32'd-372,32'd-6064,32'd1436,32'd-2749,32'd-2995,32'd3859,32'd619,32'd1166,32'd5415,32'd-4335,32'd219,32'd3046,32'd-7036,32'd-989,32'd-28,32'd-949,32'd8540,32'd-811,32'd-3098,32'd4228,32'd67,32'd-65,32'd-3984,32'd8496,32'd231,32'd-1345,32'd-1629,32'd1166,32'd-2907,32'd1046,32'd1807,32'd4196,32'd-1756,32'd-3264,32'd2666,32'd2014,32'd-2183,32'd-499,32'd4116,32'd2224,32'd-7163,32'd2213,32'd422,32'd-7285,32'd1231,32'd1849,32'd-1857,32'd600,32'd5444,32'd-4624,32'd-4709,32'd-2827,32'd2561,32'd1593,32'd2193,32'd-239,32'd3708,32'd5800,32'd2384,32'd145,32'd2507,32'd3398,32'd-2668,32'd8330,32'd5371,32'd-12255,32'd10439,32'd86,32'd-6557,32'd-2351,32'd2502,32'd-569,32'd-71,32'd13,32'd611,32'd-1937,32'd1253,32'd-7373,32'd-2014,32'd1147,32'd-390,32'd779,32'd-3793,32'd-7495,32'd3105,32'd-3864,32'd120,32'd-5195,32'd1944,32'd-199,32'd412,32'd-1334,32'd8032,32'd-59,32'd4147,32'd-1,32'd5898,32'd2460,32'd2111,32'd-6020,32'd525,32'd3183,32'd-3024,32'd-7202,32'd5092,32'd-2770,32'd-3601,32'd-765,32'd-614,32'd1469,32'd-3894,32'd6176,32'd-8515,32'd4692,32'd1324,32'd-867,32'd-3493,32'd-4641,32'd-2622,32'd2309,32'd5961,32'd-3933,32'd-5908,32'd-5249,32'd-1008,32'd563,32'd-217,32'd2980,32'd-5771,32'd-256,32'd-3574,32'd-3723,32'd-7031,32'd-2641,32'd-1616,32'd2099,32'd8012,32'd-4423,32'd6513,32'd-1706,32'd1101,32'd1416,32'd-1083,32'd-10097,32'd-3220,32'd-1420,32'd-4155,32'd1971,32'd5156,32'd2983,32'd-2724,32'd1291,32'd1236,32'd1785,32'd-660,32'd-294,32'd3642,32'd242,32'd-1186,32'd-906,32'd-288,32'd8432,32'd3405,32'd1448,32'd1199,32'd-4255,32'd-4069,32'd-411,32'd1202,32'd-2340,32'd-577,32'd1956,32'd-2161,32'd1954,32'd1446,32'd-2897,32'd5693,32'd855,32'd2976,32'd4536,32'd-5151,32'd800,32'd1583,32'd-994,32'd2386,32'd-445,32'd4973,32'd-3898,32'd-1550,32'd-3000,32'd-3093,32'd560,32'd-2810,32'd1024,32'd444,32'd-160,32'd-3344,32'd-661,32'd2019,32'd1237,32'd4187,32'd-2565,32'd1165,32'd-1955,32'd-726,32'd2419,32'd-1425,32'd1144,32'd870,32'd-30,32'd-3225,32'd1739,32'd1898,32'd-1027,32'd1545,32'd-956,32'd-2458,32'd-2347,32'd-4592,32'd-3298,32'd-7226,32'd1947,32'd-410,32'd-2829,32'd-863,32'd-1617,32'd32,32'd-7,32'd-643,32'd2019,32'd-726,32'd-5043,32'd-964,32'd1362,32'd-809,32'd-4772,32'd1330,32'd-5541,32'd-2381,32'd-3029,32'd185,32'd-2426,32'd-4313,32'd-647,32'd-1618,32'd690,32'd2832,32'd-7470,32'd-4020,32'd1883,32'd203,32'd-8193,32'd-983,32'd-7109,32'd-2536,32'd7651,32'd6596,32'd-3264,32'd-4545,32'd1257,32'd-881,32'd10380,32'd3315,32'd998,32'd507,32'd-1812,32'd-1036,32'd844,32'd5312,32'd232,32'd-2078,32'd-806,32'd-1026,32'd701,32'd-5747,32'd5922,32'd2695,32'd-3557,32'd1928,32'd-2968,32'd3430,32'd583,32'd613,32'd3425,32'd2746,32'd2045,32'd262,32'd1643,32'd480,32'd-2548,32'd4821,32'd207,32'd701,32'd1423,32'd3217,32'd-443,32'd1473,32'd2188,32'd-194,32'd-1021,32'd1734,32'd-6875,32'd-1651,32'd1704,32'd6787,32'd5317,32'd8857,32'd-2534,32'd1958,32'd1859,32'd1178,32'd2519,32'd-3896,32'd-7553,32'd-2517,32'd-6665,32'd5957,32'd-4887,32'd988,32'd-1685,32'd-2474,32'd1667,32'd-4841,32'd1883,32'd69,32'd1318,32'd-8032,32'd2110,32'd-5410,32'd4570,32'd2958,32'd581,32'd592,32'd-1066,32'd-572,32'd-160,32'd-3857,32'd31,32'd3659,32'd789};
    Wh[14]='{32'd2225,32'd-6958,32'd-1249,32'd2617,32'd1492,32'd2277,32'd-519,32'd2041,32'd-2614,32'd2968,32'd-5209,32'd89,32'd5507,32'd2071,32'd5053,32'd-8706,32'd4592,32'd2008,32'd4799,32'd5366,32'd1312,32'd2717,32'd3493,32'd48,32'd2844,32'd4707,32'd3918,32'd-520,32'd3041,32'd3188,32'd-1232,32'd3076,32'd-476,32'd-80,32'd-4572,32'd-750,32'd-3911,32'd1906,32'd890,32'd-4062,32'd7861,32'd-19,32'd596,32'd4714,32'd2546,32'd6064,32'd8183,32'd-2473,32'd-4208,32'd-1194,32'd-1162,32'd626,32'd-2056,32'd1340,32'd1066,32'd-4694,32'd1888,32'd2404,32'd-2396,32'd1017,32'd-1610,32'd3847,32'd3222,32'd2504,32'd2656,32'd891,32'd-2924,32'd1017,32'd3005,32'd4291,32'd-619,32'd-1855,32'd2851,32'd8291,32'd776,32'd5776,32'd-2368,32'd1274,32'd-3085,32'd617,32'd-950,32'd4853,32'd-1936,32'd6103,32'd2675,32'd166,32'd-4311,32'd638,32'd3129,32'd-1093,32'd-1289,32'd3937,32'd700,32'd-1572,32'd1054,32'd70,32'd3720,32'd-743,32'd2261,32'd4536,32'd-1600,32'd334,32'd2399,32'd-25,32'd5483,32'd-76,32'd3173,32'd8774,32'd1676,32'd2529,32'd3125,32'd910,32'd-14199,32'd-4072,32'd-1970,32'd-717,32'd1628,32'd-1392,32'd3686,32'd7998,32'd-294,32'd-835,32'd-6508,32'd-2261,32'd-2905,32'd4042,32'd-3225,32'd1628,32'd786,32'd6123,32'd2565,32'd-3850,32'd384,32'd914,32'd502,32'd4101,32'd1414,32'd-4284,32'd679,32'd-2541,32'd1569,32'd686,32'd-292,32'd3742,32'd-3933,32'd-3107,32'd2017,32'd-2846,32'd737,32'd-3962,32'd-285,32'd592,32'd130,32'd-982,32'd812,32'd-6811,32'd5751,32'd-1445,32'd-3676,32'd-11269,32'd684,32'd-4995,32'd-4216,32'd-6005,32'd272,32'd2597,32'd2141,32'd-3835,32'd2895,32'd-2546,32'd-1110,32'd527,32'd7978,32'd-3676,32'd-1427,32'd-98,32'd-3747,32'd-1549,32'd3425,32'd-1213,32'd-699,32'd2548,32'd3581,32'd-5253,32'd-1949,32'd-2176,32'd-192,32'd1453,32'd3417,32'd-1530,32'd-1137,32'd-791,32'd-3088,32'd-1928,32'd-3491,32'd1445,32'd-2277,32'd877,32'd7729,32'd4030,32'd-584,32'd676,32'd-1446,32'd-1022,32'd-2517,32'd52,32'd-1313,32'd4565,32'd1097,32'd-2749,32'd-215,32'd1054,32'd851,32'd-918,32'd1467,32'd-3493,32'd-408,32'd-6982,32'd1365,32'd-856,32'd-2534,32'd1713,32'd3344,32'd-4616,32'd-3395,32'd9082,32'd-3132,32'd-1855,32'd-4016,32'd2509,32'd-653,32'd-83,32'd5996,32'd3215,32'd-642,32'd8959,32'd1491,32'd-1474,32'd-2448,32'd5590,32'd-5434,32'd-3332,32'd-1604,32'd-1676,32'd1324,32'd3447,32'd-2993,32'd-1150,32'd1311,32'd-839,32'd-1452,32'd-851,32'd-6118,32'd-3054,32'd-4897,32'd445,32'd-4423,32'd-8715,32'd1448,32'd-61,32'd3352,32'd-2073,32'd-1348,32'd-876,32'd2873,32'd-911,32'd-7431,32'd-1008,32'd269,32'd-1107,32'd1137,32'd3991,32'd-1097,32'd-125,32'd-6538,32'd7573,32'd-6499,32'd-1733,32'd-4338,32'd-1218,32'd-3088,32'd-1770,32'd-980,32'd1971,32'd-926,32'd262,32'd-700,32'd3825,32'd-220,32'd-1029,32'd4604,32'd-5869,32'd4377,32'd5688,32'd4067,32'd5092,32'd-987,32'd-1805,32'd3215,32'd2790,32'd-414,32'd-2031,32'd-5708,32'd4831,32'd-4313,32'd4196,32'd2834,32'd2500,32'd-1192,32'd-5581,32'd-95,32'd1280,32'd-1322,32'd-4240,32'd3784,32'd-2624,32'd9204,32'd1401,32'd2351,32'd50,32'd-2229,32'd-1247,32'd-2069,32'd4421,32'd1585,32'd1536,32'd6621,32'd-97,32'd6591,32'd4091,32'd588,32'd2209,32'd2402,32'd-2347,32'd-1035,32'd-405,32'd2250,32'd4348,32'd-795,32'd2191,32'd-1348,32'd5166,32'd-2175,32'd-6547,32'd-2163,32'd-1152,32'd5742,32'd-7592,32'd9238,32'd-846,32'd1193,32'd998,32'd-2556,32'd-6064,32'd-996,32'd3146,32'd-1422,32'd-1171,32'd-6269,32'd849,32'd7109,32'd753,32'd-2512,32'd-1048,32'd-5429,32'd-90,32'd86,32'd3413,32'd-3649,32'd6782,32'd-2213,32'd-989,32'd7045,32'd-6186,32'd8154,32'd684,32'd1181,32'd-1573,32'd151,32'd-1816,32'd-5219,32'd5092,32'd9560,32'd-3161,32'd-5307,32'd1793,32'd2722,32'd1226,32'd688,32'd4892,32'd4733,32'd-2519,32'd-3417,32'd4467,32'd-451,32'd5380,32'd3752,32'd1165,32'd6635,32'd1414};
    Wh[15]='{32'd4309,32'd3547,32'd-3256,32'd-3666,32'd832,32'd548,32'd-4868,32'd-1104,32'd2303,32'd4172,32'd547,32'd-2004,32'd700,32'd-4577,32'd672,32'd-9145,32'd-657,32'd4169,32'd761,32'd1593,32'd781,32'd599,32'd-2052,32'd1594,32'd5830,32'd809,32'd1374,32'd2797,32'd4655,32'd139,32'd-3325,32'd6259,32'd3708,32'd-1407,32'd-5126,32'd3840,32'd-3618,32'd-1646,32'd1213,32'd6933,32'd3872,32'd3569,32'd7973,32'd-3056,32'd5556,32'd262,32'd-11201,32'd-2125,32'd-6293,32'd383,32'd2426,32'd-503,32'd-6645,32'd5927,32'd5742,32'd-599,32'd-3332,32'd6362,32'd-6572,32'd9335,32'd-5502,32'd3679,32'd-3381,32'd12070,32'd4958,32'd1593,32'd-1817,32'd-3615,32'd-4477,32'd-630,32'd-3298,32'd-484,32'd-2275,32'd252,32'd2218,32'd-1029,32'd477,32'd75,32'd-1712,32'd469,32'd-330,32'd-659,32'd-2502,32'd5136,32'd-6186,32'd475,32'd-458,32'd1898,32'd-2695,32'd2600,32'd1572,32'd5981,32'd-3496,32'd-3171,32'd-6000,32'd136,32'd-5366,32'd9594,32'd-4504,32'd9121,32'd-8408,32'd2156,32'd1729,32'd-10380,32'd-8291,32'd-2110,32'd-3747,32'd-1064,32'd5732,32'd-5336,32'd599,32'd1300,32'd5815,32'd-2105,32'd2546,32'd-6772,32'd2336,32'd1704,32'd2661,32'd84,32'd-1591,32'd-2717,32'd5791,32'd-2905,32'd5463,32'd3127,32'd-5395,32'd-7006,32'd3103,32'd-2885,32'd7631,32'd-2631,32'd3991,32'd3776,32'd13818,32'd3010,32'd11220,32'd1735,32'd1099,32'd769,32'd4323,32'd-4086,32'd8012,32'd-1100,32'd-673,32'd-378,32'd6367,32'd-8754,32'd997,32'd4562,32'd168,32'd-2890,32'd-2641,32'd-2416,32'd-5468,32'd12187,32'd503,32'd-5488,32'd1654,32'd21816,32'd2368,32'd2490,32'd7802,32'd3061,32'd-2644,32'd-1248,32'd-564,32'd1075,32'd1794,32'd-2272,32'd-1452,32'd-519,32'd-2854,32'd-4245,32'd1927,32'd4628,32'd-1544,32'd559,32'd-3654,32'd1340,32'd1966,32'd-1179,32'd-4187,32'd1209,32'd1964,32'd1690,32'd-2086,32'd-180,32'd7734,32'd3242,32'd1706,32'd2585,32'd257,32'd-3874,32'd-6372,32'd5361,32'd3820,32'd2135,32'd-3410,32'd-2426,32'd2924,32'd-4287,32'd-3972,32'd-2463,32'd-2907,32'd1472,32'd-3671,32'd-7231,32'd5136,32'd3332,32'd-9326,32'd-2379,32'd10507,32'd-878,32'd-3674,32'd-7045,32'd-121,32'd-3640,32'd7163,32'd2604,32'd1679,32'd1878,32'd4616,32'd3911,32'd2824,32'd-58,32'd3002,32'd1295,32'd2634,32'd-2346,32'd9951,32'd-2164,32'd-2398,32'd2203,32'd-2266,32'd-1608,32'd4555,32'd3337,32'd-2961,32'd-1591,32'd878,32'd674,32'd-44,32'd-3356,32'd836,32'd189,32'd3269,32'd-2495,32'd578,32'd-1954,32'd-1997,32'd2749,32'd993,32'd643,32'd734,32'd-6958,32'd2309,32'd5351,32'd576,32'd-7597,32'd-4223,32'd-2558,32'd11816,32'd-3676,32'd-6372,32'd-6479,32'd2697,32'd-611,32'd1503,32'd-328,32'd-5727,32'd-2602,32'd4084,32'd-2281,32'd2374,32'd6894,32'd-4052,32'd427,32'd-2,32'd-3017,32'd5454,32'd-4912,32'd-173,32'd9033,32'd-765,32'd-59,32'd-1962,32'd-10576,32'd249,32'd3063,32'd5800,32'd3725,32'd-61,32'd-2104,32'd-2619,32'd-5830,32'd-9,32'd543,32'd-4287,32'd4294,32'd-2531,32'd6835,32'd-4133,32'd3039,32'd-5991,32'd-5043,32'd111,32'd1704,32'd-517,32'd2027,32'd-597,32'd-3364,32'd-1800,32'd3798,32'd-1740,32'd-8330,32'd-2347,32'd284,32'd6977,32'd-3176,32'd1925,32'd1043,32'd2624,32'd-3100,32'd3964,32'd4592,32'd-1112,32'd-1813,32'd-4196,32'd366,32'd2006,32'd3591,32'd1735,32'd-1391,32'd414,32'd-402,32'd-6679,32'd-4106,32'd6372,32'd-1684,32'd-2578,32'd-1763,32'd-3527,32'd-2592,32'd-1850,32'd1022,32'd2312,32'd6674,32'd-3461,32'd-80,32'd-3095,32'd4641,32'd-1335,32'd2700,32'd7670,32'd11972,32'd5830,32'd-5585,32'd2313,32'd-5390,32'd-6665,32'd-5092,32'd8437,32'd3308,32'd4350,32'd4060,32'd-8212,32'd-464,32'd3308,32'd-7451,32'd-1143,32'd4567,32'd-2060,32'd-2814,32'd-26,32'd-1525,32'd7089,32'd-1284,32'd-4199,32'd-5380,32'd834,32'd14111,32'd-5122,32'd2714,32'd-93,32'd-707,32'd-7270,32'd-2946,32'd-2083,32'd-4846,32'd-509,32'd-3205,32'd-1385,32'd636,32'd1910,32'd-1177,32'd-3220,32'd-2446,32'd-1134,32'd1187};
    Wh[16]='{32'd2117,32'd1224,32'd-2548,32'd3327,32'd1593,32'd-1968,32'd694,32'd7031,32'd1459,32'd-1108,32'd-1901,32'd2066,32'd3347,32'd-3466,32'd-3774,32'd5478,32'd2239,32'd575,32'd4030,32'd1287,32'd-6411,32'd4602,32'd-4707,32'd1260,32'd848,32'd1904,32'd6787,32'd-3315,32'd6533,32'd-4519,32'd5307,32'd1702,32'd-418,32'd2077,32'd706,32'd1254,32'd1607,32'd34,32'd-3735,32'd4233,32'd3149,32'd4902,32'd1800,32'd2332,32'd2032,32'd-1690,32'd3325,32'd-3630,32'd-1851,32'd1920,32'd1138,32'd-5400,32'd5527,32'd1710,32'd5419,32'd-5649,32'd73,32'd-1270,32'd2047,32'd2739,32'd-5151,32'd3603,32'd5131,32'd-1822,32'd3679,32'd2770,32'd-1248,32'd-3598,32'd3745,32'd-4541,32'd2966,32'd219,32'd756,32'd184,32'd-1165,32'd6284,32'd3232,32'd1807,32'd2507,32'd-998,32'd1395,32'd6679,32'd9819,32'd-551,32'd3544,32'd-874,32'd1883,32'd5556,32'd-1823,32'd-641,32'd4040,32'd2541,32'd3449,32'd776,32'd-1403,32'd-1927,32'd-544,32'd2871,32'd5585,32'd1193,32'd-5527,32'd306,32'd589,32'd3330,32'd793,32'd4208,32'd6738,32'd1851,32'd18750,32'd-5283,32'd3828,32'd-9765,32'd3557,32'd1669,32'd2071,32'd791,32'd4846,32'd9770,32'd-748,32'd1614,32'd167,32'd16269,32'd7324,32'd7480,32'd-7021,32'd-546,32'd211,32'd1279,32'd-4519,32'd2829,32'd103,32'd726,32'd-2597,32'd4868,32'd6845,32'd8515,32'd16728,32'd-2215,32'd2028,32'd1094,32'd8203,32'd1560,32'd-5771,32'd240,32'd169,32'd2917,32'd9101,32'd-11718,32'd346,32'd-1854,32'd6748,32'd1458,32'd653,32'd3989,32'd-4594,32'd3918,32'd8813,32'd1048,32'd-5659,32'd2122,32'd932,32'd717,32'd-204,32'd735,32'd1711,32'd-5419,32'd-312,32'd4814,32'd-5961,32'd2178,32'd-1833,32'd-6337,32'd-297,32'd1724,32'd3088,32'd2978,32'd455,32'd-5283,32'd-875,32'd-3703,32'd5615,32'd3620,32'd-2188,32'd-4580,32'd-5747,32'd4970,32'd-2717,32'd4545,32'd-692,32'd-1396,32'd-4956,32'd-2144,32'd5961,32'd-6127,32'd-4858,32'd10224,32'd4089,32'd-5087,32'd11357,32'd1981,32'd-3505,32'd123,32'd73,32'd-8930,32'd4414,32'd-1185,32'd-4282,32'd-3212,32'd977,32'd2357,32'd-9350,32'd-240,32'd2124,32'd703,32'd-428,32'd-2307,32'd1456,32'd7963,32'd-1628,32'd-1130,32'd-3212,32'd-4702,32'd712,32'd-4150,32'd3183,32'd-4792,32'd-5385,32'd2404,32'd-7861,32'd661,32'd-141,32'd304,32'd-3508,32'd923,32'd1593,32'd-4548,32'd-817,32'd-927,32'd1,32'd58,32'd956,32'd1495,32'd-4042,32'd3640,32'd2612,32'd1152,32'd-3388,32'd392,32'd-6113,32'd-963,32'd-5449,32'd-4902,32'd2269,32'd2766,32'd186,32'd-341,32'd-379,32'd-3659,32'd4235,32'd-2338,32'd-2622,32'd-1065,32'd2839,32'd-5375,32'd-9326,32'd-5883,32'd795,32'd-1074,32'd-917,32'd-3544,32'd865,32'd428,32'd-4462,32'd-181,32'd-5712,32'd-3554,32'd-3405,32'd-11767,32'd-2210,32'd-4196,32'd-928,32'd2534,32'd-1641,32'd-321,32'd-2612,32'd-3623,32'd-2941,32'd-7177,32'd-761,32'd-2293,32'd15937,32'd-2744,32'd-2408,32'd-5717,32'd2416,32'd1351,32'd-3654,32'd-7758,32'd-2080,32'd-3471,32'd-2998,32'd-335,32'd3063,32'd-2924,32'd2119,32'd-1185,32'd300,32'd297,32'd-2697,32'd-3371,32'd5253,32'd-5029,32'd-3007,32'd-5571,32'd-2177,32'd1162,32'd-2563,32'd3947,32'd-576,32'd4528,32'd5737,32'd265,32'd-3183,32'd-8061,32'd-2114,32'd-1259,32'd2995,32'd5234,32'd-1795,32'd2795,32'd-745,32'd-769,32'd-1573,32'd-3679,32'd4875,32'd-2222,32'd-91,32'd2587,32'd2041,32'd-2966,32'd3269,32'd-981,32'd-206,32'd1508,32'd-1138,32'd-468,32'd1209,32'd1596,32'd-793,32'd3305,32'd-433,32'd3330,32'd2498,32'd-3852,32'd6127,32'd-248,32'd1601,32'd-5493,32'd2403,32'd4602,32'd-2141,32'd7,32'd-1280,32'd-3928,32'd1505,32'd4357,32'd-3850,32'd2324,32'd2875,32'd-8627,32'd-896,32'd-2932,32'd2180,32'd-6748,32'd809,32'd-212,32'd7651,32'd-231,32'd-806,32'd4287,32'd949,32'd6108,32'd-2053,32'd-3117,32'd8173,32'd-6713,32'd-6225,32'd2646,32'd1223,32'd4350,32'd2070,32'd195,32'd3984,32'd400,32'd-5463,32'd-4006,32'd-3093,32'd-154,32'd4042,32'd-5336};
    Wh[17]='{32'd2614,32'd1950,32'd188,32'd4067,32'd76,32'd2514,32'd-6132,32'd960,32'd5883,32'd2138,32'd4638,32'd5039,32'd-2008,32'd993,32'd4313,32'd-1335,32'd3933,32'd8251,32'd2434,32'd212,32'd1370,32'd2773,32'd1927,32'd856,32'd867,32'd1562,32'd2363,32'd-1771,32'd739,32'd-4343,32'd-1693,32'd-2983,32'd-1418,32'd-3269,32'd2619,32'd170,32'd-214,32'd1640,32'd523,32'd602,32'd-631,32'd-1494,32'd3457,32'd-3806,32'd-355,32'd-4052,32'd-2727,32'd4689,32'd6171,32'd2456,32'd1584,32'd2546,32'd-3032,32'd-6909,32'd-2856,32'd2673,32'd1658,32'd968,32'd2092,32'd-684,32'd4350,32'd-2670,32'd-4702,32'd-32,32'd1130,32'd3195,32'd-1209,32'd3635,32'd1870,32'd391,32'd378,32'd-856,32'd947,32'd1656,32'd-1088,32'd-218,32'd-4140,32'd-274,32'd-33,32'd-1311,32'd-475,32'd-870,32'd-4855,32'd-461,32'd3154,32'd2941,32'd2512,32'd68,32'd-61,32'd-3942,32'd1933,32'd-1732,32'd533,32'd-5283,32'd-2066,32'd429,32'd-2858,32'd673,32'd-3542,32'd2203,32'd-7905,32'd5097,32'd1157,32'd1593,32'd-2934,32'd-1464,32'd-3642,32'd2145,32'd-1433,32'd-9384,32'd8632,32'd2802,32'd3486,32'd-51,32'd3864,32'd-1993,32'd7250,32'd13554,32'd-8437,32'd-3281,32'd1424,32'd6533,32'd11660,32'd1938,32'd2044,32'd-13574,32'd-475,32'd-1124,32'd-1329,32'd4775,32'd3146,32'd3310,32'd244,32'd1828,32'd-1074,32'd5415,32'd-2810,32'd5859,32'd1575,32'd-422,32'd6484,32'd662,32'd659,32'd-3747,32'd-4694,32'd3232,32'd10029,32'd-3964,32'd-2556,32'd149,32'd6630,32'd2009,32'd-922,32'd149,32'd3310,32'd-1624,32'd741,32'd-2204,32'd5170,32'd7480,32'd2425,32'd-1290,32'd-3493,32'd5400,32'd-1955,32'd1213,32'd-1169,32'd3198,32'd-1510,32'd662,32'd2247,32'd5166,32'd2236,32'd98,32'd1148,32'd-1005,32'd1705,32'd-961,32'd-6625,32'd-3117,32'd2751,32'd-5883,32'd273,32'd1907,32'd-7358,32'd-336,32'd-71,32'd4870,32'd-2749,32'd-5600,32'd260,32'd-1650,32'd-344,32'd-646,32'd-587,32'd2910,32'd4697,32'd1630,32'd4814,32'd4099,32'd4738,32'd125,32'd-2497,32'd-1706,32'd4421,32'd376,32'd1429,32'd-295,32'd6884,32'd4143,32'd4328,32'd193,32'd10000,32'd5932,32'd-601,32'd-995,32'd1325,32'd740,32'd5952,32'd1145,32'd240,32'd-5117,32'd-4184,32'd235,32'd-1014,32'd-2380,32'd1701,32'd2302,32'd2320,32'd2368,32'd1630,32'd5717,32'd-1726,32'd4199,32'd-1197,32'd1806,32'd-3557,32'd-776,32'd620,32'd-125,32'd1746,32'd-3771,32'd-457,32'd1585,32'd1801,32'd4431,32'd-4833,32'd-1981,32'd-4138,32'd1954,32'd-4060,32'd-72,32'd2127,32'd4538,32'd363,32'd224,32'd2020,32'd1704,32'd540,32'd989,32'd4089,32'd1309,32'd3825,32'd-4738,32'd640,32'd1374,32'd-153,32'd2199,32'd-2452,32'd764,32'd3574,32'd-634,32'd-374,32'd-2951,32'd-1375,32'd-383,32'd7705,32'd-1124,32'd2205,32'd3708,32'd807,32'd1905,32'd2517,32'd-590,32'd1579,32'd-319,32'd-1361,32'd4428,32'd-3312,32'd-2347,32'd4743,32'd-5195,32'd-2683,32'd-5805,32'd-5532,32'd2467,32'd-2866,32'd-1525,32'd-4108,32'd-1130,32'd6762,32'd3605,32'd-2180,32'd6181,32'd-260,32'd527,32'd70,32'd2362,32'd983,32'd-5068,32'd1091,32'd2293,32'd-3068,32'd-3793,32'd1373,32'd6005,32'd-1220,32'd3881,32'd7094,32'd-3952,32'd-1936,32'd-41,32'd-932,32'd-2968,32'd-1040,32'd1398,32'd659,32'd6855,32'd-4201,32'd3496,32'd499,32'd-1927,32'd1551,32'd-1588,32'd-5009,32'd-4770,32'd1772,32'd4594,32'd1737,32'd3598,32'd-1229,32'd-2280,32'd2507,32'd1729,32'd1323,32'd-3063,32'd-867,32'd-425,32'd-3583,32'd-1127,32'd-1550,32'd3527,32'd1524,32'd858,32'd3903,32'd-4169,32'd3342,32'd-6923,32'd1765,32'd1148,32'd7568,32'd5126,32'd343,32'd-4418,32'd3378,32'd5800,32'd-2668,32'd2321,32'd4116,32'd708,32'd492,32'd-3869,32'd2619,32'd-1777,32'd4616,32'd344,32'd1856,32'd6967,32'd2268,32'd4748,32'd4492,32'd-8989,32'd-1392,32'd-4250,32'd4130,32'd-4919,32'd137,32'd1005,32'd-1978,32'd1639,32'd2265,32'd-2624,32'd7978,32'd-6591,32'd249,32'd-1867,32'd-3449,32'd4570,32'd-1190,32'd1394};
    Wh[18]='{32'd183,32'd-7089,32'd-76,32'd-3771,32'd-880,32'd-2636,32'd-9,32'd-1289,32'd-4899,32'd-223,32'd4978,32'd-1962,32'd-4587,32'd-617,32'd-2553,32'd-881,32'd5410,32'd-4694,32'd-48,32'd3103,32'd-302,32'd377,32'd1414,32'd-3710,32'd-931,32'd-2592,32'd378,32'd-723,32'd-1231,32'd-294,32'd-1267,32'd2480,32'd-5561,32'd2436,32'd2622,32'd1873,32'd-1733,32'd64,32'd-1427,32'd2724,32'd-1589,32'd1020,32'd-1645,32'd1409,32'd576,32'd-1281,32'd-1284,32'd599,32'd5566,32'd-4423,32'd-1116,32'd3066,32'd-236,32'd-538,32'd-628,32'd-1105,32'd1929,32'd-1834,32'd-283,32'd-3808,32'd1226,32'd-2072,32'd2387,32'd-1473,32'd-2142,32'd1435,32'd-299,32'd2851,32'd-2707,32'd-1617,32'd-4877,32'd4113,32'd-2491,32'd5747,32'd572,32'd-2263,32'd-895,32'd-3479,32'd562,32'd2298,32'd-1398,32'd1181,32'd-5947,32'd1317,32'd141,32'd-1047,32'd-534,32'd1851,32'd-3288,32'd-12,32'd-775,32'd-611,32'd-1513,32'd-1067,32'd-471,32'd1834,32'd484,32'd11054,32'd4709,32'd931,32'd-2541,32'd-2021,32'd1738,32'd1849,32'd-6083,32'd429,32'd-237,32'd2470,32'd-6113,32'd5434,32'd-8154,32'd5439,32'd-2836,32'd-2225,32'd3652,32'd-1527,32'd-186,32'd-4587,32'd-2773,32'd3081,32'd-2126,32'd2626,32'd1600,32'd3227,32'd-5390,32'd-822,32'd4428,32'd-2814,32'd-2285,32'd2597,32'd1489,32'd-2905,32'd-3269,32'd-1197,32'd-5410,32'd-2614,32'd-5957,32'd323,32'd4052,32'd3666,32'd1856,32'd-965,32'd1348,32'd-2666,32'd-3996,32'd3681,32'd-3732,32'd4245,32'd-1216,32'd-2717,32'd2410,32'd1923,32'd-3430,32'd2413,32'd3579,32'd-731,32'd-6806,32'd958,32'd-4614,32'd6728,32'd-1901,32'd528,32'd2076,32'd161,32'd-2220,32'd4572,32'd12,32'd1030,32'd2263,32'd-1059,32'd2053,32'd-4821,32'd-6625,32'd4809,32'd-1370,32'd-3913,32'd-2861,32'd-2556,32'd-4685,32'd-759,32'd710,32'd2824,32'd6337,32'd-1799,32'd7133,32'd1990,32'd-2056,32'd2849,32'd-3100,32'd3476,32'd3471,32'd2143,32'd-4040,32'd-4133,32'd-1488,32'd-8950,32'd-4443,32'd3125,32'd-1374,32'd264,32'd1589,32'd1514,32'd1779,32'd-293,32'd-2519,32'd-1251,32'd2130,32'd1021,32'd7905,32'd-284,32'd1787,32'd-4328,32'd308,32'd670,32'd1658,32'd5058,32'd107,32'd-2447,32'd3566,32'd2797,32'd118,32'd-469,32'd-3845,32'd367,32'd-3027,32'd681,32'd-1591,32'd-365,32'd3210,32'd7138,32'd4079,32'd3569,32'd1644,32'd-326,32'd-8,32'd-4326,32'd1270,32'd-1315,32'd2089,32'd-9760,32'd5439,32'd-3378,32'd10126,32'd-2202,32'd96,32'd550,32'd-2846,32'd316,32'd5166,32'd437,32'd-3354,32'd-174,32'd432,32'd-3996,32'd2897,32'd1784,32'd1497,32'd-1026,32'd-2541,32'd7050,32'd2270,32'd3193,32'd1121,32'd3356,32'd5268,32'd3603,32'd348,32'd-2668,32'd1525,32'd-517,32'd2464,32'd-3146,32'd3115,32'd-3894,32'd542,32'd-1155,32'd-2670,32'd-1124,32'd2282,32'd4990,32'd-3029,32'd-149,32'd4768,32'd62,32'd-1893,32'd3974,32'd1853,32'd2343,32'd-3247,32'd2152,32'd-491,32'd-550,32'd-849,32'd-2512,32'd-2376,32'd-1579,32'd3857,32'd-2058,32'd-57,32'd-1789,32'd1663,32'd-1610,32'd214,32'd-1490,32'd-1943,32'd7114,32'd4343,32'd2224,32'd878,32'd522,32'd1278,32'd-3933,32'd1820,32'd-3081,32'd1184,32'd1212,32'd-920,32'd121,32'd2458,32'd2260,32'd-1579,32'd5004,32'd1064,32'd1478,32'd-786,32'd1766,32'd4279,32'd744,32'd-289,32'd1903,32'd2132,32'd285,32'd-7114,32'd2653,32'd46,32'd2536,32'd-4665,32'd238,32'd-7519,32'd-2105,32'd1340,32'd-5224,32'd6157,32'd2524,32'd-6748,32'd-751,32'd-2822,32'd1683,32'd-1403,32'd-344,32'd2753,32'd1572,32'd-3813,32'd1986,32'd820,32'd-3464,32'd-604,32'd-1437,32'd-2496,32'd2858,32'd-2432,32'd-4216,32'd2224,32'd-3728,32'd-461,32'd784,32'd5000,32'd-3845,32'd-1072,32'd2700,32'd3723,32'd5053,32'd-1583,32'd-1064,32'd941,32'd-1712,32'd-3186,32'd-3466,32'd388,32'd599,32'd-2248,32'd156,32'd1687,32'd-2956,32'd-146,32'd-1021,32'd2037,32'd-1649,32'd-711,32'd3095,32'd-6030,32'd1953,32'd-7377,32'd4460,32'd2150,32'd2807,32'd2105,32'd1992,32'd3117,32'd761};
    Wh[19]='{32'd-1257,32'd-6694,32'd81,32'd5019,32'd-1503,32'd116,32'd2597,32'd-728,32'd-83,32'd-44,32'd3078,32'd3115,32'd539,32'd-4023,32'd7460,32'd-6928,32'd-1152,32'd4453,32'd276,32'd1459,32'd-842,32'd-2004,32'd1170,32'd-378,32'd-4475,32'd546,32'd3784,32'd2097,32'd2741,32'd3041,32'd-2308,32'd5102,32'd-5458,32'd-2524,32'd-4304,32'd-359,32'd-6181,32'd736,32'd-411,32'd735,32'd-1859,32'd-6235,32'd-1115,32'd1804,32'd10527,32'd-613,32'd-1767,32'd2391,32'd3574,32'd2268,32'd2470,32'd-3454,32'd7612,32'd1473,32'd1488,32'd-718,32'd-1568,32'd934,32'd48,32'd-1984,32'd1203,32'd4072,32'd260,32'd-697,32'd-2336,32'd7524,32'd-1439,32'd-1467,32'd774,32'd-575,32'd609,32'd3564,32'd-2810,32'd-2946,32'd-2841,32'd-783,32'd-1960,32'd-955,32'd2910,32'd1629,32'd-414,32'd-3718,32'd-3872,32'd1705,32'd701,32'd-3537,32'd-3308,32'd1214,32'd-34,32'd-2768,32'd-3969,32'd-4226,32'd-1030,32'd-2014,32'd-8779,32'd-41,32'd-1571,32'd-446,32'd3728,32'd-1818,32'd-2336,32'd1802,32'd-4157,32'd10195,32'd1800,32'd-1545,32'd7714,32'd10693,32'd-291,32'd-424,32'd1500,32'd-12275,32'd-1555,32'd3278,32'd5317,32'd3344,32'd4594,32'd7846,32'd190,32'd-47,32'd-33,32'd-3200,32'd3557,32'd1669,32'd-2773,32'd3415,32'd-3442,32'd-3498,32'd7963,32'd-17890,32'd6206,32'd-776,32'd-3640,32'd-606,32'd4501,32'd1413,32'd-1976,32'd-3515,32'd1502,32'd1165,32'd2482,32'd3493,32'd8134,32'd-2180,32'd1635,32'd-3483,32'd3190,32'd6030,32'd2539,32'd-3081,32'd1673,32'd4394,32'd3491,32'd1129,32'd-4108,32'd8183,32'd-5937,32'd-4340,32'd3208,32'd5371,32'd6528,32'd3784,32'd-113,32'd-699,32'd-167,32'd-6176,32'd2382,32'd-866,32'd-3486,32'd-895,32'd-3117,32'd-1295,32'd-2344,32'd2026,32'd-875,32'd2807,32'd3269,32'd-5034,32'd-1156,32'd1865,32'd3881,32'd-563,32'd6757,32'd9638,32'd5786,32'd5751,32'd2218,32'd10107,32'd36,32'd-5434,32'd1226,32'd-2100,32'd586,32'd-590,32'd-2388,32'd4973,32'd-476,32'd-4711,32'd-5942,32'd1226,32'd2663,32'd1490,32'd3188,32'd3305,32'd650,32'd327,32'd1834,32'd6245,32'd-3657,32'd-2927,32'd-2163,32'd2700,32'd4038,32'd-1257,32'd580,32'd5649,32'd6684,32'd-3942,32'd65,32'd-1534,32'd1646,32'd4184,32'd5639,32'd227,32'd-127,32'd1729,32'd6508,32'd-159,32'd-1022,32'd-2351,32'd894,32'd4807,32'd3715,32'd3234,32'd2500,32'd4045,32'd1287,32'd1937,32'd8857,32'd-6557,32'd-2836,32'd8090,32'd5244,32'd-3049,32'd-2802,32'd-1517,32'd1864,32'd789,32'd4658,32'd-2011,32'd-618,32'd182,32'd2102,32'd-1549,32'd-281,32'd-404,32'd2337,32'd-776,32'd-2490,32'd185,32'd-2421,32'd-4470,32'd1890,32'd4282,32'd491,32'd3020,32'd-1547,32'd-1319,32'd1287,32'd-1466,32'd-7724,32'd5263,32'd-1315,32'd-424,32'd-1009,32'd-2066,32'd-609,32'd1109,32'd-253,32'd1949,32'd-2279,32'd1679,32'd2421,32'd-210,32'd3425,32'd-2158,32'd1247,32'd1386,32'd-4626,32'd1234,32'd-8129,32'd-542,32'd2622,32'd-940,32'd3283,32'd1376,32'd-219,32'd1593,32'd6855,32'd-1519,32'd-3847,32'd-3867,32'd-5048,32'd-815,32'd-644,32'd-6323,32'd6215,32'd2083,32'd5742,32'd-1015,32'd7749,32'd-1364,32'd1972,32'd-1809,32'd-232,32'd-2098,32'd1718,32'd2227,32'd1032,32'd-159,32'd-3076,32'd5356,32'd3515,32'd-755,32'd769,32'd4328,32'd8383,32'd-2597,32'd2617,32'd591,32'd-3911,32'd6372,32'd-1336,32'd-1181,32'd-827,32'd7939,32'd-154,32'd-160,32'd-682,32'd2629,32'd-4709,32'd6899,32'd-242,32'd4863,32'd-331,32'd-5039,32'd3093,32'd3229,32'd-1385,32'd-839,32'd-620,32'd757,32'd-5683,32'd-2978,32'd-5156,32'd3425,32'd-1,32'd-13076,32'd-12929,32'd601,32'd-1192,32'd1128,32'd1469,32'd-3352,32'd-2225,32'd1158,32'd4206,32'd1044,32'd-973,32'd424,32'd7983,32'd2098,32'd-5351,32'd-6411,32'd-3239,32'd1860,32'd1899,32'd661,32'd4174,32'd4206,32'd-435,32'd5317,32'd5927,32'd110,32'd-95,32'd-7773,32'd-4245,32'd-5620,32'd-402,32'd-1579,32'd-9389,32'd6513,32'd-1066,32'd2275,32'd2841,32'd-4052,32'd-4082,32'd-898,32'd8388,32'd-1330};
    Wh[20]='{32'd-498,32'd-6962,32'd-2366,32'd-1527,32'd-14,32'd1022,32'd3635,32'd2658,32'd1043,32'd-2495,32'd-2297,32'd2177,32'd-621,32'd3083,32'd-210,32'd-1916,32'd-911,32'd1638,32'd-1871,32'd1039,32'd-2941,32'd-2004,32'd1859,32'd-1906,32'd-311,32'd-690,32'd620,32'd-2192,32'd1304,32'd-1672,32'd-544,32'd26,32'd-5737,32'd378,32'd-2971,32'd-2849,32'd-4797,32'd-1130,32'd617,32'd-539,32'd856,32'd-1726,32'd3156,32'd-2414,32'd4482,32'd2517,32'd4372,32'd1226,32'd-4248,32'd2092,32'd1975,32'd-1813,32'd1353,32'd34,32'd4826,32'd1254,32'd251,32'd-1361,32'd-3977,32'd4519,32'd3298,32'd-3112,32'd3288,32'd1004,32'd3530,32'd-326,32'd3964,32'd-2595,32'd-1224,32'd1879,32'd2907,32'd2895,32'd-1861,32'd2561,32'd-2639,32'd1635,32'd-1456,32'd-1459,32'd4057,32'd578,32'd-2963,32'd-5385,32'd1721,32'd-3908,32'd4035,32'd-1804,32'd-112,32'd1282,32'd1998,32'd1220,32'd-2285,32'd-5366,32'd1638,32'd-939,32'd-3913,32'd-414,32'd444,32'd-3537,32'd-1945,32'd-1520,32'd-2998,32'd-3911,32'd-3779,32'd-2761,32'd2285,32'd-1602,32'd40,32'd-2056,32'd-1049,32'd2182,32'd-1380,32'd5258,32'd-253,32'd-3681,32'd-1893,32'd-1665,32'd1270,32'd5517,32'd-756,32'd2832,32'd983,32'd-2104,32'd-1936,32'd-3105,32'd-1290,32'd246,32'd-1455,32'd-12,32'd2222,32'd13486,32'd-3842,32'd-1629,32'd-2431,32'd2822,32'd2091,32'd-2379,32'd1397,32'd364,32'd-1533,32'd1564,32'd352,32'd484,32'd-1160,32'd2312,32'd4038,32'd2003,32'd-3073,32'd5639,32'd1813,32'd-1439,32'd1027,32'd341,32'd5512,32'd-5229,32'd-3493,32'd-1423,32'd-35,32'd-2083,32'd2587,32'd-6152,32'd-3999,32'd-384,32'd1060,32'd-2963,32'd-2526,32'd-3554,32'd-6494,32'd1705,32'd-2685,32'd-6,32'd-3400,32'd-8193,32'd-3720,32'd7670,32'd1562,32'd-1877,32'd-3269,32'd1627,32'd1799,32'd2187,32'd1766,32'd-2824,32'd-3215,32'd2678,32'd2244,32'd2326,32'd872,32'd1560,32'd-3159,32'd3947,32'd-2963,32'd127,32'd-6708,32'd1835,32'd-656,32'd916,32'd176,32'd-1396,32'd-363,32'd-2454,32'd-930,32'd2751,32'd349,32'd1652,32'd-1374,32'd65,32'd1356,32'd2585,32'd-840,32'd242,32'd-9794,32'd-2583,32'd-2368,32'd-300,32'd687,32'd1993,32'd5864,32'd2053,32'd-6181,32'd-1199,32'd-317,32'd2054,32'd-4331,32'd2077,32'd-177,32'd-3100,32'd-5786,32'd742,32'd660,32'd-2034,32'd-1483,32'd6625,32'd2871,32'd-1070,32'd2277,32'd1614,32'd2993,32'd-505,32'd-1876,32'd-2271,32'd357,32'd6723,32'd-4309,32'd469,32'd4636,32'd1828,32'd-3293,32'd2293,32'd-1113,32'd-4487,32'd-1860,32'd-242,32'd-332,32'd-3859,32'd681,32'd4121,32'd-3847,32'd-743,32'd306,32'd-2778,32'd-1106,32'd-4470,32'd1783,32'd-370,32'd3535,32'd1818,32'd2464,32'd-983,32'd245,32'd900,32'd3029,32'd-2543,32'd-4130,32'd1492,32'd39,32'd3190,32'd1029,32'd-1342,32'd-7192,32'd-1240,32'd-3452,32'd-6289,32'd1163,32'd5537,32'd2307,32'd6059,32'd1191,32'd1323,32'd4125,32'd-2622,32'd-3459,32'd-2015,32'd-1888,32'd390,32'd5737,32'd99,32'd-4504,32'd2553,32'd-2690,32'd-3845,32'd-643,32'd-3383,32'd411,32'd-3166,32'd-2041,32'd-4174,32'd1129,32'd7421,32'd1611,32'd-2644,32'd-2739,32'd-131,32'd1335,32'd3134,32'd-299,32'd3071,32'd-4829,32'd1763,32'd-6391,32'd3203,32'd-6459,32'd268,32'd-1588,32'd-445,32'd-2641,32'd-604,32'd-562,32'd-3200,32'd3242,32'd640,32'd-4104,32'd-1391,32'd5976,32'd-1854,32'd-3715,32'd-2038,32'd3051,32'd62,32'd-1829,32'd1010,32'd-3347,32'd404,32'd-484,32'd2924,32'd1050,32'd1773,32'd-1329,32'd-1660,32'd-5786,32'd919,32'd2368,32'd3059,32'd-825,32'd289,32'd-765,32'd120,32'd-6733,32'd-10175,32'd-1818,32'd-4008,32'd-2573,32'd-5258,32'd3747,32'd-362,32'd855,32'd-3103,32'd744,32'd597,32'd-327,32'd-3725,32'd-560,32'd-1779,32'd-6484,32'd-2290,32'd-7651,32'd-823,32'd3032,32'd1571,32'd5483,32'd-2536,32'd15,32'd-2052,32'd-1683,32'd5541,32'd-1485,32'd1194,32'd174,32'd2590,32'd-924,32'd-1008,32'd1781,32'd2519,32'd1336,32'd2561,32'd6796,32'd-8198,32'd-1058,32'd3278,32'd-6162,32'd764};
    Wh[21]='{32'd-440,32'd-3913,32'd5195,32'd-854,32'd-2685,32'd-252,32'd-528,32'd-2573,32'd2376,32'd266,32'd2270,32'd-2502,32'd-295,32'd1602,32'd-6494,32'd2104,32'd1832,32'd-731,32'd-1517,32'd-603,32'd-2410,32'd-5268,32'd-278,32'd-3986,32'd-1395,32'd-36,32'd-3676,32'd-844,32'd809,32'd1220,32'd1915,32'd7431,32'd-2022,32'd-2191,32'd-3024,32'd-2043,32'd-1380,32'd1926,32'd1706,32'd1981,32'd-1165,32'd-1008,32'd-740,32'd-785,32'd2425,32'd-2553,32'd-4289,32'd1888,32'd-2143,32'd793,32'd7729,32'd1719,32'd12578,32'd896,32'd1059,32'd-1716,32'd1295,32'd2144,32'd-2985,32'd710,32'd-2607,32'd2893,32'd-1436,32'd-3383,32'd-583,32'd1243,32'd-2489,32'd751,32'd1436,32'd269,32'd-2578,32'd-644,32'd653,32'd-1083,32'd215,32'd1594,32'd-5444,32'd1336,32'd2160,32'd1069,32'd2103,32'd-1958,32'd-535,32'd634,32'd3176,32'd-5820,32'd-84,32'd-2519,32'd-1705,32'd-2646,32'd3198,32'd935,32'd-2093,32'd-675,32'd-3325,32'd1,32'd-922,32'd-5146,32'd-2202,32'd-2487,32'd855,32'd2468,32'd-2106,32'd5561,32'd1420,32'd1600,32'd-485,32'd1425,32'd-2761,32'd4467,32'd383,32'd-3640,32'd-5458,32'd1800,32'd1488,32'd174,32'd805,32'd2875,32'd2646,32'd-2749,32'd-1578,32'd-4399,32'd6469,32'd-2351,32'd3371,32'd-3354,32'd-2186,32'd488,32'd3349,32'd-2558,32'd1705,32'd-1262,32'd401,32'd-2326,32'd-3066,32'd-1495,32'd-2269,32'd-396,32'd680,32'd1166,32'd297,32'd1787,32'd-3540,32'd318,32'd-4096,32'd-556,32'd-1334,32'd1967,32'd3522,32'd406,32'd-49,32'd1796,32'd-2697,32'd-3310,32'd-2255,32'd4218,32'd1715,32'd-1712,32'd-2490,32'd8100,32'd5502,32'd3977,32'd-790,32'd5039,32'd659,32'd7016,32'd-1032,32'd-3381,32'd1202,32'd228,32'd-5410,32'd-3701,32'd7187,32'd3845,32'd4953,32'd587,32'd2103,32'd938,32'd2102,32'd764,32'd214,32'd-3002,32'd1774,32'd92,32'd5830,32'd514,32'd886,32'd-653,32'd-10703,32'd4848,32'd-1315,32'd-129,32'd-731,32'd538,32'd-2302,32'd-7631,32'd-2890,32'd-936,32'd3081,32'd-292,32'd237,32'd1867,32'd1160,32'd-633,32'd-5712,32'd885,32'd338,32'd5507,32'd1256,32'd-2312,32'd847,32'd-3432,32'd4960,32'd1068,32'd5292,32'd-7099,32'd1589,32'd1977,32'd192,32'd149,32'd-266,32'd3322,32'd-1960,32'd-624,32'd-1811,32'd-1365,32'd514,32'd1499,32'd1239,32'd453,32'd351,32'd2690,32'd2634,32'd-566,32'd-1669,32'd-2919,32'd6787,32'd1571,32'd1883,32'd2131,32'd-3666,32'd4782,32'd2727,32'd-944,32'd-568,32'd1809,32'd1271,32'd3178,32'd-2048,32'd1597,32'd382,32'd-4013,32'd2714,32'd-1395,32'd-1591,32'd-3361,32'd-4624,32'd3742,32'd1341,32'd-2442,32'd-536,32'd-4384,32'd4123,32'd-5698,32'd3833,32'd848,32'd-2047,32'd-3662,32'd-586,32'd318,32'd486,32'd510,32'd2420,32'd-1080,32'd428,32'd-4624,32'd-778,32'd-2296,32'd-1702,32'd2442,32'd1352,32'd-1871,32'd598,32'd-3642,32'd-1323,32'd-1542,32'd1358,32'd-7558,32'd-2038,32'd-1533,32'd1926,32'd-2416,32'd-7104,32'd-1466,32'd-2393,32'd-2070,32'd-73,32'd5390,32'd1572,32'd-4064,32'd-3105,32'd5654,32'd576,32'd2010,32'd-4357,32'd1052,32'd1627,32'd357,32'd-178,32'd-833,32'd3237,32'd-238,32'd-5185,32'd-3620,32'd4375,32'd-869,32'd6542,32'd96,32'd946,32'd-3764,32'd-6230,32'd-2810,32'd2705,32'd-1367,32'd-5405,32'd2895,32'd1138,32'd-1300,32'd-2526,32'd1546,32'd5034,32'd-753,32'd1256,32'd2081,32'd-2354,32'd-9272,32'd-4367,32'd4301,32'd-2854,32'd2153,32'd889,32'd3947,32'd-1016,32'd4904,32'd-1268,32'd298,32'd10029,32'd-1811,32'd724,32'd2570,32'd4714,32'd4291,32'd-1013,32'd-546,32'd-2575,32'd-1057,32'd-4875,32'd-838,32'd-6240,32'd-869,32'd2042,32'd-3193,32'd-1645,32'd-4382,32'd2521,32'd-33,32'd-30,32'd-1966,32'd3830,32'd-1602,32'd5898,32'd-6625,32'd-4912,32'd-3481,32'd-3098,32'd-678,32'd1846,32'd4072,32'd-1696,32'd-7299,32'd-933,32'd315,32'd3232,32'd-2607,32'd-3723,32'd-1019,32'd556,32'd-6923,32'd2210,32'd-3283,32'd729,32'd-2016,32'd4182,32'd-415,32'd2653,32'd-4235,32'd-233,32'd-6,32'd1230,32'd-757};
    Wh[22]='{32'd1689,32'd550,32'd-933,32'd4160,32'd-120,32'd-799,32'd5444,32'd2768,32'd270,32'd-171,32'd1372,32'd7592,32'd737,32'd1856,32'd-3129,32'd-2054,32'd1534,32'd-187,32'd2761,32'd1884,32'd-1009,32'd2661,32'd-694,32'd-1347,32'd-924,32'd-390,32'd-1595,32'd44,32'd2602,32'd-540,32'd509,32'd10302,32'd-2792,32'd1997,32'd1552,32'd-4089,32'd-1678,32'd5375,32'd2225,32'd-731,32'd4326,32'd910,32'd-5112,32'd-572,32'd3317,32'd4162,32'd5825,32'd8427,32'd1557,32'd-1732,32'd2558,32'd2233,32'd-2634,32'd-957,32'd-1608,32'd-2399,32'd-5605,32'd2286,32'd2597,32'd189,32'd3122,32'd1960,32'd206,32'd-1589,32'd-1502,32'd158,32'd-2026,32'd-551,32'd-803,32'd-559,32'd-2797,32'd3986,32'd1330,32'd2398,32'd-3618,32'd6958,32'd1076,32'd1066,32'd-3684,32'd6889,32'd-802,32'd-2839,32'd-2086,32'd5087,32'd-6391,32'd559,32'd913,32'd-293,32'd3012,32'd-965,32'd-1022,32'd-1301,32'd4345,32'd-688,32'd4206,32'd-999,32'd-2056,32'd327,32'd2949,32'd-17,32'd2639,32'd-1612,32'd1611,32'd6645,32'd-1297,32'd-2800,32'd1607,32'd-599,32'd136,32'd-142,32'd484,32'd-2548,32'd-6401,32'd2083,32'd59,32'd-1021,32'd-2156,32'd2459,32'd1416,32'd-905,32'd-1462,32'd-2048,32'd-6040,32'd7392,32'd881,32'd-2127,32'd-1252,32'd841,32'd1334,32'd1453,32'd4633,32'd-754,32'd-166,32'd-802,32'd-4455,32'd-1629,32'd-9760,32'd2249,32'd-2568,32'd-62,32'd895,32'd-51,32'd4165,32'd-1011,32'd-1350,32'd-388,32'd-1927,32'd90,32'd770,32'd-1325,32'd-957,32'd123,32'd-1511,32'd2047,32'd3232,32'd-1154,32'd-282,32'd2210,32'd-1036,32'd-195,32'd-7456,32'd-1356,32'd1833,32'd-2294,32'd-4716,32'd4035,32'd2456,32'd-532,32'd-223,32'd-726,32'd6518,32'd-2858,32'd729,32'd4306,32'd-2731,32'd120,32'd-3735,32'd-1669,32'd1333,32'd-1405,32'd-734,32'd702,32'd4340,32'd-1616,32'd-2362,32'd-7241,32'd5083,32'd963,32'd-3369,32'd-1174,32'd1076,32'd-2486,32'd1233,32'd-2382,32'd-1343,32'd-5458,32'd-4228,32'd538,32'd-298,32'd-1386,32'd831,32'd-2121,32'd-862,32'd4680,32'd-1614,32'd-1275,32'd996,32'd-1435,32'd165,32'd2753,32'd3879,32'd2858,32'd-269,32'd-1024,32'd2519,32'd1054,32'd1623,32'd-1109,32'd3742,32'd1683,32'd-2109,32'd5502,32'd2017,32'd-2766,32'd3100,32'd2059,32'd2719,32'd-2298,32'd1676,32'd2629,32'd3886,32'd-558,32'd5966,32'd-941,32'd916,32'd-929,32'd-695,32'd222,32'd4194,32'd-283,32'd489,32'd-1481,32'd643,32'd-6171,32'd-562,32'd1613,32'd2358,32'd-4396,32'd1489,32'd842,32'd1413,32'd-1578,32'd-531,32'd-1593,32'd1949,32'd2264,32'd960,32'd-509,32'd-725,32'd6342,32'd-3449,32'd-2431,32'd-5639,32'd2456,32'd2067,32'd-1896,32'd2082,32'd2343,32'd-1412,32'd-3293,32'd4787,32'd-3422,32'd932,32'd4309,32'd-398,32'd-9267,32'd-1235,32'd-4443,32'd2059,32'd4594,32'd-2008,32'd1341,32'd4277,32'd2663,32'd246,32'd1119,32'd-384,32'd4992,32'd1491,32'd-366,32'd10,32'd-994,32'd1146,32'd-2337,32'd515,32'd6250,32'd708,32'd-878,32'd-347,32'd-597,32'd-1314,32'd-8085,32'd150,32'd2651,32'd-560,32'd-295,32'd4477,32'd3937,32'd-1052,32'd3664,32'd-4169,32'd-2910,32'd-2434,32'd-2489,32'd-3479,32'd1256,32'd-5063,32'd1132,32'd1412,32'd3830,32'd6723,32'd5429,32'd-2700,32'd-3215,32'd334,32'd1407,32'd1850,32'd-1517,32'd-1398,32'd-1048,32'd355,32'd-228,32'd3012,32'd-2443,32'd-2539,32'd-2863,32'd6577,32'd7890,32'd-1481,32'd5239,32'd20,32'd4470,32'd1517,32'd5478,32'd86,32'd-679,32'd-1540,32'd-30,32'd2128,32'd1409,32'd2766,32'd445,32'd1678,32'd-5146,32'd-2373,32'd3544,32'd-140,32'd3205,32'd373,32'd1320,32'd2707,32'd4384,32'd503,32'd133,32'd-6118,32'd4194,32'd1246,32'd3549,32'd1773,32'd1868,32'd1722,32'd-2834,32'd-2841,32'd2858,32'd-2106,32'd3403,32'd-1220,32'd-3178,32'd2287,32'd311,32'd3466,32'd3393,32'd7807,32'd-1773,32'd-6059,32'd2514,32'd6250,32'd2137,32'd2185,32'd-3298,32'd-241,32'd2729,32'd1687,32'd-3579,32'd1052,32'd4221,32'd-76,32'd-892,32'd8149,32'd-1372};
    Wh[23]='{32'd2824,32'd1776,32'd1765,32'd-4050,32'd414,32'd-2800,32'd5068,32'd-4,32'd1783,32'd-1641,32'd1015,32'd3476,32'd-1402,32'd-525,32'd4211,32'd-2060,32'd5732,32'd4553,32'd2196,32'd741,32'd-70,32'd2159,32'd-5385,32'd-3122,32'd980,32'd-4023,32'd-2077,32'd-721,32'd-1679,32'd3498,32'd2156,32'd2171,32'd1766,32'd2541,32'd-1459,32'd-4809,32'd662,32'd-1934,32'd2922,32'd6894,32'd4057,32'd1557,32'd-1015,32'd3417,32'd469,32'd-1047,32'd48,32'd-816,32'd2524,32'd-2722,32'd-2531,32'd2583,32'd-5732,32'd-1124,32'd431,32'd4040,32'd2700,32'd1669,32'd4091,32'd6367,32'd2440,32'd-166,32'd6821,32'd515,32'd-770,32'd2878,32'd-4865,32'd1813,32'd2954,32'd2590,32'd373,32'd2670,32'd3833,32'd4377,32'd-1196,32'd927,32'd2343,32'd1793,32'd354,32'd-3808,32'd1047,32'd-4138,32'd-1069,32'd2712,32'd1909,32'd1530,32'd-492,32'd-1265,32'd252,32'd478,32'd2731,32'd-1221,32'd725,32'd2717,32'd1329,32'd-3327,32'd2310,32'd-1762,32'd339,32'd2751,32'd-2241,32'd4538,32'd1624,32'd3054,32'd569,32'd91,32'd6005,32'd7,32'd6738,32'd-225,32'd-3969,32'd-1586,32'd-140,32'd7900,32'd527,32'd143,32'd-2445,32'd619,32'd3933,32'd-4814,32'd-605,32'd-1706,32'd-5532,32'd-1975,32'd-656,32'd-8911,32'd5063,32'd803,32'd1378,32'd-11093,32'd-1324,32'd2366,32'd-1993,32'd-3303,32'd-3979,32'd-4050,32'd3881,32'd-78,32'd383,32'd1633,32'd-4904,32'd2551,32'd1000,32'd-804,32'd3261,32'd-4396,32'd1021,32'd-3513,32'd2585,32'd1867,32'd-1340,32'd2474,32'd624,32'd-92,32'd1420,32'd425,32'd7153,32'd2298,32'd1190,32'd-5922,32'd1992,32'd-4614,32'd459,32'd-8007,32'd6196,32'd1816,32'd1032,32'd-493,32'd352,32'd1939,32'd-651,32'd2078,32'd-352,32'd1666,32'd2043,32'd-3505,32'd-1958,32'd2861,32'd-4477,32'd1772,32'd-1695,32'd-5366,32'd5214,32'd-3273,32'd3220,32'd-709,32'd-136,32'd-1232,32'd-3334,32'd2465,32'd-4807,32'd-1146,32'd-4528,32'd2795,32'd-3479,32'd-2164,32'd-2985,32'd-291,32'd5527,32'd239,32'd-3774,32'd1564,32'd1433,32'd-2215,32'd-928,32'd-1568,32'd444,32'd2219,32'd1217,32'd666,32'd-3815,32'd1656,32'd523,32'd-1300,32'd-791,32'd4174,32'd-2780,32'd3168,32'd970,32'd-787,32'd2077,32'd2954,32'd6679,32'd6381,32'd532,32'd1738,32'd3176,32'd312,32'd-3486,32'd3669,32'd-1051,32'd-4421,32'd1892,32'd-527,32'd6123,32'd4416,32'd905,32'd-2448,32'd828,32'd1944,32'd7622,32'd-2790,32'd722,32'd325,32'd-1254,32'd1026,32'd4272,32'd-847,32'd1370,32'd-42,32'd-1118,32'd2954,32'd-2244,32'd-1206,32'd-488,32'd1119,32'd5502,32'd-110,32'd5590,32'd715,32'd1385,32'd3037,32'd623,32'd-4291,32'd-6484,32'd2337,32'd-2069,32'd-62,32'd872,32'd1221,32'd-2500,32'd1336,32'd4165,32'd893,32'd-5468,32'd-6889,32'd3615,32'd1859,32'd-1101,32'd1168,32'd2529,32'd308,32'd-6376,32'd2290,32'd68,32'd1354,32'd-1856,32'd5400,32'd-3164,32'd693,32'd6542,32'd233,32'd74,32'd2612,32'd2770,32'd3935,32'd6508,32'd5844,32'd-2946,32'd-3041,32'd-438,32'd-397,32'd5224,32'd-3129,32'd3198,32'd7309,32'd196,32'd-1812,32'd1396,32'd669,32'd4106,32'd1484,32'd2502,32'd2454,32'd-1326,32'd5180,32'd1420,32'd3054,32'd-81,32'd3166,32'd3833,32'd1411,32'd2790,32'd4047,32'd1176,32'd-369,32'd8989,32'd-1116,32'd-92,32'd509,32'd4960,32'd1545,32'd1705,32'd-1903,32'd6298,32'd8417,32'd-2231,32'd1660,32'd-4042,32'd-4997,32'd2235,32'd972,32'd-3872,32'd1243,32'd4025,32'd3403,32'd-10781,32'd-1882,32'd-148,32'd-957,32'd-493,32'd952,32'd-2250,32'd573,32'd1762,32'd-2829,32'd6791,32'd2968,32'd4772,32'd-907,32'd-2600,32'd2739,32'd1459,32'd-2714,32'd-4987,32'd12314,32'd-3415,32'd-5048,32'd411,32'd2937,32'd-1162,32'd-51,32'd2202,32'd4729,32'd-5561,32'd2066,32'd-4150,32'd1832,32'd2408,32'd5278,32'd6987,32'd-386,32'd-2873,32'd85,32'd2364,32'd1156,32'd-96,32'd6738,32'd3103,32'd61,32'd698,32'd-4770,32'd6723,32'd-2042,32'd1497,32'd-3522,32'd6479,32'd2810,32'd9570,32'd346};
    Wh[24]='{32'd-942,32'd2512,32'd771,32'd-1721,32'd2481,32'd-1436,32'd2556,32'd-4997,32'd7177,32'd3352,32'd-415,32'd188,32'd1139,32'd-3745,32'd4541,32'd3935,32'd224,32'd1478,32'd-1524,32'd407,32'd-1323,32'd983,32'd-1829,32'd1766,32'd1508,32'd-247,32'd-2824,32'd2517,32'd-1163,32'd-1950,32'd-2042,32'd-781,32'd478,32'd-707,32'd892,32'd3276,32'd2937,32'd2219,32'd-5688,32'd88,32'd-1253,32'd-1484,32'd-10205,32'd4255,32'd-4533,32'd-2380,32'd-2458,32'd1291,32'd-1055,32'd-3493,32'd1987,32'd-3183,32'd-3022,32'd-6542,32'd3095,32'd-2081,32'd7226,32'd-3024,32'd650,32'd7729,32'd-1437,32'd1612,32'd-1940,32'd4489,32'd5439,32'd-1248,32'd-2807,32'd181,32'd855,32'd1333,32'd-2915,32'd975,32'd-4519,32'd413,32'd1842,32'd-403,32'd667,32'd786,32'd420,32'd-217,32'd3708,32'd512,32'd-3300,32'd1718,32'd-612,32'd350,32'd112,32'd419,32'd1341,32'd-318,32'd2778,32'd3481,32'd490,32'd-1281,32'd-2380,32'd1300,32'd377,32'd1002,32'd2458,32'd-354,32'd-344,32'd29,32'd2135,32'd-537,32'd-3923,32'd149,32'd-2390,32'd-4379,32'd2440,32'd-900,32'd-211,32'd1634,32'd2354,32'd-3859,32'd2011,32'd-1386,32'd-679,32'd3215,32'd8720,32'd3457,32'd-3740,32'd809,32'd2514,32'd3937,32'd-2121,32'd-2629,32'd1339,32'd-1551,32'd3952,32'd-1629,32'd652,32'd3046,32'd-1317,32'd4326,32'd-1920,32'd4853,32'd7861,32'd-1429,32'd-3342,32'd-2308,32'd386,32'd-731,32'd-1211,32'd-188,32'd390,32'd-1572,32'd-2832,32'd-8139,32'd-409,32'd3999,32'd2332,32'd-1503,32'd6909,32'd3557,32'd158,32'd-566,32'd-5708,32'd958,32'd-6806,32'd-1652,32'd-1386,32'd-1423,32'd-2741,32'd7070,32'd-1590,32'd-1156,32'd4172,32'd3527,32'd3007,32'd-523,32'd5312,32'd-2315,32'd-1099,32'd-2502,32'd-1003,32'd52,32'd2130,32'd-264,32'd-2753,32'd489,32'd-4189,32'd-406,32'd835,32'd2072,32'd-1385,32'd-2551,32'd-3481,32'd-461,32'd1784,32'd-1027,32'd-1077,32'd-3161,32'd-2282,32'd1406,32'd-534,32'd4978,32'd5097,32'd4218,32'd-144,32'd-2436,32'd-2272,32'd-969,32'd2539,32'd1619,32'd2130,32'd-1055,32'd1567,32'd2578,32'd-2663,32'd2172,32'd2836,32'd7768,32'd-438,32'd1418,32'd558,32'd-2492,32'd-1964,32'd3254,32'd-996,32'd-1947,32'd-375,32'd1004,32'd1900,32'd700,32'd-147,32'd-1856,32'd4033,32'd-483,32'd3876,32'd-1474,32'd1328,32'd-10009,32'd1213,32'd677,32'd5844,32'd-392,32'd-4208,32'd-955,32'd2336,32'd5859,32'd2841,32'd-3491,32'd-2185,32'd3371,32'd1785,32'd1270,32'd2025,32'd0,32'd3857,32'd-5429,32'd-3947,32'd3698,32'd-4831,32'd4829,32'd8403,32'd5361,32'd1865,32'd-4780,32'd2802,32'd-1418,32'd187,32'd2104,32'd2172,32'd2673,32'd-7407,32'd4340,32'd561,32'd2614,32'd1376,32'd107,32'd-1932,32'd3894,32'd-2207,32'd1914,32'd-1097,32'd-2993,32'd8754,32'd-561,32'd1345,32'd1075,32'd5175,32'd-501,32'd3784,32'd-3796,32'd1920,32'd4091,32'd2016,32'd3547,32'd-5654,32'd5927,32'd4204,32'd237,32'd-268,32'd-881,32'd-3059,32'd2685,32'd-1715,32'd167,32'd144,32'd2224,32'd-1531,32'd-1801,32'd5004,32'd139,32'd3134,32'd100,32'd4489,32'd-1739,32'd947,32'd2832,32'd789,32'd-334,32'd295,32'd-187,32'd147,32'd-784,32'd419,32'd2558,32'd-1385,32'd988,32'd4042,32'd-1269,32'd-2247,32'd-375,32'd4931,32'd1295,32'd1506,32'd663,32'd-2180,32'd-499,32'd569,32'd-308,32'd266,32'd53,32'd-2912,32'd205,32'd506,32'd-3251,32'd4458,32'd1806,32'd3986,32'd1068,32'd-927,32'd209,32'd-3425,32'd1392,32'd4025,32'd4184,32'd-3461,32'd-556,32'd2639,32'd-2352,32'd-191,32'd2419,32'd652,32'd2929,32'd2125,32'd1436,32'd-155,32'd-3698,32'd437,32'd-343,32'd1295,32'd6791,32'd3706,32'd4152,32'd-7080,32'd3710,32'd1632,32'd2185,32'd-6254,32'd302,32'd4204,32'd647,32'd-1142,32'd-1270,32'd-477,32'd-1106,32'd2595,32'd3078,32'd5532,32'd-1469,32'd2283,32'd-1542,32'd5698,32'd-3015,32'd2102,32'd2849,32'd1039,32'd1727,32'd3520,32'd-2292,32'd3566,32'd-10507,32'd-7470,32'd3896,32'd-83,32'd1595,32'd6743,32'd-632};
    Wh[25]='{32'd-64,32'd-494,32'd-1726,32'd38,32'd-1181,32'd473,32'd187,32'd1046,32'd-3044,32'd798,32'd-3015,32'd4372,32'd3845,32'd-3063,32'd2727,32'd2573,32'd-3476,32'd415,32'd-4309,32'd825,32'd1301,32'd-2856,32'd1649,32'd1132,32'd3466,32'd3032,32'd-5825,32'd-3330,32'd393,32'd-1430,32'd3356,32'd-4860,32'd-991,32'd1209,32'd-2814,32'd186,32'd123,32'd2683,32'd-785,32'd-3051,32'd-6538,32'd-1080,32'd1017,32'd-4638,32'd-1623,32'd-5048,32'd-54,32'd-2739,32'd-1297,32'd4562,32'd-2341,32'd2895,32'd5185,32'd5327,32'd-1823,32'd-6079,32'd3054,32'd-388,32'd1873,32'd1135,32'd-365,32'd-4418,32'd-180,32'd330,32'd-376,32'd-2509,32'd3193,32'd1082,32'd-1667,32'd-6562,32'd-6000,32'd-2705,32'd-5952,32'd1652,32'd1810,32'd5458,32'd2047,32'd2298,32'd-2130,32'd-1129,32'd-1083,32'd1222,32'd-1938,32'd1270,32'd3754,32'd2158,32'd574,32'd-5541,32'd-47,32'd4125,32'd-2839,32'd-6782,32'd4301,32'd-4643,32'd-1804,32'd2001,32'd-296,32'd-967,32'd-2291,32'd-2810,32'd-1067,32'd-5268,32'd822,32'd-8100,32'd-1027,32'd-196,32'd2583,32'd-698,32'd13164,32'd-4858,32'd250,32'd4228,32'd4338,32'd-2692,32'd-2264,32'd-2634,32'd-1879,32'd3618,32'd-1481,32'd-235,32'd574,32'd502,32'd2668,32'd-2053,32'd-1556,32'd-6088,32'd5185,32'd-1572,32'd6206,32'd2286,32'd960,32'd-348,32'd-2128,32'd-2651,32'd1066,32'd-433,32'd5712,32'd-5917,32'd-1966,32'd170,32'd6079,32'd-333,32'd-2100,32'd-1260,32'd830,32'd1625,32'd-1002,32'd-121,32'd3488,32'd2612,32'd-303,32'd-3447,32'd-3439,32'd5776,32'd-4240,32'd-3972,32'd-2103,32'd723,32'd-3481,32'd1542,32'd2399,32'd758,32'd715,32'd902,32'd-3715,32'd-4777,32'd-377,32'd-3176,32'd-3212,32'd779,32'd1376,32'd776,32'd-4633,32'd1005,32'd1992,32'd4704,32'd1441,32'd238,32'd853,32'd-562,32'd-2670,32'd-1802,32'd-1395,32'd2526,32'd-3110,32'd2137,32'd-4726,32'd3017,32'd2474,32'd-4379,32'd-2322,32'd-823,32'd7773,32'd2092,32'd1923,32'd4396,32'd317,32'd387,32'd-3906,32'd3237,32'd-392,32'd-805,32'd328,32'd-139,32'd4960,32'd-396,32'd-2919,32'd-3818,32'd-4267,32'd-6186,32'd44,32'd-839,32'd-1024,32'd-1636,32'd225,32'd2482,32'd-3767,32'd-3356,32'd-1138,32'd-1691,32'd-2966,32'd23,32'd-3359,32'd-1577,32'd-1580,32'd-2697,32'd-2272,32'd470,32'd2939,32'd626,32'd3554,32'd451,32'd-1190,32'd-1297,32'd-3925,32'd3081,32'd911,32'd-5327,32'd2729,32'd-1781,32'd-229,32'd240,32'd-47,32'd947,32'd2587,32'd311,32'd-4367,32'd-4768,32'd-361,32'd-1025,32'd1756,32'd-2349,32'd563,32'd-4353,32'd-1143,32'd-132,32'd-1149,32'd-2773,32'd-1402,32'd-2347,32'd949,32'd3747,32'd-2464,32'd4023,32'd-552,32'd376,32'd3229,32'd-2866,32'd308,32'd2558,32'd4365,32'd-1094,32'd-795,32'd-543,32'd2014,32'd7050,32'd-3215,32'd2927,32'd-55,32'd-2521,32'd-3967,32'd-969,32'd-1293,32'd1229,32'd-1054,32'd-5239,32'd-1635,32'd-5756,32'd424,32'd2357,32'd-2614,32'd-1529,32'd-37,32'd15,32'd-2492,32'd1291,32'd1131,32'd137,32'd-2744,32'd4523,32'd-1734,32'd631,32'd-745,32'd-1273,32'd3769,32'd-3061,32'd-2158,32'd-447,32'd-1551,32'd-5771,32'd-504,32'd-1015,32'd1340,32'd2958,32'd-3891,32'd374,32'd-8652,32'd-232,32'd-2033,32'd5493,32'd-209,32'd-203,32'd-3479,32'd-1459,32'd-5668,32'd-948,32'd-2310,32'd-3205,32'd4567,32'd-4057,32'd2432,32'd591,32'd1586,32'd1883,32'd-6318,32'd-193,32'd887,32'd-2373,32'd4072,32'd4470,32'd-988,32'd-2314,32'd3850,32'd-6933,32'd-1627,32'd-1302,32'd-63,32'd3610,32'd3359,32'd1102,32'd-2749,32'd5517,32'd-1740,32'd374,32'd-4555,32'd3325,32'd764,32'd2010,32'd1374,32'd2315,32'd-405,32'd-4497,32'd2102,32'd3564,32'd1573,32'd2878,32'd631,32'd-191,32'd1430,32'd-4440,32'd-2197,32'd-5561,32'd-1112,32'd1489,32'd2661,32'd-2441,32'd5043,32'd1472,32'd-3793,32'd-1768,32'd-4160,32'd-1679,32'd-1995,32'd-1711,32'd-3894,32'd-2291,32'd-2849,32'd-4963,32'd-3581,32'd-3452,32'd1140,32'd1776,32'd-786,32'd-823,32'd4094,32'd1077,32'd1337,32'd-911,32'd91,32'd143};
    Wh[26]='{32'd-913,32'd6176,32'd2734,32'd-1777,32'd2149,32'd-1712,32'd-430,32'd-1312,32'd-1325,32'd-939,32'd2014,32'd-730,32'd2034,32'd1665,32'd-3662,32'd-473,32'd905,32'd3312,32'd2144,32'd-788,32'd-242,32'd3920,32'd-1934,32'd807,32'd-487,32'd-23,32'd3347,32'd-2304,32'd5634,32'd-8261,32'd-1876,32'd-2966,32'd-2071,32'd3833,32'd4130,32'd-1138,32'd2128,32'd328,32'd137,32'd1096,32'd37,32'd3122,32'd-2158,32'd1148,32'd533,32'd-68,32'd2318,32'd1274,32'd-3239,32'd2000,32'd1840,32'd-1406,32'd-3200,32'd-2861,32'd-1800,32'd2539,32'd3144,32'd-5937,32'd-4272,32'd4211,32'd241,32'd-6733,32'd852,32'd-384,32'd3330,32'd-18,32'd-375,32'd-602,32'd2639,32'd1293,32'd2148,32'd-1291,32'd-2846,32'd-2084,32'd2673,32'd-1827,32'd2746,32'd1750,32'd1713,32'd-1225,32'd-156,32'd-1510,32'd3078,32'd1078,32'd-1727,32'd-2834,32'd940,32'd-2239,32'd-252,32'd-326,32'd2905,32'd-120,32'd-1237,32'd-3149,32'd-1183,32'd2196,32'd-467,32'd-595,32'd1060,32'd-1507,32'd-1892,32'd462,32'd1479,32'd-1850,32'd2985,32'd-244,32'd3164,32'd-3859,32'd4577,32'd-2602,32'd-1038,32'd3371,32'd-7797,32'd-3820,32'd4797,32'd-1611,32'd6303,32'd8852,32'd4055,32'd-1950,32'd716,32'd5302,32'd-4797,32'd1340,32'd1516,32'd-91,32'd-7905,32'd2966,32'd-3896,32'd-2352,32'd-1183,32'd3730,32'd-1246,32'd493,32'd38,32'd1470,32'd4855,32'd1102,32'd-337,32'd-5185,32'd-1748,32'd1069,32'd-3823,32'd2595,32'd-29,32'd-13,32'd2061,32'd322,32'd-2288,32'd1879,32'd4602,32'd-693,32'd-3957,32'd-1230,32'd986,32'd-7231,32'd-3898,32'd3081,32'd-3205,32'd-2442,32'd-9184,32'd-1419,32'd-3955,32'd3547,32'd2644,32'd3012,32'd-2419,32'd-1706,32'd687,32'd-2719,32'd-1319,32'd5048,32'd-4687,32'd1036,32'd3723,32'd1900,32'd5195,32'd-2362,32'd368,32'd-3183,32'd130,32'd3107,32'd-2758,32'd521,32'd-3579,32'd-320,32'd-4006,32'd-3566,32'd-3920,32'd2448,32'd789,32'd-3732,32'd2536,32'd-2749,32'd872,32'd3835,32'd-541,32'd-2318,32'd7324,32'd-386,32'd-1556,32'd2907,32'd-1851,32'd263,32'd772,32'd-849,32'd239,32'd-1889,32'd440,32'd239,32'd-5268,32'd-1112,32'd-1478,32'd939,32'd925,32'd1205,32'd-611,32'd-905,32'd-5908,32'd-5893,32'd1394,32'd1354,32'd2175,32'd1871,32'd-4699,32'd-2398,32'd-3039,32'd645,32'd1357,32'd2247,32'd-314,32'd1414,32'd-4423,32'd-1203,32'd-492,32'd2778,32'd2106,32'd-1483,32'd-1582,32'd130,32'd-4191,32'd2410,32'd-6577,32'd-2890,32'd65,32'd281,32'd-7451,32'd-2412,32'd-3681,32'd-4299,32'd-1240,32'd-2692,32'd1663,32'd-4865,32'd-3454,32'd-5400,32'd-605,32'd1013,32'd1156,32'd542,32'd372,32'd2486,32'd-1447,32'd-2492,32'd-3010,32'd-628,32'd1148,32'd517,32'd880,32'd-2561,32'd-3767,32'd179,32'd-2100,32'd3435,32'd-5776,32'd-1682,32'd859,32'd-559,32'd1181,32'd212,32'd3430,32'd-4472,32'd-2836,32'd-3115,32'd581,32'd-1890,32'd-2113,32'd1959,32'd-656,32'd-5371,32'd3759,32'd600,32'd-6284,32'd-2130,32'd62,32'd-709,32'd-3999,32'd-2083,32'd-9741,32'd-2834,32'd2044,32'd326,32'd-4101,32'd1672,32'd1437,32'd809,32'd881,32'd-1595,32'd3496,32'd2009,32'd-1212,32'd-473,32'd-556,32'd-2088,32'd-2834,32'd-3420,32'd902,32'd-328,32'd-1354,32'd7451,32'd20,32'd-4702,32'd-2604,32'd475,32'd-374,32'd565,32'd9008,32'd466,32'd-6015,32'd-834,32'd-807,32'd2753,32'd-3132,32'd-2587,32'd334,32'd3515,32'd-1373,32'd-5629,32'd-1030,32'd1928,32'd2036,32'd-5708,32'd1549,32'd1362,32'd-917,32'd1367,32'd3752,32'd-4841,32'd-969,32'd-3664,32'd-1428,32'd-3361,32'd1427,32'd535,32'd-1842,32'd-3774,32'd-3249,32'd5810,32'd833,32'd-2208,32'd1614,32'd-1865,32'd-3798,32'd1101,32'd1247,32'd-3862,32'd-560,32'd9057,32'd2270,32'd2110,32'd-177,32'd-494,32'd-2788,32'd498,32'd985,32'd-1364,32'd2534,32'd1781,32'd2220,32'd-3188,32'd-1333,32'd2153,32'd-2717,32'd2264,32'd1807,32'd-3505,32'd-1115,32'd4587,32'd1933,32'd-2008,32'd3459,32'd5434,32'd-5688,32'd3662,32'd-191,32'd816,32'd6455,32'd-3041,32'd8374,32'd-1425};
    Wh[27]='{32'd-648,32'd2390,32'd1024,32'd-643,32'd1619,32'd-969,32'd-5517,32'd-4270,32'd42,32'd2335,32'd-497,32'd-321,32'd1280,32'd387,32'd4313,32'd-4350,32'd-817,32'd-3317,32'd-1868,32'd-1706,32'd1350,32'd-3798,32'd-876,32'd1176,32'd2578,32'd551,32'd-508,32'd-1008,32'd-1871,32'd3007,32'd2,32'd-947,32'd-851,32'd-1545,32'd4416,32'd1884,32'd1944,32'd825,32'd-1625,32'd-3020,32'd2531,32'd4409,32'd-1726,32'd3833,32'd3750,32'd880,32'd-5234,32'd612,32'd-304,32'd-2885,32'd-350,32'd4567,32'd-3068,32'd-2163,32'd-3125,32'd-586,32'd2666,32'd-578,32'd-1085,32'd-2185,32'd-2995,32'd1650,32'd832,32'd1671,32'd-425,32'd-3293,32'd-233,32'd1711,32'd1180,32'd-359,32'd-1942,32'd918,32'd-907,32'd-776,32'd2849,32'd3229,32'd-1222,32'd-6059,32'd-497,32'd-4050,32'd-2058,32'd2761,32'd-1215,32'd3505,32'd446,32'd1772,32'd1555,32'd-2553,32'd-2746,32'd-1412,32'd1477,32'd1119,32'd-888,32'd781,32'd-3996,32'd-17,32'd-1469,32'd-2435,32'd2001,32'd757,32'd-1594,32'd-2196,32'd-775,32'd-1058,32'd-614,32'd494,32'd783,32'd-5629,32'd1616,32'd750,32'd237,32'd621,32'd231,32'd1551,32'd-1728,32'd-1707,32'd-2009,32'd-4130,32'd4313,32'd-25,32'd-837,32'd-444,32'd-1066,32'd2924,32'd-376,32'd-1888,32'd4328,32'd-1716,32'd-95,32'd-6489,32'd-345,32'd2495,32'd-615,32'd232,32'd-4956,32'd-1657,32'd2587,32'd-1202,32'd4509,32'd1146,32'd2814,32'd1837,32'd-1755,32'd-4079,32'd218,32'd1739,32'd-2340,32'd564,32'd2238,32'd-3225,32'd3242,32'd594,32'd-2297,32'd-2993,32'd1368,32'd3017,32'd2003,32'd-513,32'd2006,32'd-2800,32'd1936,32'd45,32'd-2497,32'd-599,32'd-1918,32'd154,32'd699,32'd1756,32'd899,32'd-665,32'd67,32'd2214,32'd-2054,32'd-4382,32'd138,32'd1105,32'd2189,32'd1016,32'd-2641,32'd669,32'd-2487,32'd-3625,32'd-1024,32'd4978,32'd62,32'd3312,32'd3212,32'd3286,32'd1783,32'd-3288,32'd2695,32'd1813,32'd3630,32'd-5522,32'd-3645,32'd-2202,32'd-3601,32'd626,32'd-5537,32'd2016,32'd3513,32'd-4741,32'd156,32'd-1967,32'd1172,32'd394,32'd3278,32'd-3125,32'd-3632,32'd1370,32'd5068,32'd1031,32'd2239,32'd-2440,32'd2384,32'd-254,32'd-2253,32'd2172,32'd2856,32'd-4711,32'd1627,32'd699,32'd1983,32'd453,32'd-1177,32'd3710,32'd1614,32'd182,32'd1520,32'd4062,32'd1273,32'd-5590,32'd1540,32'd-993,32'd-9599,32'd-3205,32'd-313,32'd81,32'd-2429,32'd-203,32'd1098,32'd-7187,32'd2052,32'd-4890,32'd-3063,32'd1083,32'd-2810,32'd-1071,32'd4104,32'd3977,32'd3315,32'd4152,32'd-1282,32'd3823,32'd-5732,32'd-2478,32'd993,32'd1446,32'd3059,32'd3276,32'd1017,32'd2749,32'd1291,32'd-1942,32'd-1209,32'd2463,32'd1228,32'd-2141,32'd-921,32'd-546,32'd3701,32'd4321,32'd410,32'd-673,32'd596,32'd53,32'd2797,32'd3730,32'd6088,32'd-1480,32'd-158,32'd-4133,32'd-907,32'd-881,32'd-87,32'd3090,32'd614,32'd314,32'd6191,32'd3259,32'd2995,32'd1599,32'd2364,32'd-1600,32'd-3376,32'd-3256,32'd-2553,32'd1918,32'd1527,32'd1224,32'd2,32'd1490,32'd2834,32'd1536,32'd957,32'd2739,32'd2015,32'd-4184,32'd-2487,32'd5317,32'd-819,32'd-476,32'd4001,32'd821,32'd2292,32'd2194,32'd-579,32'd-4687,32'd1716,32'd721,32'd996,32'd-999,32'd54,32'd-1447,32'd-1683,32'd-2230,32'd362,32'd5288,32'd809,32'd-321,32'd2895,32'd4453,32'd1171,32'd4301,32'd655,32'd3483,32'd-2497,32'd291,32'd2871,32'd5375,32'd3430,32'd2917,32'd-3686,32'd-8120,32'd238,32'd5004,32'd-1084,32'd1447,32'd5747,32'd-265,32'd-2512,32'd1610,32'd637,32'd1538,32'd-668,32'd-603,32'd523,32'd9589,32'd2617,32'd377,32'd189,32'd4838,32'd1702,32'd1296,32'd97,32'd-2414,32'd4387,32'd4042,32'd4821,32'd4343,32'd-6489,32'd4340,32'd4250,32'd2093,32'd2910,32'd704,32'd1201,32'd-648,32'd2291,32'd1083,32'd-155,32'd-100,32'd593,32'd3615,32'd2680,32'd149,32'd566,32'd-339,32'd3190,32'd-1503,32'd650,32'd2199,32'd783,32'd-7475,32'd-883,32'd1459,32'd-1734,32'd1684,32'd2191,32'd1264};
    Wh[28]='{32'd-1152,32'd1925,32'd-1087,32'd3854,32'd-2073,32'd1480,32'd10009,32'd-2333,32'd4963,32'd-2003,32'd6044,32'd-4870,32'd2692,32'd2680,32'd3623,32'd5429,32'd-2192,32'd-2426,32'd4055,32'd4040,32'd3835,32'd455,32'd805,32'd-186,32'd2993,32'd3156,32'd6694,32'd-731,32'd9360,32'd1702,32'd2595,32'd-69,32'd1406,32'd173,32'd-3125,32'd3664,32'd-5585,32'd1501,32'd-3186,32'd-2048,32'd7182,32'd3469,32'd1773,32'd-330,32'd-1093,32'd-429,32'd5170,32'd-2602,32'd4406,32'd-3994,32'd7192,32'd-2512,32'd-1242,32'd-5727,32'd2059,32'd1098,32'd-4062,32'd1237,32'd2543,32'd-3508,32'd-5595,32'd-4130,32'd3310,32'd277,32'd1333,32'd4895,32'd-2479,32'd-1624,32'd-3237,32'd-1403,32'd3662,32'd4499,32'd-1340,32'd1704,32'd597,32'd-2043,32'd-1326,32'd5312,32'd3847,32'd1896,32'd1778,32'd4001,32'd3298,32'd382,32'd380,32'd-1843,32'd2135,32'd4111,32'd2973,32'd287,32'd-935,32'd-5009,32'd-4399,32'd-4572,32'd4826,32'd2609,32'd4274,32'd-483,32'd5678,32'd-1445,32'd-17,32'd3691,32'd1108,32'd-3349,32'd2531,32'd-800,32'd2053,32'd3286,32'd-7734,32'd-3535,32'd-6196,32'd-2561,32'd-2961,32'd-894,32'd-2651,32'd-837,32'd748,32'd5073,32'd-2597,32'd2839,32'd650,32'd-164,32'd7651,32'd4826,32'd-7202,32'd-6157,32'd1144,32'd-948,32'd-11074,32'd1531,32'd10917,32'd2514,32'd-1514,32'd-2327,32'd2048,32'd-3725,32'd-722,32'd-3325,32'd-5073,32'd1302,32'd-3911,32'd557,32'd4592,32'd-580,32'd979,32'd-4301,32'd5278,32'd-9511,32'd-3476,32'd-5156,32'd498,32'd3813,32'd-2712,32'd-3156,32'd6909,32'd1633,32'd-3171,32'd-1303,32'd-2145,32'd6704,32'd-2597,32'd3081,32'd1166,32'd8730,32'd-3386,32'd-5356,32'd3403,32'd2126,32'd432,32'd-1089,32'd-573,32'd-1098,32'd-6899,32'd1796,32'd2120,32'd-2343,32'd-1499,32'd2160,32'd-2446,32'd2985,32'd726,32'd196,32'd529,32'd7509,32'd-1318,32'd3300,32'd2473,32'd2249,32'd-9345,32'd114,32'd-974,32'd-287,32'd10849,32'd-2272,32'd1243,32'd3400,32'd1468,32'd20,32'd1940,32'd4038,32'd-852,32'd3820,32'd1405,32'd-6,32'd3525,32'd2680,32'd304,32'd3520,32'd-1771,32'd1948,32'd-2646,32'd379,32'd2014,32'd1613,32'd5024,32'd3503,32'd6367,32'd2468,32'd5048,32'd3598,32'd2133,32'd-1374,32'd4426,32'd-2222,32'd1528,32'd-494,32'd1466,32'd1987,32'd-7851,32'd-369,32'd4187,32'd2580,32'd3608,32'd2644,32'd3227,32'd-1890,32'd-4645,32'd2418,32'd685,32'd-1934,32'd-5893,32'd4204,32'd-296,32'd147,32'd-4340,32'd918,32'd-2215,32'd-4606,32'd5307,32'd-3476,32'd2531,32'd-1922,32'd3024,32'd-3503,32'd-2272,32'd527,32'd5449,32'd-5771,32'd1842,32'd3239,32'd1883,32'd1997,32'd273,32'd1586,32'd2687,32'd6645,32'd-212,32'd2052,32'd791,32'd-2797,32'd2072,32'd-6669,32'd947,32'd-392,32'd-5053,32'd3188,32'd-3977,32'd2846,32'd4570,32'd3107,32'd-430,32'd-1384,32'd4902,32'd-2377,32'd5957,32'd-1008,32'd3403,32'd722,32'd-1857,32'd-2673,32'd567,32'd-3740,32'd-1881,32'd-1665,32'd2067,32'd9516,32'd-7817,32'd-2308,32'd2409,32'd4404,32'd-4301,32'd6284,32'd-1849,32'd459,32'd-299,32'd-3181,32'd11298,32'd449,32'd3464,32'd-13,32'd-1433,32'd-1057,32'd11191,32'd-3947,32'd578,32'd-6313,32'd-1578,32'd-1602,32'd11640,32'd14677,32'd-2016,32'd-166,32'd-2722,32'd1453,32'd3342,32'd89,32'd-4470,32'd-3588,32'd1375,32'd3015,32'd3181,32'd-3122,32'd1293,32'd-3718,32'd-6367,32'd3249,32'd1169,32'd-728,32'd8784,32'd-1022,32'd1694,32'd-7651,32'd-4882,32'd-3554,32'd1290,32'd3354,32'd6347,32'd3666,32'd1403,32'd-3520,32'd-143,32'd2401,32'd-2629,32'd-3156,32'd-1691,32'd4821,32'd-1135,32'd-1444,32'd4123,32'd1506,32'd2792,32'd6293,32'd232,32'd512,32'd2375,32'd-4372,32'd-5732,32'd1950,32'd657,32'd-6289,32'd-3881,32'd2807,32'd-2580,32'd-1340,32'd816,32'd5913,32'd2995,32'd929,32'd-1336,32'd2163,32'd-1112,32'd2176,32'd4838,32'd-7661,32'd-3615,32'd-3659,32'd1666,32'd2128,32'd921,32'd-1632,32'd-1523,32'd2425,32'd755,32'd-3020,32'd3535,32'd1214,32'd-440,32'd1475,32'd2814,32'd-277};
    Wh[29]='{32'd-936,32'd5561,32'd1749,32'd2658,32'd-318,32'd-3571,32'd-1483,32'd-21,32'd528,32'd401,32'd8593,32'd2302,32'd7368,32'd2370,32'd-2320,32'd4426,32'd3981,32'd802,32'd400,32'd-2983,32'd-1540,32'd-6689,32'd4160,32'd7089,32'd90,32'd-1341,32'd2504,32'd-3120,32'd245,32'd-3771,32'd-3913,32'd-1202,32'd3696,32'd811,32'd-2587,32'd-1114,32'd-4719,32'd1524,32'd-2741,32'd1445,32'd-3508,32'd-5986,32'd1759,32'd-1795,32'd-2683,32'd-1302,32'd8676,32'd-3649,32'd-2248,32'd4367,32'd-5146,32'd2812,32'd-2249,32'd-1560,32'd-591,32'd-690,32'd3930,32'd-13007,32'd2978,32'd-1798,32'd-1875,32'd-5234,32'd3481,32'd-1280,32'd4462,32'd-1878,32'd2902,32'd1085,32'd-2954,32'd-154,32'd-6596,32'd-5781,32'd-411,32'd-2580,32'd-888,32'd5097,32'd-855,32'd-1627,32'd-5952,32'd1907,32'd552,32'd-8364,32'd5644,32'd2152,32'd348,32'd-436,32'd-589,32'd-563,32'd-3122,32'd-15263,32'd-117,32'd-217,32'd-154,32'd-2990,32'd123,32'd1900,32'd398,32'd3691,32'd777,32'd316,32'd-3317,32'd338,32'd1912,32'd15712,32'd-2279,32'd-2482,32'd2392,32'd3872,32'd772,32'd576,32'd2880,32'd-7636,32'd6420,32'd-620,32'd3012,32'd1043,32'd-4140,32'd257,32'd2512,32'd225,32'd-2934,32'd-9189,32'd-3598,32'd-2502,32'd681,32'd16250,32'd-3037,32'd-1903,32'd878,32'd-6005,32'd-12724,32'd605,32'd-9086,32'd-69,32'd3732,32'd10068,32'd-5639,32'd-4331,32'd4938,32'd1467,32'd-4533,32'd785,32'd723,32'd-1093,32'd2922,32'd2272,32'd-717,32'd4582,32'd4804,32'd-6611,32'd-1171,32'd3103,32'd-2922,32'd3063,32'd-2993,32'd1333,32'd-195,32'd3662,32'd-4118,32'd2320,32'd1557,32'd-484,32'd1696,32'd4921,32'd3312,32'd-28,32'd3498,32'd2639,32'd3610,32'd316,32'd-4218,32'd-2790,32'd616,32'd-121,32'd-8403,32'd-654,32'd968,32'd6567,32'd5498,32'd2451,32'd1811,32'd5361,32'd-1461,32'd-3107,32'd3134,32'd3466,32'd5371,32'd1975,32'd1132,32'd-5698,32'd806,32'd-285,32'd-5854,32'd-539,32'd6484,32'd-5004,32'd-64,32'd499,32'd5205,32'd-603,32'd-814,32'd1337,32'd-867,32'd-6562,32'd-1844,32'd-2763,32'd408,32'd4851,32'd-1252,32'd-1633,32'd-1257,32'd-372,32'd-10605,32'd975,32'd3000,32'd850,32'd-961,32'd-73,32'd-2480,32'd-2902,32'd1668,32'd3410,32'd-5834,32'd-1595,32'd2407,32'd-3659,32'd-4926,32'd-820,32'd-3059,32'd-5966,32'd-9018,32'd-1045,32'd4414,32'd-5014,32'd-3015,32'd1352,32'd-1302,32'd1932,32'd1218,32'd723,32'd-292,32'd1770,32'd-527,32'd-5883,32'd1132,32'd38,32'd4599,32'd-3400,32'd831,32'd1848,32'd-1765,32'd-3105,32'd1518,32'd-5297,32'd-6733,32'd671,32'd1835,32'd-9775,32'd1945,32'd-3325,32'd-9746,32'd11,32'd847,32'd-2294,32'd3476,32'd714,32'd-473,32'd-2137,32'd1342,32'd-4421,32'd-4362,32'd-3520,32'd-357,32'd-609,32'd1185,32'd-7202,32'd265,32'd-3476,32'd1240,32'd-1776,32'd618,32'd3977,32'd6132,32'd-5683,32'd-2575,32'd-10556,32'd-739,32'd-1527,32'd-3937,32'd1697,32'd-6899,32'd-4138,32'd231,32'd626,32'd-158,32'd1168,32'd1708,32'd-9658,32'd559,32'd271,32'd-1979,32'd-10996,32'd2282,32'd-791,32'd-760,32'd-2578,32'd3618,32'd-2963,32'd-3371,32'd-2293,32'd-3234,32'd-3444,32'd-4355,32'd2028,32'd-7768,32'd-1414,32'd11337,32'd-909,32'd4582,32'd6396,32'd-69,32'd5585,32'd-5195,32'd-1795,32'd237,32'd1878,32'd1462,32'd-1427,32'd-1748,32'd-933,32'd-5634,32'd2325,32'd-4926,32'd-9360,32'd-359,32'd4003,32'd-635,32'd-4934,32'd-1319,32'd204,32'd1295,32'd2362,32'd4069,32'd1853,32'd6254,32'd-2634,32'd1403,32'd-7495,32'd-1752,32'd3125,32'd6586,32'd-2279,32'd-6,32'd3769,32'd-1095,32'd1953,32'd2932,32'd-5458,32'd-1120,32'd5366,32'd-3515,32'd4301,32'd-2424,32'd-3562,32'd-6049,32'd-6757,32'd-732,32'd-4226,32'd-2932,32'd1362,32'd985,32'd58,32'd-4567,32'd1823,32'd-2673,32'd-51,32'd-1711,32'd-358,32'd-600,32'd-1911,32'd-3652,32'd1271,32'd2082,32'd-2391,32'd2419,32'd2078,32'd948,32'd-513,32'd-1027,32'd3327,32'd-7060,32'd4814,32'd-5991,32'd963,32'd-8666,32'd3535,32'd2587,32'd241,32'd2150,32'd-5634};
    Wh[30]='{32'd2841,32'd-913,32'd228,32'd2937,32'd2810,32'd-2393,32'd1484,32'd-4790,32'd-1542,32'd-287,32'd1950,32'd2257,32'd-2170,32'd1286,32'd4855,32'd-682,32'd-2958,32'd-429,32'd1789,32'd1782,32'd1739,32'd-2401,32'd-6767,32'd-574,32'd2001,32'd1456,32'd3376,32'd-748,32'd1100,32'd-2047,32'd-2271,32'd6118,32'd36,32'd1350,32'd-1784,32'd1456,32'd905,32'd-1291,32'd1049,32'd3598,32'd-147,32'd-713,32'd-3068,32'd877,32'd-3581,32'd1004,32'd2795,32'd-1290,32'd745,32'd-4479,32'd-3249,32'd2941,32'd-4335,32'd-2963,32'd-935,32'd4978,32'd-1428,32'd2736,32'd-3745,32'd-555,32'd2736,32'd551,32'd-2321,32'd1907,32'd5698,32'd1071,32'd245,32'd1166,32'd-1976,32'd357,32'd3498,32'd-229,32'd3442,32'd-1578,32'd2111,32'd-830,32'd3796,32'd1617,32'd-4294,32'd-551,32'd456,32'd-530,32'd-2064,32'd-1234,32'd-4533,32'd854,32'd3513,32'd779,32'd3920,32'd1832,32'd1086,32'd-282,32'd4228,32'd-97,32'd-1099,32'd514,32'd-710,32'd3937,32'd-1523,32'd2169,32'd-1960,32'd1330,32'd-1529,32'd13427,32'd4011,32'd336,32'd-1412,32'd-1855,32'd3129,32'd5151,32'd-4423,32'd-1693,32'd-1868,32'd5615,32'd948,32'd4343,32'd-2717,32'd1556,32'd-1820,32'd-3566,32'd-1959,32'd-287,32'd1909,32'd-5976,32'd746,32'd-2541,32'd-4396,32'd1439,32'd-3015,32'd3989,32'd-7382,32'd764,32'd-1398,32'd-3928,32'd-5302,32'd-6708,32'd-2360,32'd3569,32'd-3776,32'd375,32'd-2546,32'd1306,32'd-3925,32'd2327,32'd7207,32'd-4365,32'd2539,32'd-3674,32'd-234,32'd2968,32'd-1790,32'd-3674,32'd-751,32'd1658,32'd6523,32'd5537,32'd-3762,32'd-411,32'd-1027,32'd-637,32'd886,32'd2183,32'd-12,32'd-7822,32'd-1782,32'd5400,32'd-1640,32'd-3547,32'd1851,32'd-981,32'd43,32'd-1434,32'd7905,32'd1000,32'd-527,32'd1149,32'd-5571,32'd47,32'd1296,32'd-2714,32'd-814,32'd3630,32'd-1431,32'd-2509,32'd-953,32'd949,32'd1861,32'd5937,32'd-4882,32'd-1215,32'd-1116,32'd2705,32'd1669,32'd-3457,32'd-2286,32'd-2546,32'd2308,32'd-2666,32'd-1402,32'd-7075,32'd1066,32'd493,32'd1333,32'd-1597,32'd-637,32'd-39,32'd-561,32'd5922,32'd-2005,32'd2836,32'd4401,32'd3442,32'd2371,32'd-2370,32'd2147,32'd884,32'd579,32'd1500,32'd2775,32'd2292,32'd2194,32'd5146,32'd3281,32'd-2003,32'd3225,32'd-1077,32'd736,32'd497,32'd2675,32'd442,32'd-485,32'd2406,32'd3132,32'd2376,32'd-470,32'd1111,32'd-1181,32'd462,32'd-123,32'd3789,32'd3166,32'd2600,32'd3942,32'd18,32'd-2751,32'd957,32'd3823,32'd-5332,32'd646,32'd439,32'd-777,32'd1074,32'd822,32'd5786,32'd-2678,32'd613,32'd-431,32'd1876,32'd1804,32'd5937,32'd5776,32'd-4277,32'd-4489,32'd-616,32'd-1400,32'd2476,32'd25,32'd3552,32'd-914,32'd-1085,32'd2492,32'd2783,32'd-419,32'd819,32'd1627,32'd223,32'd-442,32'd2093,32'd-31,32'd3789,32'd1489,32'd616,32'd-2152,32'd-3425,32'd2484,32'd3381,32'd800,32'd2966,32'd-137,32'd-1691,32'd2692,32'd-6450,32'd4028,32'd1419,32'd-665,32'd5058,32'd-393,32'd692,32'd-14,32'd-2363,32'd3305,32'd690,32'd4604,32'd4716,32'd2373,32'd4482,32'd-141,32'd-487,32'd505,32'd-914,32'd-1623,32'd1914,32'd75,32'd-4421,32'd316,32'd4514,32'd6616,32'd-1314,32'd-152,32'd-2617,32'd3825,32'd632,32'd-3950,32'd-1711,32'd4660,32'd2829,32'd-1722,32'd1392,32'd465,32'd127,32'd-2272,32'd1423,32'd-180,32'd4050,32'd-135,32'd2587,32'd4035,32'd-22,32'd-250,32'd2326,32'd2434,32'd2314,32'd-2403,32'd-755,32'd1729,32'd2062,32'd2531,32'd-797,32'd2200,32'd-717,32'd7495,32'd753,32'd1761,32'd-978,32'd-1702,32'd731,32'd475,32'd1822,32'd-1704,32'd3352,32'd8505,32'd2130,32'd-1146,32'd-1695,32'd-2180,32'd-524,32'd1562,32'd-162,32'd-1835,32'd-1057,32'd4975,32'd1342,32'd-55,32'd421,32'd4914,32'd2773,32'd-218,32'd-1157,32'd-653,32'd1326,32'd2946,32'd359,32'd-733,32'd3876,32'd-2670,32'd-2636,32'd5952,32'd3693,32'd1235,32'd-2670,32'd233,32'd-3603,32'd807,32'd3793,32'd-1730,32'd4838,32'd-4177,32'd1403,32'd406,32'd-1301};
    Wh[31]='{32'd539,32'd-75,32'd-380,32'd-2418,32'd94,32'd-226,32'd149,32'd9624,32'd-2604,32'd-4133,32'd2220,32'd542,32'd1148,32'd-1866,32'd-2122,32'd-1556,32'd1905,32'd11,32'd655,32'd3796,32'd-242,32'd-1456,32'd-1267,32'd-4123,32'd-1196,32'd1150,32'd4909,32'd3117,32'd93,32'd1767,32'd722,32'd-7895,32'd701,32'd309,32'd2277,32'd1662,32'd-2387,32'd852,32'd1315,32'd2592,32'd5664,32'd405,32'd-2766,32'd2983,32'd199,32'd725,32'd-2739,32'd3825,32'd-888,32'd1553,32'd1135,32'd3803,32'd2734,32'd3376,32'd1651,32'd4868,32'd1328,32'd-208,32'd-1611,32'd5419,32'd1617,32'd-345,32'd2254,32'd3903,32'd3037,32'd2137,32'd-6826,32'd-4020,32'd2231,32'd2320,32'd-5200,32'd8481,32'd-1021,32'd4260,32'd-5039,32'd7714,32'd841,32'd3264,32'd-608,32'd2324,32'd-247,32'd2561,32'd8789,32'd-5869,32'd-5122,32'd5092,32'd-3283,32'd-2213,32'd-1152,32'd2573,32'd-244,32'd5991,32'd4157,32'd664,32'd3317,32'd3117,32'd-1005,32'd-2047,32'd164,32'd-3576,32'd-2431,32'd-6250,32'd791,32'd-154,32'd-2807,32'd555,32'd-3784,32'd-3991,32'd-1447,32'd-3808,32'd-2968,32'd10253,32'd-5815,32'd-2895,32'd-946,32'd-3764,32'd616,32'd5595,32'd8925,32'd-2447,32'd3112,32'd7343,32'd-2382,32'd6757,32'd7939,32'd-7807,32'd7705,32'd-26,32'd-6293,32'd-2269,32'd1713,32'd6206,32'd-5263,32'd3793,32'd306,32'd-4538,32'd474,32'd2517,32'd-4821,32'd4157,32'd-1004,32'd404,32'd-3449,32'd-4189,32'd-3732,32'd1241,32'd252,32'd993,32'd4648,32'd-2807,32'd-1966,32'd-4953,32'd-3557,32'd-866,32'd-4108,32'd-6074,32'd4367,32'd-415,32'd67,32'd-11083,32'd-4162,32'd1357,32'd-2770,32'd717,32'd715,32'd10224,32'd3845,32'd6025,32'd-1813,32'd1673,32'd-1859,32'd2456,32'd-258,32'd2266,32'd-4638,32'd-3166,32'd-1790,32'd-3176,32'd-4353,32'd1656,32'd3793,32'd-6918,32'd1166,32'd-1413,32'd-5136,32'd-1862,32'd5283,32'd329,32'd3051,32'd3859,32'd-1761,32'd-5537,32'd-5395,32'd-2663,32'd-1348,32'd4804,32'd-1705,32'd-4211,32'd909,32'd206,32'd18,32'd-3239,32'd1761,32'd-3022,32'd-5517,32'd957,32'd484,32'd408,32'd2225,32'd-3828,32'd-4770,32'd-3950,32'd-651,32'd6411,32'd-1239,32'd-885,32'd-1308,32'd3881,32'd-92,32'd-339,32'd5068,32'd5839,32'd-4411,32'd-1771,32'd-1988,32'd2282,32'd-4780,32'd4453,32'd3232,32'd-2351,32'd-2304,32'd-1182,32'd-5478,32'd-1646,32'd3955,32'd1176,32'd-2307,32'd-1748,32'd-3103,32'd-1113,32'd833,32'd115,32'd-3698,32'd1639,32'd-1759,32'd1691,32'd-1566,32'd-5297,32'd-3818,32'd-1087,32'd-4042,32'd2690,32'd1840,32'd-4025,32'd-1428,32'd941,32'd602,32'd-2368,32'd-2658,32'd-3537,32'd1169,32'd-353,32'd7070,32'd-3640,32'd3220,32'd-2976,32'd-1072,32'd1212,32'd-730,32'd1264,32'd10,32'd-1883,32'd-747,32'd-4047,32'd1211,32'd3149,32'd1202,32'd-7895,32'd2023,32'd2010,32'd3234,32'd-1424,32'd1793,32'd4665,32'd-4265,32'd-3559,32'd3320,32'd254,32'd58,32'd1018,32'd4902,32'd-812,32'd3251,32'd-2673,32'd-230,32'd-5102,32'd3222,32'd4226,32'd-2453,32'd-761,32'd1401,32'd4172,32'd1336,32'd4741,32'd878,32'd6845,32'd2858,32'd4885,32'd1451,32'd116,32'd-1259,32'd-4438,32'd-3071,32'd-2427,32'd1503,32'd-296,32'd-489,32'd-4003,32'd6694,32'd3935,32'd3095,32'd-806,32'd-138,32'd-5942,32'd1375,32'd-5405,32'd-1636,32'd2104,32'd1159,32'd597,32'd-7207,32'd4643,32'd2958,32'd-1050,32'd78,32'd-2132,32'd-3413,32'd5214,32'd-5366,32'd-3688,32'd-960,32'd-3249,32'd1188,32'd5253,32'd1555,32'd4497,32'd-2917,32'd-3239,32'd-4323,32'd-21,32'd5000,32'd3825,32'd-781,32'd-5341,32'd-2563,32'd1392,32'd-7001,32'd-2307,32'd7148,32'd-3750,32'd1323,32'd761,32'd3129,32'd412,32'd-2136,32'd-2464,32'd-3515,32'd-634,32'd3911,32'd-3930,32'd-497,32'd-4030,32'd4909,32'd681,32'd-2185,32'd-3020,32'd6669,32'd-2614,32'd4704,32'd4362,32'd6518,32'd-5546,32'd5307,32'd2460,32'd3061,32'd5146,32'd38,32'd5883,32'd-280,32'd10322,32'd3283,32'd1042,32'd-6440,32'd-482,32'd3806,32'd529,32'd-2069,32'd-54,32'd-2362,32'd-1672};
    Wh[32]='{32'd-2254,32'd-9633,32'd-1667,32'd-3422,32'd1873,32'd-1373,32'd772,32'd-6318,32'd5107,32'd40,32'd-3620,32'd-3527,32'd-7890,32'd3659,32'd434,32'd4008,32'd2807,32'd-574,32'd-3225,32'd-1120,32'd935,32'd1166,32'd-222,32'd1320,32'd-506,32'd-3088,32'd-112,32'd-657,32'd-10244,32'd-802,32'd-2875,32'd-5727,32'd-2880,32'd-1596,32'd3681,32'd-2277,32'd605,32'd-1353,32'd-4235,32'd963,32'd-10537,32'd-1495,32'd-9594,32'd-5488,32'd-4587,32'd6010,32'd-2998,32'd-2573,32'd2717,32'd555,32'd7290,32'd-793,32'd-4399,32'd-2783,32'd-958,32'd-3395,32'd-2602,32'd-787,32'd-6240,32'd2749,32'd-414,32'd-5419,32'd-313,32'd-3188,32'd-2702,32'd1743,32'd-2373,32'd-3342,32'd-4692,32'd-5024,32'd1510,32'd-1442,32'd-5966,32'd1379,32'd-3598,32'd-5766,32'd4606,32'd-4914,32'd4348,32'd1857,32'd-218,32'd-2200,32'd-1267,32'd480,32'd-407,32'd-839,32'd-2702,32'd3515,32'd-3828,32'd1984,32'd-2775,32'd-1990,32'd-10175,32'd1496,32'd-2609,32'd-1243,32'd-1251,32'd1708,32'd206,32'd-7617,32'd2474,32'd5585,32'd303,32'd2880,32'd1403,32'd3049,32'd5092,32'd5146,32'd2727,32'd-1483,32'd-4064,32'd5820,32'd13310,32'd-3818,32'd-4580,32'd1973,32'd1450,32'd10849,32'd5068,32'd12,32'd3256,32'd3173,32'd-72,32'd4289,32'd5639,32'd-8432,32'd6953,32'd-677,32'd5771,32'd-2756,32'd-2729,32'd-1000,32'd-6044,32'd5673,32'd4230,32'd-6176,32'd-316,32'd3137,32'd2377,32'd3281,32'd123,32'd-1625,32'd-687,32'd132,32'd-1165,32'd-3847,32'd3654,32'd2283,32'd-4809,32'd3347,32'd-2048,32'd-1017,32'd2255,32'd-5258,32'd1938,32'd-16103,32'd3049,32'd-603,32'd6440,32'd-25097,32'd12089,32'd2846,32'd232,32'd3676,32'd2469,32'd-13076,32'd-4694,32'd-552,32'd3784,32'd-482,32'd-659,32'd1279,32'd-8217,32'd2072,32'd1518,32'd1342,32'd-507,32'd889,32'd498,32'd-2147,32'd5786,32'd-2546,32'd-1247,32'd20,32'd2626,32'd-253,32'd-2893,32'd7065,32'd11572,32'd2687,32'd3093,32'd-764,32'd8750,32'd329,32'd1049,32'd-935,32'd2553,32'd145,32'd-45,32'd-150,32'd3786,32'd575,32'd1138,32'd4191,32'd-2631,32'd-253,32'd3969,32'd-2512,32'd674,32'd6977,32'd-3945,32'd1201,32'd5668,32'd2822,32'd7182,32'd5483,32'd5922,32'd2844,32'd-1198,32'd3681,32'd682,32'd221,32'd-1412,32'd1563,32'd2489,32'd2736,32'd-5854,32'd1065,32'd3166,32'd772,32'd-2846,32'd2812,32'd4704,32'd979,32'd-708,32'd6757,32'd-1744,32'd-314,32'd-6660,32'd1228,32'd6142,32'd-257,32'd-744,32'd-9023,32'd9125,32'd4558,32'd629,32'd3417,32'd-6567,32'd-1077,32'd-669,32'd1571,32'd3906,32'd4714,32'd3750,32'd2580,32'd996,32'd2435,32'd-4038,32'd-8564,32'd-1237,32'd5249,32'd1058,32'd569,32'd867,32'd-553,32'd1953,32'd-2463,32'd-2420,32'd678,32'd357,32'd9047,32'd-2580,32'd-41,32'd-1489,32'd-276,32'd4125,32'd1845,32'd3168,32'd-368,32'd1757,32'd1390,32'd-446,32'd6250,32'd-1334,32'd2556,32'd-4504,32'd583,32'd2998,32'd3312,32'd-1839,32'd4145,32'd-2286,32'd2827,32'd1491,32'd-796,32'd-6333,32'd1661,32'd-3615,32'd3891,32'd5649,32'd2849,32'd-2678,32'd7866,32'd1418,32'd-10898,32'd-2299,32'd-2126,32'd-701,32'd-2056,32'd-6264,32'd-4736,32'd4516,32'd9746,32'd-6191,32'd2541,32'd3525,32'd-2410,32'd-9897,32'd3190,32'd-2858,32'd2636,32'd-2954,32'd947,32'd1251,32'd2434,32'd-5053,32'd-2250,32'd-4477,32'd-1943,32'd-734,32'd-629,32'd1171,32'd3754,32'd3710,32'd13935,32'd980,32'd-7895,32'd-2453,32'd5458,32'd-3554,32'd868,32'd1004,32'd-3527,32'd-676,32'd4602,32'd495,32'd3874,32'd-16113,32'd-148,32'd5117,32'd-1025,32'd-1614,32'd-1337,32'd3666,32'd-900,32'd-3803,32'd2556,32'd-6748,32'd-857,32'd6733,32'd-2044,32'd3291,32'd1890,32'd3095,32'd-196,32'd-4516,32'd1468,32'd111,32'd-1268,32'd-350,32'd2150,32'd-10048,32'd3732,32'd5034,32'd-3095,32'd1995,32'd1052,32'd-86,32'd1473,32'd668,32'd7548,32'd-4035,32'd3657,32'd-3251,32'd-253,32'd-5117,32'd-2369,32'd1844,32'd-2846,32'd2164,32'd-4,32'd-7500,32'd798,32'd-6113,32'd-2102,32'd-5195,32'd9028,32'd3627,32'd3188};
    Wh[33]='{32'd717,32'd-8090,32'd-857,32'd-1063,32'd2651,32'd-261,32'd6816,32'd3991,32'd-2824,32'd-1931,32'd-1209,32'd-4699,32'd-3244,32'd-1467,32'd-2910,32'd3208,32'd-4694,32'd3498,32'd-317,32'd-2573,32'd926,32'd3002,32'd-1690,32'd-2056,32'd-1042,32'd-2902,32'd-2152,32'd1023,32'd-7866,32'd3967,32'd391,32'd-1594,32'd1396,32'd-3605,32'd-4741,32'd-687,32'd-248,32'd101,32'd-4523,32'd5058,32'd-303,32'd1402,32'd-5263,32'd-521,32'd4323,32'd3562,32'd3752,32'd7099,32'd-3000,32'd-2714,32'd2199,32'd5952,32'd-64,32'd-5947,32'd963,32'd3173,32'd115,32'd3232,32'd-247,32'd-12832,32'd1756,32'd-155,32'd-2330,32'd-1015,32'd-1097,32'd2115,32'd1628,32'd-3627,32'd4501,32'd-3757,32'd1959,32'd306,32'd2292,32'd-1171,32'd703,32'd3405,32'd-5000,32'd-1387,32'd4343,32'd-1749,32'd-1340,32'd2344,32'd3952,32'd-637,32'd5180,32'd1926,32'd-4541,32'd819,32'd2998,32'd245,32'd-462,32'd-2475,32'd2181,32'd-12539,32'd-2315,32'd1483,32'd-3168,32'd-2384,32'd2429,32'd1661,32'd1007,32'd1270,32'd-809,32'd-5351,32'd2990,32'd2242,32'd-59,32'd5244,32'd-8657,32'd5581,32'd3132,32'd8847,32'd-2003,32'd2575,32'd3657,32'd3078,32'd-3139,32'd-5092,32'd2386,32'd-3295,32'd2880,32'd626,32'd-5156,32'd-5180,32'd-3146,32'd-2471,32'd650,32'd231,32'd-6108,32'd1970,32'd1857,32'd3757,32'd2426,32'd-9028,32'd2641,32'd-1727,32'd-1601,32'd1527,32'd-3967,32'd-2045,32'd-4899,32'd1606,32'd-5024,32'd8198,32'd5205,32'd-1159,32'd-1751,32'd-689,32'd-1008,32'd-4433,32'd-1026,32'd190,32'd-4433,32'd-3786,32'd-1009,32'd-1657,32'd-2756,32'd-3105,32'd-5126,32'd-1525,32'd-12988,32'd-221,32'd-885,32'd-2751,32'd42,32'd6997,32'd769,32'd-5917,32'd-431,32'd1195,32'd2150,32'd2161,32'd1837,32'd-536,32'd1027,32'd-3122,32'd-3969,32'd-160,32'd1962,32'd-883,32'd3942,32'd-2381,32'd-2614,32'd540,32'd585,32'd-2551,32'd-4887,32'd5048,32'd-6982,32'd2475,32'd-1109,32'd157,32'd-483,32'd-3605,32'd5424,32'd-13427,32'd-622,32'd5708,32'd5781,32'd4384,32'd1339,32'd1503,32'd-2077,32'd-5488,32'd-6044,32'd492,32'd-61,32'd-257,32'd1384,32'd-1718,32'd-97,32'd-1756,32'd-6762,32'd8017,32'd-486,32'd448,32'd2143,32'd2531,32'd-613,32'd1264,32'd855,32'd2489,32'd-7680,32'd1560,32'd-2065,32'd-6440,32'd-2526,32'd-2844,32'd-6835,32'd133,32'd247,32'd5034,32'd1373,32'd93,32'd1386,32'd347,32'd2922,32'd-2071,32'd-3400,32'd3435,32'd-2912,32'd1290,32'd-1671,32'd6601,32'd1260,32'd962,32'd1732,32'd5522,32'd-3095,32'd1567,32'd-2849,32'd-2239,32'd-4226,32'd2578,32'd-428,32'd6093,32'd-6806,32'd1345,32'd-4877,32'd8427,32'd1992,32'd-506,32'd-2561,32'd-771,32'd5825,32'd-2443,32'd-640,32'd-3701,32'd-372,32'd-1462,32'd6953,32'd-3669,32'd733,32'd-5952,32'd1536,32'd-2078,32'd-4523,32'd2524,32'd-4340,32'd130,32'd-4138,32'd-1607,32'd-1900,32'd-3789,32'd-4760,32'd3532,32'd-3251,32'd-496,32'd-1994,32'd-2454,32'd-1921,32'd1198,32'd-6171,32'd-2268,32'd-2663,32'd4294,32'd268,32'd2429,32'd5488,32'd129,32'd5751,32'd-3708,32'd-4890,32'd-661,32'd-746,32'd-6445,32'd7299,32'd916,32'd435,32'd-421,32'd-3879,32'd-1779,32'd-5073,32'd5712,32'd-4660,32'd-250,32'd450,32'd1525,32'd-1569,32'd1220,32'd-8325,32'd3562,32'd562,32'd921,32'd5053,32'd-1805,32'd-1662,32'd-2719,32'd-1258,32'd4873,32'd5068,32'd2424,32'd6586,32'd-428,32'd-2182,32'd-8295,32'd1154,32'd720,32'd2022,32'd1039,32'd1938,32'd-5664,32'd18,32'd7,32'd179,32'd-6064,32'd9467,32'd108,32'd1960,32'd-223,32'd4252,32'd2156,32'd3544,32'd-4699,32'd4458,32'd-505,32'd-3383,32'd-424,32'd8178,32'd-245,32'd-2539,32'd-5947,32'd-324,32'd577,32'd4904,32'd-5092,32'd4938,32'd-4821,32'd-3000,32'd406,32'd-1849,32'd-2788,32'd2893,32'd-3586,32'd-53,32'd-6279,32'd5615,32'd-7436,32'd3242,32'd2419,32'd-1455,32'd-5996,32'd11816,32'd517,32'd-6323,32'd4179,32'd-2407,32'd1278,32'd1646,32'd4445,32'd2956,32'd4992,32'd2910,32'd-88,32'd1030,32'd4433,32'd-3989,32'd6596,32'd-1168,32'd1612};
    Wh[34]='{32'd-3029,32'd339,32'd415,32'd178,32'd717,32'd-122,32'd1199,32'd2863,32'd1738,32'd2692,32'd1136,32'd1916,32'd-4658,32'd1738,32'd2170,32'd-2829,32'd4169,32'd2624,32'd470,32'd2617,32'd3244,32'd-1595,32'd-1428,32'd-445,32'd-3376,32'd67,32'd-173,32'd-3193,32'd2368,32'd-5668,32'd2449,32'd1622,32'd1115,32'd-2995,32'd7207,32'd317,32'd-12773,32'd3664,32'd232,32'd5063,32'd792,32'd-1094,32'd9,32'd-516,32'd-4055,32'd2675,32'd-6762,32'd1462,32'd-1763,32'd587,32'd4833,32'd2492,32'd4450,32'd58,32'd6435,32'd-5693,32'd2067,32'd4187,32'd-1448,32'd1955,32'd2783,32'd-2309,32'd3730,32'd1069,32'd1623,32'd3669,32'd-3901,32'd4218,32'd-3298,32'd-3837,32'd6816,32'd1990,32'd1729,32'd-2272,32'd-1778,32'd8598,32'd-1005,32'd4238,32'd6586,32'd2683,32'd5688,32'd2651,32'd-1335,32'd5878,32'd565,32'd6806,32'd-3149,32'd1530,32'd-2927,32'd4116,32'd-833,32'd7651,32'd3447,32'd4218,32'd42,32'd-191,32'd-1295,32'd4372,32'd1403,32'd2133,32'd-1236,32'd1422,32'd5239,32'd1029,32'd-4677,32'd1762,32'd737,32'd6660,32'd-10712,32'd2086,32'd-1312,32'd2192,32'd1154,32'd4621,32'd-2026,32'd-2211,32'd923,32'd687,32'd3405,32'd-109,32'd717,32'd-2709,32'd-574,32'd1232,32'd-1320,32'd-7675,32'd1114,32'd-5566,32'd146,32'd-2233,32'd-1519,32'd-74,32'd3354,32'd897,32'd22675,32'd2147,32'd-9228,32'd6464,32'd-2785,32'd-43,32'd6406,32'd1959,32'd7465,32'd61,32'd-4279,32'd-5737,32'd-568,32'd-5087,32'd-2247,32'd2468,32'd-1586,32'd2558,32'd-2132,32'd4318,32'd-7182,32'd1776,32'd2023,32'd-1024,32'd1372,32'd5288,32'd-3205,32'd477,32'd3769,32'd5263,32'd714,32'd-5869,32'd2355,32'd-3806,32'd4267,32'd-2370,32'd9853,32'd16,32'd-6430,32'd-1235,32'd805,32'd360,32'd6684,32'd-3942,32'd2958,32'd-5229,32'd1392,32'd-1857,32'd963,32'd-1699,32'd267,32'd-1975,32'd1010,32'd-515,32'd-6708,32'd1571,32'd3073,32'd3603,32'd172,32'd539,32'd-476,32'd8002,32'd5341,32'd1470,32'd-1719,32'd-4868,32'd-3981,32'd-1450,32'd-412,32'd870,32'd787,32'd-1044,32'd-1229,32'd1796,32'd-1602,32'd4121,32'd-5756,32'd1101,32'd-4504,32'd-1821,32'd-2851,32'd3466,32'd2108,32'd-4199,32'd1427,32'd5014,32'd1226,32'd5219,32'd5219,32'd1054,32'd2153,32'd2479,32'd4792,32'd-596,32'd-4128,32'd1800,32'd507,32'd1892,32'd1578,32'd2624,32'd15458,32'd16767,32'd-865,32'd1450,32'd-273,32'd-2861,32'd-6259,32'd-118,32'd-2951,32'd2861,32'd1354,32'd3232,32'd3347,32'd-745,32'd-4333,32'd-2868,32'd-122,32'd797,32'd-3571,32'd-1851,32'd1611,32'd-11064,32'd-2271,32'd4636,32'd-1412,32'd-8256,32'd340,32'd-1796,32'd1379,32'd-1431,32'd4230,32'd8666,32'd-6152,32'd-2604,32'd808,32'd-2333,32'd-4077,32'd3107,32'd262,32'd1130,32'd-2369,32'd-1508,32'd394,32'd-2360,32'd-10742,32'd1100,32'd7011,32'd-5322,32'd-5502,32'd-1069,32'd-676,32'd-2683,32'd-4169,32'd-340,32'd3681,32'd2178,32'd938,32'd1718,32'd3803,32'd-2105,32'd-5141,32'd905,32'd393,32'd-728,32'd2529,32'd-4877,32'd-7749,32'd3864,32'd3901,32'd1658,32'd551,32'd-578,32'd422,32'd1531,32'd7319,32'd-2420,32'd-3469,32'd-1939,32'd4311,32'd3000,32'd237,32'd-10605,32'd9780,32'd4724,32'd6997,32'd1979,32'd-1367,32'd4689,32'd4304,32'd282,32'd1198,32'd1256,32'd3430,32'd-1275,32'd2145,32'd-2570,32'd-3139,32'd-4780,32'd2827,32'd-7480,32'd-5922,32'd5292,32'd1006,32'd994,32'd1610,32'd-3872,32'd-6782,32'd740,32'd-6127,32'd-6752,32'd-4455,32'd6723,32'd5258,32'd-778,32'd733,32'd-5830,32'd11064,32'd-245,32'd1234,32'd-3481,32'd-2526,32'd9072,32'd2082,32'd-2188,32'd-9091,32'd-1218,32'd-4750,32'd-402,32'd7705,32'd2436,32'd195,32'd-511,32'd3786,32'd2004,32'd781,32'd-3588,32'd2580,32'd-3598,32'd-692,32'd-4208,32'd3613,32'd-1578,32'd6918,32'd-2427,32'd-3305,32'd546,32'd56,32'd7871,32'd2324,32'd1336,32'd-3151,32'd4431,32'd-8212,32'd6826,32'd968,32'd4777,32'd-1539,32'd-4028,32'd4199,32'd-2364,32'd-10771,32'd6826,32'd-896,32'd-100,32'd-2174,32'd-1105};
    Wh[35]='{32'd-3591,32'd-3715,32'd-1462,32'd-1607,32'd-1612,32'd659,32'd-1298,32'd4685,32'd-3417,32'd-2731,32'd4160,32'd352,32'd-991,32'd-795,32'd-112,32'd953,32'd-4291,32'd767,32'd-2381,32'd4997,32'd-599,32'd3791,32'd346,32'd-768,32'd546,32'd-2034,32'd1171,32'd1133,32'd-2070,32'd152,32'd664,32'd1756,32'd-3620,32'd-550,32'd-1790,32'd-979,32'd-2434,32'd-1721,32'd-2341,32'd1445,32'd-4458,32'd1102,32'd1369,32'd1612,32'd4433,32'd-3505,32'd-2191,32'd98,32'd1402,32'd4294,32'd-3745,32'd-3630,32'd2226,32'd1155,32'd-498,32'd-3769,32'd-2841,32'd252,32'd101,32'd-8549,32'd-2946,32'd-2391,32'd292,32'd-1887,32'd1165,32'd377,32'd567,32'd-3803,32'd1296,32'd-2734,32'd4274,32'd3054,32'd-2283,32'd-2932,32'd-1034,32'd2819,32'd340,32'd-1809,32'd1466,32'd-1973,32'd-2661,32'd671,32'd1593,32'd1206,32'd638,32'd1619,32'd1950,32'd-2985,32'd-4033,32'd3908,32'd-5180,32'd-6459,32'd-2890,32'd1373,32'd-509,32'd4775,32'd-971,32'd4050,32'd1757,32'd-938,32'd3903,32'd-1667,32'd-2912,32'd-7763,32'd3745,32'd-186,32'd-4545,32'd-3974,32'd-4655,32'd-355,32'd1225,32'd3696,32'd5268,32'd2587,32'd-2073,32'd-4079,32'd2,32'd2144,32'd-3852,32'd-1373,32'd-2561,32'd4938,32'd7656,32'd177,32'd-5546,32'd-5957,32'd6757,32'd4035,32'd2866,32'd-1435,32'd8486,32'd-3103,32'd-1831,32'd-3833,32'd-2152,32'd2644,32'd7177,32'd-3249,32'd-286,32'd3176,32'd-1068,32'd2188,32'd-1420,32'd-1389,32'd1606,32'd1955,32'd8032,32'd0,32'd-204,32'd-1904,32'd5107,32'd1925,32'd5747,32'd-1289,32'd-3977,32'd2993,32'd-4233,32'd287,32'd-526,32'd-3085,32'd-4787,32'd2049,32'd502,32'd-141,32'd2790,32'd-6083,32'd-2105,32'd602,32'd-383,32'd1185,32'd-1417,32'd1137,32'd-8242,32'd-10,32'd-162,32'd-880,32'd803,32'd641,32'd982,32'd3981,32'd5976,32'd-1851,32'd-4211,32'd1997,32'd-566,32'd3872,32'd-2229,32'd1778,32'd807,32'd2071,32'd-5585,32'd-1348,32'd-693,32'd3679,32'd528,32'd3176,32'd148,32'd-9282,32'd7924,32'd5800,32'd3376,32'd-601,32'd1259,32'd5415,32'd-3771,32'd1472,32'd-1003,32'd-4455,32'd-9599,32'd-1496,32'd-2167,32'd-3764,32'd-2340,32'd3264,32'd-1025,32'd-5253,32'd3344,32'd-1489,32'd-1481,32'd-2897,32'd1951,32'd-1135,32'd-601,32'd4865,32'd-1091,32'd-2055,32'd1550,32'd189,32'd-3293,32'd1250,32'd255,32'd-2536,32'd-7500,32'd3886,32'd-3583,32'd881,32'd-429,32'd-97,32'd2536,32'd-1209,32'd-2568,32'd3203,32'd-6127,32'd-393,32'd-4323,32'd2634,32'd-5717,32'd-1572,32'd-544,32'd1687,32'd-4150,32'd1970,32'd-1838,32'd1063,32'd1953,32'd-2493,32'd973,32'd-2805,32'd-3288,32'd3391,32'd-713,32'd-2722,32'd-2458,32'd1739,32'd-4843,32'd-3027,32'd-944,32'd529,32'd-900,32'd-357,32'd-113,32'd-55,32'd-2524,32'd4384,32'd-2824,32'd217,32'd-1572,32'd-2069,32'd85,32'd-725,32'd1079,32'd-946,32'd-914,32'd2824,32'd-1124,32'd-3212,32'd4167,32'd-1547,32'd4660,32'd1546,32'd9741,32'd-1978,32'd-471,32'd1812,32'd2421,32'd-2573,32'd-4965,32'd-12,32'd3898,32'd-359,32'd1439,32'd-1195,32'd2086,32'd-2454,32'd-2338,32'd-3193,32'd339,32'd-9672,32'd-1019,32'd-3459,32'd4206,32'd-2941,32'd-3640,32'd858,32'd1183,32'd-3933,32'd3632,32'd508,32'd-4333,32'd511,32'd-18,32'd-1033,32'd-2670,32'd5195,32'd1569,32'd1700,32'd-500,32'd3010,32'd-648,32'd809,32'd-1875,32'd749,32'd-8,32'd-1178,32'd1106,32'd1882,32'd-960,32'd1090,32'd434,32'd2497,32'd-332,32'd-5576,32'd1594,32'd2440,32'd1078,32'd-3618,32'd4465,32'd-2298,32'd158,32'd3488,32'd-707,32'd-4057,32'd5166,32'd-3300,32'd1001,32'd2995,32'd-935,32'd1903,32'd803,32'd3649,32'd-803,32'd-938,32'd-2568,32'd-1522,32'd449,32'd-4538,32'd4504,32'd-540,32'd2856,32'd-955,32'd-3588,32'd-1822,32'd-7568,32'd5708,32'd-1311,32'd-7451,32'd3869,32'd-1445,32'd5087,32'd-1661,32'd322,32'd827,32'd-900,32'd-916,32'd-3974,32'd4350,32'd-1479,32'd-1239,32'd-3137,32'd-1799,32'd1683,32'd2690,32'd-1745,32'd-465,32'd9501,32'd-3354,32'd-2377,32'd-2995,32'd737,32'd-4853};
    Wh[36]='{32'd-516,32'd-556,32'd-1314,32'd-4350,32'd129,32'd1223,32'd5541,32'd-522,32'd-768,32'd-2680,32'd-4250,32'd-4724,32'd1738,32'd-1331,32'd-2418,32'd-866,32'd-2824,32'd241,32'd-4145,32'd-693,32'd-608,32'd291,32'd-4887,32'd-502,32'd-3801,32'd-1185,32'd422,32'd-2155,32'd-9296,32'd-3034,32'd4143,32'd-2568,32'd-2978,32'd2678,32'd-12958,32'd-919,32'd4218,32'd1364,32'd-5458,32'd-1328,32'd3969,32'd-1746,32'd239,32'd-5253,32'd635,32'd-2868,32'd-9741,32'd377,32'd-1341,32'd3596,32'd-2636,32'd-3398,32'd2426,32'd-1199,32'd2661,32'd1159,32'd1265,32'd2673,32'd-509,32'd8583,32'd261,32'd-3449,32'd-3354,32'd3464,32'd1611,32'd-3647,32'd3918,32'd-2463,32'd-1217,32'd-869,32'd651,32'd-858,32'd1190,32'd2116,32'd-5571,32'd3269,32'd630,32'd-2193,32'd2478,32'd-2496,32'd-394,32'd2158,32'd2827,32'd2770,32'd-574,32'd-1055,32'd-855,32'd1859,32'd1206,32'd2097,32'd3300,32'd-4008,32'd2851,32'd-933,32'd-5527,32'd-1474,32'd-2902,32'd-2890,32'd2023,32'd-5390,32'd354,32'd-1269,32'd-95,32'd3088,32'd2553,32'd-2065,32'd2766,32'd1306,32'd7954,32'd2558,32'd4074,32'd4160,32'd975,32'd1101,32'd117,32'd4077,32'd6713,32'd3188,32'd65,32'd-1657,32'd1171,32'd-877,32'd-4907,32'd1933,32'd-4848,32'd-6308,32'd1865,32'd-1779,32'd-178,32'd-1400,32'd-2462,32'd1296,32'd-2629,32'd3371,32'd11474,32'd386,32'd4660,32'd4462,32'd-603,32'd3364,32'd-707,32'd3457,32'd-1071,32'd-160,32'd-354,32'd1766,32'd773,32'd4265,32'd1673,32'd5805,32'd240,32'd764,32'd-1097,32'd4460,32'd-6723,32'd2088,32'd1145,32'd-1910,32'd-1051,32'd-1185,32'd-10722,32'd-2203,32'd4831,32'd-4016,32'd5625,32'd-561,32'd3974,32'd-671,32'd-2805,32'd-3857,32'd-5229,32'd-3015,32'd2453,32'd1053,32'd-252,32'd2592,32'd-4938,32'd-613,32'd3305,32'd-7753,32'd-2988,32'd2910,32'd-1662,32'd-1021,32'd372,32'd-1567,32'd-4050,32'd3798,32'd-2800,32'd6665,32'd-3964,32'd-14,32'd578,32'd3842,32'd-5097,32'd6699,32'd3107,32'd2792,32'd2230,32'd879,32'd-4150,32'd2446,32'd1076,32'd2517,32'd-980,32'd-1518,32'd2044,32'd3156,32'd-1477,32'd-274,32'd-4052,32'd-1337,32'd-1403,32'd2675,32'd-1491,32'd-3955,32'd275,32'd4414,32'd-2956,32'd-7089,32'd-131,32'd-1633,32'd-8305,32'd-3471,32'd-1629,32'd351,32'd387,32'd-1198,32'd-1483,32'd970,32'd848,32'd-92,32'd-1187,32'd-1219,32'd3654,32'd597,32'd-2084,32'd-4257,32'd-3044,32'd-6376,32'd-2127,32'd3286,32'd-7373,32'd5009,32'd-197,32'd-3330,32'd-226,32'd-3525,32'd-259,32'd-1750,32'd-7358,32'd-4707,32'd1058,32'd-2766,32'd-4902,32'd-2011,32'd99,32'd368,32'd-34,32'd-4985,32'd-4833,32'd-4494,32'd-2758,32'd-9521,32'd-5517,32'd-4345,32'd-1505,32'd187,32'd-3247,32'd-953,32'd-5800,32'd2122,32'd-2410,32'd-1782,32'd-3183,32'd-548,32'd-2468,32'd-3293,32'd-1308,32'd-3984,32'd4553,32'd200,32'd-2296,32'd1951,32'd140,32'd6528,32'd466,32'd-3183,32'd-3403,32'd-4372,32'd-98,32'd8520,32'd3366,32'd-582,32'd1776,32'd560,32'd-528,32'd-2253,32'd1224,32'd1347,32'd-3557,32'd-2746,32'd-130,32'd-4433,32'd2196,32'd-5068,32'd3427,32'd-1656,32'd-1940,32'd-8559,32'd2958,32'd-1949,32'd822,32'd2893,32'd-2656,32'd-5815,32'd-2773,32'd2187,32'd44,32'd-6333,32'd-5024,32'd-3928,32'd-4736,32'd-3652,32'd-825,32'd-1301,32'd2880,32'd-1691,32'd-1078,32'd-3842,32'd-3337,32'd-3232,32'd-2675,32'd-8876,32'd-6508,32'd-7412,32'd617,32'd-6289,32'd-1217,32'd-3854,32'd7451,32'd68,32'd-4721,32'd6293,32'd-285,32'd-4387,32'd3803,32'd1431,32'd364,32'd-1947,32'd-2993,32'd-4641,32'd355,32'd-2521,32'd-1937,32'd791,32'd-865,32'd1857,32'd-2381,32'd-5415,32'd-4265,32'd-1734,32'd397,32'd-2690,32'd1907,32'd-6826,32'd3750,32'd3503,32'd1020,32'd-7924,32'd-1788,32'd6083,32'd-5317,32'd-7343,32'd-2995,32'd-5756,32'd4621,32'd-2792,32'd-5795,32'd-4589,32'd4550,32'd7016,32'd1373,32'd4174,32'd-5180,32'd-1992,32'd643,32'd-287,32'd-2052,32'd508,32'd-323,32'd2071,32'd-2081,32'd441,32'd-1688,32'd789,32'd662,32'd-4541,32'd-1185,32'd-4638};
    Wh[37]='{32'd-1599,32'd117,32'd-391,32'd-3774,32'd1353,32'd-654,32'd-1260,32'd1148,32'd3220,32'd897,32'd722,32'd263,32'd467,32'd-2312,32'd-2209,32'd-1433,32'd-7011,32'd-843,32'd1945,32'd2448,32'd1173,32'd-297,32'd-6660,32'd466,32'd-341,32'd2619,32'd946,32'd2442,32'd1334,32'd-2761,32'd874,32'd493,32'd-4628,32'd-4638,32'd776,32'd-2729,32'd-797,32'd-3828,32'd-147,32'd-2944,32'd-4536,32'd-2495,32'd6284,32'd1791,32'd364,32'd46,32'd-6875,32'd-1890,32'd-853,32'd1251,32'd2556,32'd-3476,32'd3056,32'd2832,32'd4941,32'd-548,32'd-2266,32'd369,32'd-5175,32'd-2663,32'd779,32'd888,32'd-5825,32'd-216,32'd-276,32'd1812,32'd-1628,32'd-5620,32'd912,32'd-649,32'd3466,32'd-999,32'd-1632,32'd223,32'd-2756,32'd3828,32'd-3098,32'd-57,32'd2519,32'd-426,32'd-3002,32'd-5410,32'd-358,32'd-5668,32'd1326,32'd-3012,32'd1745,32'd2261,32'd-523,32'd4147,32'd-2451,32'd-7065,32'd-208,32'd-608,32'd4855,32'd3676,32'd-1856,32'd33,32'd-1149,32'd-2103,32'd591,32'd780,32'd2631,32'd256,32'd-98,32'd-2519,32'd3049,32'd-1939,32'd4548,32'd-2388,32'd-2805,32'd202,32'd-1239,32'd-3393,32'd3303,32'd-3803,32'd-785,32'd2115,32'd-2910,32'd550,32'd3264,32'd2110,32'd-1883,32'd-628,32'd2705,32'd-932,32'd-4030,32'd-2241,32'd-1541,32'd10488,32'd-2617,32'd-3059,32'd1263,32'd-2459,32'd3476,32'd3095,32'd1200,32'd1605,32'd-3845,32'd-1899,32'd-441,32'd-2919,32'd2475,32'd-188,32'd4086,32'd-1584,32'd549,32'd1777,32'd-139,32'd2027,32'd3066,32'd4028,32'd255,32'd3283,32'd-8022,32'd-1446,32'd1254,32'd-2763,32'd3100,32'd-1248,32'd-4548,32'd-4560,32'd2293,32'd-4189,32'd3696,32'd3974,32'd1242,32'd1297,32'd-2536,32'd375,32'd-2978,32'd-3273,32'd3911,32'd856,32'd3852,32'd3144,32'd1597,32'd-3059,32'd1311,32'd-2153,32'd1325,32'd-4353,32'd-96,32'd-2325,32'd3630,32'd-2932,32'd-2036,32'd-4851,32'd-1008,32'd2421,32'd-3781,32'd3569,32'd-2775,32'd1440,32'd2374,32'd2445,32'd596,32'd-1101,32'd2812,32'd4201,32'd429,32'd2135,32'd-993,32'd-733,32'd564,32'd74,32'd655,32'd-2163,32'd539,32'd77,32'd-2788,32'd-3476,32'd-2326,32'd837,32'd3933,32'd-5727,32'd1752,32'd1516,32'd-2548,32'd662,32'd-1467,32'd3005,32'd-2379,32'd2198,32'd-80,32'd-3774,32'd-4326,32'd-1204,32'd-208,32'd242,32'd-611,32'd5253,32'd-3505,32'd1362,32'd-3940,32'd1067,32'd-7299,32'd814,32'd-1402,32'd-190,32'd718,32'd5136,32'd-4606,32'd3222,32'd1185,32'd-3059,32'd-3852,32'd-624,32'd-346,32'd-3293,32'd-123,32'd-3190,32'd-572,32'd-3098,32'd3369,32'd-1784,32'd-3359,32'd468,32'd-3618,32'd1151,32'd-6406,32'd-637,32'd1314,32'd-2316,32'd-2144,32'd-1757,32'd-3034,32'd4724,32'd477,32'd-41,32'd-3576,32'd-114,32'd-1433,32'd-283,32'd-84,32'd-2910,32'd-442,32'd-2038,32'd-2265,32'd-3540,32'd-460,32'd1511,32'd-2685,32'd2376,32'd-694,32'd5019,32'd-1959,32'd-464,32'd2379,32'd-1820,32'd-3330,32'd-1301,32'd1501,32'd1196,32'd3024,32'd521,32'd2263,32'd4431,32'd-3027,32'd-2348,32'd-739,32'd-2219,32'd-6049,32'd-3669,32'd1695,32'd-6308,32'd847,32'd1677,32'd1262,32'd122,32'd936,32'd-2213,32'd2521,32'd-5170,32'd-2427,32'd98,32'd505,32'd1411,32'd739,32'd-1943,32'd-3903,32'd-3354,32'd-4121,32'd-2169,32'd1657,32'd1228,32'd-1555,32'd-3969,32'd-5488,32'd-1166,32'd-3493,32'd-2919,32'd1599,32'd-2192,32'd1552,32'd-4282,32'd-2773,32'd2312,32'd5439,32'd868,32'd-2983,32'd2265,32'd3281,32'd7465,32'd-1121,32'd-5839,32'd2614,32'd-3671,32'd-4729,32'd370,32'd-709,32'd1257,32'd14,32'd859,32'd416,32'd-975,32'd-5332,32'd-6025,32'd-2243,32'd-247,32'd-1423,32'd1092,32'd-3027,32'd-3740,32'd3332,32'd-817,32'd-4458,32'd4919,32'd-803,32'd-9169,32'd9853,32'd-5576,32'd-4548,32'd-2932,32'd-6748,32'd1846,32'd-853,32'd3366,32'd5498,32'd-2075,32'd301,32'd1047,32'd-1242,32'd-2443,32'd-6455,32'd-1586,32'd345,32'd-1325,32'd1796,32'd-1021,32'd2529,32'd-3168,32'd2646,32'd413,32'd4338,32'd-4836,32'd35,32'd5014,32'd-3564,32'd-1566};
    Wh[38]='{32'd1875,32'd-481,32'd2773,32'd1027,32'd-3027,32'd486,32'd-249,32'd-3732,32'd-2369,32'd419,32'd-3813,32'd1235,32'd1894,32'd1466,32'd-4584,32'd-1103,32'd-560,32'd4489,32'd-6738,32'd2500,32'd1034,32'd634,32'd2291,32'd181,32'd33,32'd-2773,32'd-125,32'd-3010,32'd3012,32'd1606,32'd1756,32'd3183,32'd-1246,32'd1113,32'd173,32'd-2137,32'd245,32'd-2495,32'd614,32'd2218,32'd2539,32'd450,32'd5625,32'd2626,32'd3215,32'd2211,32'd-4633,32'd603,32'd-2683,32'd1035,32'd-5761,32'd2182,32'd3183,32'd1054,32'd-2829,32'd-159,32'd3273,32'd-190,32'd-3925,32'd2362,32'd-2062,32'd1574,32'd-1057,32'd-2316,32'd12,32'd390,32'd4057,32'd-5375,32'd-833,32'd-3247,32'd-1080,32'd-2785,32'd603,32'd1490,32'd1627,32'd2966,32'd-1978,32'd-1510,32'd-875,32'd-6386,32'd2127,32'd-8896,32'd2110,32'd12,32'd-1682,32'd-2325,32'd1295,32'd-808,32'd-4187,32'd-2238,32'd2775,32'd-812,32'd1978,32'd-5336,32'd5483,32'd938,32'd-5800,32'd936,32'd-3972,32'd-336,32'd-2307,32'd145,32'd713,32'd5615,32'd-5454,32'd4138,32'd-453,32'd2670,32'd1079,32'd1300,32'd-781,32'd-1500,32'd2753,32'd-5161,32'd3144,32'd5136,32'd4631,32'd-531,32'd-4450,32'd4523,32'd3171,32'd2160,32'd2910,32'd2302,32'd-533,32'd642,32'd593,32'd-3791,32'd812,32'd3361,32'd-3786,32'd-1862,32'd-2600,32'd1342,32'd-2604,32'd-898,32'd6684,32'd127,32'd-3454,32'd-1699,32'd5395,32'd-1495,32'd12167,32'd-1092,32'd-1192,32'd335,32'd-2048,32'd-1411,32'd4460,32'd878,32'd-3459,32'd5820,32'd-1510,32'd3107,32'd3061,32'd1867,32'd2059,32'd-2326,32'd3605,32'd1535,32'd-4870,32'd-8007,32'd1384,32'd-1287,32'd-1566,32'd2658,32'd-2895,32'd2895,32'd-1100,32'd3166,32'd-2413,32'd4904,32'd-5219,32'd-690,32'd-964,32'd-1141,32'd-1005,32'd-1798,32'd6689,32'd717,32'd-4350,32'd-6250,32'd560,32'd-1024,32'd408,32'd-1496,32'd8100,32'd-3874,32'd1822,32'd-9624,32'd773,32'd2056,32'd790,32'd2734,32'd-897,32'd-3078,32'd-1429,32'd-2531,32'd-90,32'd61,32'd-2287,32'd-1524,32'd-2819,32'd-2539,32'd-2612,32'd167,32'd756,32'd458,32'd-3715,32'd3581,32'd-785,32'd404,32'd-2121,32'd-166,32'd1204,32'd1634,32'd2104,32'd307,32'd2220,32'd-5048,32'd-2019,32'd-5102,32'd441,32'd-5122,32'd-1864,32'd-3361,32'd-4645,32'd587,32'd4252,32'd-6186,32'd416,32'd-1158,32'd-4223,32'd-2155,32'd-2856,32'd-6508,32'd-522,32'd-1540,32'd-5014,32'd1512,32'd-2075,32'd1611,32'd-2119,32'd-9052,32'd-665,32'd-1877,32'd7192,32'd-6787,32'd-404,32'd1995,32'd-144,32'd1607,32'd2050,32'd-3283,32'd-1361,32'd-5239,32'd375,32'd729,32'd667,32'd-115,32'd-3818,32'd1402,32'd4645,32'd-3830,32'd-709,32'd-1473,32'd-61,32'd1010,32'd-3386,32'd-2675,32'd773,32'd5249,32'd-1955,32'd741,32'd-1702,32'd-802,32'd3110,32'd-2683,32'd1790,32'd-353,32'd-1080,32'd-3383,32'd1042,32'd937,32'd-2203,32'd-2880,32'd2149,32'd-716,32'd8,32'd2890,32'd-1702,32'd-5136,32'd-2497,32'd3054,32'd3320,32'd550,32'd-2164,32'd-3017,32'd1741,32'd1308,32'd-1234,32'd226,32'd5517,32'd-626,32'd-839,32'd-5986,32'd-2161,32'd2363,32'd-272,32'd-1610,32'd-631,32'd-2302,32'd2705,32'd695,32'd-5146,32'd-468,32'd3269,32'd-2429,32'd3256,32'd-3410,32'd-1198,32'd369,32'd1384,32'd-5483,32'd2313,32'd896,32'd382,32'd-2690,32'd-1101,32'd1505,32'd196,32'd222,32'd3457,32'd-6469,32'd-5019,32'd371,32'd-1881,32'd-1365,32'd1612,32'd-1875,32'd4326,32'd-1928,32'd-1100,32'd547,32'd-406,32'd-2148,32'd-2486,32'd4196,32'd5146,32'd3676,32'd-315,32'd-6220,32'd3645,32'd-2844,32'd-2288,32'd-1384,32'd6049,32'd3891,32'd-2622,32'd-1697,32'd-1300,32'd4531,32'd1556,32'd-4758,32'd712,32'd-1545,32'd1684,32'd-4516,32'd2919,32'd-7602,32'd-2073,32'd2666,32'd-2622,32'd-11220,32'd-122,32'd377,32'd-1293,32'd1323,32'd-3833,32'd2509,32'd1280,32'd2739,32'd3449,32'd966,32'd-2797,32'd5751,32'd2384,32'd750,32'd-2822,32'd4296,32'd-226,32'd5053,32'd4631,32'd1877,32'd-1171,32'd4370,32'd-2362,32'd5083,32'd4121,32'd1915};
    Wh[39]='{32'd2780,32'd217,32'd-290,32'd-1810,32'd-843,32'd-810,32'd3095,32'd1645,32'd-4274,32'd2252,32'd3767,32'd91,32'd-5761,32'd928,32'd-1567,32'd-1006,32'd4770,32'd-1829,32'd1606,32'd755,32'd4221,32'd-878,32'd1145,32'd-3178,32'd-1385,32'd-1076,32'd-285,32'd1801,32'd-2819,32'd2413,32'd1876,32'd4213,32'd5458,32'd5991,32'd995,32'd-4213,32'd-1518,32'd1060,32'd72,32'd2778,32'd2117,32'd-931,32'd-1328,32'd-373,32'd4599,32'd1933,32'd-2095,32'd-2551,32'd331,32'd-531,32'd1971,32'd502,32'd4855,32'd-8471,32'd1793,32'd3398,32'd3454,32'd2261,32'd3486,32'd-1166,32'd819,32'd2015,32'd-1450,32'd-1904,32'd7910,32'd2817,32'd1228,32'd7290,32'd-3659,32'd5161,32'd-639,32'd2390,32'd6523,32'd448,32'd5341,32'd-386,32'd-1898,32'd39,32'd-3073,32'd-3557,32'd-70,32'd-76,32'd4228,32'd-6289,32'd6064,32'd-4411,32'd2592,32'd3637,32'd-3640,32'd2198,32'd2,32'd5029,32'd2961,32'd5878,32'd1196,32'd283,32'd1870,32'd-834,32'd-2454,32'd-443,32'd-6489,32'd2346,32'd2214,32'd-4440,32'd-5390,32'd-545,32'd4079,32'd1613,32'd-1672,32'd5771,32'd2836,32'd-1429,32'd-8735,32'd1932,32'd3635,32'd-2474,32'd1247,32'd-8554,32'd792,32'd4648,32'd1652,32'd-7465,32'd-3020,32'd-807,32'd-110,32'd-659,32'd-4028,32'd-2423,32'd7524,32'd-349,32'd-9711,32'd-4777,32'd1054,32'd-3874,32'd-3173,32'd-3576,32'd-2408,32'd2148,32'd4709,32'd-2829,32'd-5361,32'd1887,32'd975,32'd-1352,32'd1051,32'd-2844,32'd-3933,32'd-1665,32'd-277,32'd-1901,32'd9116,32'd-2012,32'd5297,32'd114,32'd3425,32'd-344,32'd1457,32'd-4353,32'd-2403,32'd-1281,32'd-5688,32'd310,32'd-2061,32'd4284,32'd5136,32'd2482,32'd113,32'd-709,32'd4304,32'd367,32'd-4692,32'd-1384,32'd8188,32'd-4411,32'd-3715,32'd2048,32'd-2973,32'd105,32'd-6982,32'd3093,32'd-3786,32'd15175,32'd-903,32'd-5483,32'd-1065,32'd-6220,32'd-1075,32'd-60,32'd-5786,32'd5180,32'd3356,32'd2873,32'd533,32'd5747,32'd3571,32'd-11220,32'd-3288,32'd7182,32'd2399,32'd794,32'd-1771,32'd3210,32'd482,32'd-1961,32'd880,32'd194,32'd-1684,32'd2459,32'd2541,32'd6152,32'd8671,32'd2773,32'd481,32'd-453,32'd8686,32'd18,32'd-2719,32'd966,32'd-709,32'd4025,32'd936,32'd2115,32'd4707,32'd5141,32'd6059,32'd-3156,32'd3813,32'd-1783,32'd-1772,32'd320,32'd2397,32'd-4150,32'd-1461,32'd-88,32'd-509,32'd-2183,32'd-303,32'd553,32'd4526,32'd2293,32'd2092,32'd-2553,32'd5068,32'd4223,32'd56,32'd172,32'd851,32'd4343,32'd3588,32'd-1679,32'd2381,32'd-300,32'd1252,32'd-1016,32'd-2211,32'd-1046,32'd-3320,32'd113,32'd-897,32'd5605,32'd2474,32'd2590,32'd258,32'd5546,32'd2878,32'd304,32'd2132,32'd-2019,32'd-1472,32'd1529,32'd1284,32'd-2553,32'd-3708,32'd-213,32'd3776,32'd-327,32'd-4609,32'd-44,32'd3215,32'd-1157,32'd-4128,32'd-4,32'd1865,32'd-601,32'd3039,32'd1949,32'd43,32'd-3400,32'd-1834,32'd983,32'd-3632,32'd7309,32'd-650,32'd975,32'd-3486,32'd11083,32'd530,32'd3723,32'd2117,32'd-5991,32'd-158,32'd-3093,32'd-8056,32'd3613,32'd-1859,32'd6577,32'd-5498,32'd1424,32'd2446,32'd-820,32'd3950,32'd3908,32'd-1892,32'd3188,32'd-3862,32'd2854,32'd-4025,32'd-4184,32'd4301,32'd5014,32'd5351,32'd2248,32'd-167,32'd562,32'd709,32'd-1671,32'd122,32'd-741,32'd234,32'd242,32'd3564,32'd-4467,32'd-3784,32'd481,32'd615,32'd2261,32'd-7221,32'd5581,32'd-1398,32'd-732,32'd85,32'd3876,32'd2349,32'd-3198,32'd-4934,32'd1793,32'd-748,32'd4440,32'd7304,32'd-3486,32'd-1183,32'd8779,32'd-4306,32'd3164,32'd-3222,32'd-3364,32'd3630,32'd-1668,32'd-4135,32'd5410,32'd1497,32'd-6855,32'd1794,32'd572,32'd-6083,32'd-1809,32'd-495,32'd-7929,32'd512,32'd938,32'd-581,32'd-6210,32'd1492,32'd891,32'd-1159,32'd472,32'd-5415,32'd-2268,32'd1467,32'd407,32'd-4121,32'd-6376,32'd985,32'd-4301,32'd-3342,32'd-3190,32'd1143,32'd-3691,32'd-2895,32'd-2436,32'd-1909,32'd-1577,32'd9062,32'd3249,32'd2756,32'd-3198,32'd-24,32'd2330,32'd3647,32'd913};
    Wh[40]='{32'd914,32'd4023,32'd2384,32'd-2541,32'd-3142,32'd2746,32'd1883,32'd6098,32'd1859,32'd-1303,32'd3374,32'd2017,32'd799,32'd138,32'd6386,32'd-513,32'd-1429,32'd-150,32'd402,32'd-2561,32'd25,32'd965,32'd2402,32'd-32,32'd-343,32'd-3654,32'd701,32'd480,32'd-2305,32'd-982,32'd-1611,32'd-3085,32'd4880,32'd-421,32'd-2216,32'd6835,32'd206,32'd-1119,32'd-4672,32'd2297,32'd532,32'd3896,32'd-2277,32'd-1596,32'd4680,32'd1420,32'd1767,32'd3730,32'd4052,32'd747,32'd-2761,32'd2486,32'd1003,32'd-3640,32'd-3818,32'd5664,32'd180,32'd3071,32'd-1741,32'd1030,32'd1099,32'd2966,32'd3881,32'd-1641,32'd-1945,32'd-3022,32'd-383,32'd5854,32'd-2148,32'd755,32'd-7290,32'd-2414,32'd1909,32'd5722,32'd4213,32'd2851,32'd-1577,32'd1839,32'd-4167,32'd2171,32'd2707,32'd-126,32'd3093,32'd4638,32'd-1273,32'd476,32'd3391,32'd-1362,32'd5429,32'd-1884,32'd2254,32'd-1267,32'd-4147,32'd-243,32'd1470,32'd-1761,32'd-1411,32'd-1351,32'd707,32'd2126,32'd-3417,32'd482,32'd-3107,32'd1539,32'd-2856,32'd-1021,32'd-2114,32'd748,32'd-4780,32'd455,32'd-3613,32'd2277,32'd4829,32'd4287,32'd3483,32'd127,32'd-3715,32'd-1300,32'd-3588,32'd-5126,32'd-601,32'd-1242,32'd2705,32'd3818,32'd-1248,32'd2856,32'd1076,32'd-1636,32'd-568,32'd2746,32'd209,32'd2303,32'd-2412,32'd1346,32'd820,32'd-1516,32'd4025,32'd-4282,32'd2330,32'd-1389,32'd-4218,32'd-2575,32'd2595,32'd-1158,32'd3203,32'd-2661,32'd-1370,32'd-935,32'd-2980,32'd-1805,32'd-3454,32'd764,32'd4016,32'd-2915,32'd-687,32'd8496,32'd-4182,32'd1011,32'd-238,32'd12773,32'd1759,32'd2145,32'd1233,32'd-3837,32'd-2968,32'd178,32'd1163,32'd4699,32'd-1643,32'd18,32'd-134,32'd1114,32'd3090,32'd1933,32'd-919,32'd-1314,32'd-649,32'd-3073,32'd1778,32'd737,32'd-4272,32'd-994,32'd-1716,32'd6235,32'd-3830,32'd983,32'd449,32'd6,32'd-4592,32'd-886,32'd972,32'd1949,32'd1193,32'd-397,32'd-3583,32'd-838,32'd-1817,32'd-1811,32'd-1939,32'd5131,32'd1309,32'd-5576,32'd1041,32'd-1081,32'd-1959,32'd1562,32'd-3898,32'd-3288,32'd5146,32'd-1547,32'd-1331,32'd3959,32'd150,32'd-4526,32'd-852,32'd602,32'd-981,32'd4042,32'd5380,32'd2514,32'd694,32'd-1851,32'd-360,32'd1194,32'd-520,32'd-4404,32'd2053,32'd-169,32'd4594,32'd-597,32'd-605,32'd-2225,32'd-3588,32'd591,32'd-4028,32'd-2309,32'd-1210,32'd-2609,32'd-585,32'd-2519,32'd-1290,32'd-4016,32'd-783,32'd-1437,32'd-1129,32'd240,32'd7080,32'd-2092,32'd389,32'd-48,32'd2000,32'd-73,32'd-598,32'd-1038,32'd-2839,32'd-1939,32'd3400,32'd-3195,32'd2541,32'd-1014,32'd3164,32'd207,32'd-3027,32'd508,32'd-1423,32'd-2739,32'd1737,32'd1333,32'd766,32'd-313,32'd-1959,32'd-4499,32'd1181,32'd-539,32'd3676,32'd-1644,32'd-1778,32'd1301,32'd1117,32'd2313,32'd7211,32'd623,32'd-1940,32'd1813,32'd1124,32'd827,32'd2297,32'd-89,32'd2025,32'd-2646,32'd715,32'd-259,32'd871,32'd-2243,32'd-2731,32'd4838,32'd-831,32'd1285,32'd-845,32'd-2568,32'd759,32'd-4392,32'd10253,32'd-88,32'd-5117,32'd4614,32'd591,32'd2524,32'd7939,32'd-2158,32'd110,32'd-2318,32'd5849,32'd-3876,32'd-2585,32'd2281,32'd-3911,32'd2312,32'd1218,32'd1853,32'd-954,32'd4050,32'd-2663,32'd457,32'd-615,32'd-6210,32'd-1268,32'd3156,32'd-5102,32'd-626,32'd-4379,32'd-2230,32'd21,32'd-600,32'd853,32'd13,32'd1688,32'd2656,32'd-466,32'd1047,32'd3903,32'd2548,32'd-3994,32'd4846,32'd7177,32'd-181,32'd-9316,32'd2407,32'd0,32'd-2856,32'd-540,32'd-1933,32'd312,32'd826,32'd1055,32'd4526,32'd7319,32'd-3554,32'd603,32'd-2397,32'd-3745,32'd-2619,32'd4479,32'd-6718,32'd1251,32'd1827,32'd8276,32'd-7504,32'd6049,32'd1268,32'd-360,32'd4018,32'd-1506,32'd5317,32'd1542,32'd2242,32'd-4216,32'd2022,32'd-2648,32'd238,32'd8037,32'd1209,32'd5854,32'd4162,32'd2305,32'd2717,32'd2731,32'd600,32'd2027,32'd4775,32'd-76,32'd2563,32'd-3605,32'd-379,32'd11972,32'd-466,32'd1926,32'd1861,32'd-31,32'd-985};
    Wh[41]='{32'd2856,32'd-838,32'd-584,32'd591,32'd2692,32'd1584,32'd552,32'd-7509,32'd2844,32'd2137,32'd-2320,32'd2235,32'd1314,32'd1677,32'd1763,32'd588,32'd-7045,32'd1612,32'd-2443,32'd-1882,32'd1872,32'd2653,32'd-465,32'd-2471,32'd-1315,32'd-3789,32'd-2084,32'd-432,32'd-4265,32'd-482,32'd2288,32'd-4155,32'd-7578,32'd1223,32'd2746,32'd-2436,32'd-69,32'd-1199,32'd1958,32'd-1950,32'd-2373,32'd-2792,32'd2114,32'd-8012,32'd-561,32'd3361,32'd-1690,32'd1942,32'd-1892,32'd17,32'd119,32'd7011,32'd-454,32'd-870,32'd4365,32'd-5195,32'd-1383,32'd-1280,32'd-2785,32'd6562,32'd-3798,32'd-1840,32'd823,32'd1483,32'd-400,32'd-831,32'd1933,32'd-172,32'd3735,32'd157,32'd2810,32'd-2381,32'd-852,32'd-3867,32'd-1234,32'd3403,32'd476,32'd-4843,32'd2775,32'd2000,32'd1535,32'd2687,32'd-2076,32'd-4379,32'd-1868,32'd-3911,32'd-3002,32'd-4345,32'd1311,32'd8198,32'd1422,32'd2512,32'd-3181,32'd637,32'd1514,32'd1478,32'd4624,32'd70,32'd-2902,32'd-2155,32'd-6533,32'd2462,32'd936,32'd-9301,32'd11591,32'd-378,32'd-2058,32'd4624,32'd-2724,32'd-2993,32'd-3515,32'd4331,32'd9570,32'd-3830,32'd-134,32'd960,32'd-2161,32'd220,32'd1737,32'd-4797,32'd-1495,32'd-4848,32'd-11650,32'd-3259,32'd975,32'd-3278,32'd3479,32'd2683,32'd434,32'd-1437,32'd1214,32'd-5234,32'd-55,32'd-6684,32'd-3706,32'd-5253,32'd1904,32'd-2600,32'd-1539,32'd1148,32'd-623,32'd126,32'd2366,32'd-723,32'd2363,32'd-4445,32'd1909,32'd-11201,32'd-4953,32'd2973,32'd4604,32'd-650,32'd1517,32'd-996,32'd104,32'd-1931,32'd-3776,32'd-3662,32'd858,32'd-12988,32'd9311,32'd273,32'd-1224,32'd1303,32'd-1506,32'd-397,32'd-3156,32'd-777,32'd1926,32'd4584,32'd-2056,32'd-2176,32'd-4831,32'd-6391,32'd-6547,32'd-191,32'd-2565,32'd9033,32'd2492,32'd-3476,32'd8007,32'd5615,32'd-381,32'd-2612,32'd1232,32'd-2246,32'd3813,32'd3073,32'd3171,32'd2727,32'd1856,32'd942,32'd2998,32'd-2203,32'd-1961,32'd-545,32'd-147,32'd3041,32'd413,32'd-1193,32'd1777,32'd-2727,32'd1745,32'd7290,32'd741,32'd2431,32'd-1865,32'd2375,32'd-3295,32'd4208,32'd3146,32'd-6323,32'd5122,32'd7509,32'd4819,32'd2739,32'd1474,32'd573,32'd-3305,32'd3579,32'd-174,32'd228,32'd2429,32'd2130,32'd1735,32'd2727,32'd-256,32'd-1315,32'd2600,32'd-1093,32'd1205,32'd874,32'd2130,32'd6835,32'd-102,32'd-3352,32'd-1216,32'd4692,32'd5517,32'd5463,32'd-600,32'd-2824,32'd4990,32'd2673,32'd-1689,32'd678,32'd-7719,32'd-5058,32'd3215,32'd1966,32'd4172,32'd1573,32'd1551,32'd9,32'd-2397,32'd-884,32'd-4079,32'd4692,32'd-3518,32'd-3107,32'd-2556,32'd2445,32'd-7436,32'd1956,32'd-1375,32'd3041,32'd1704,32'd1056,32'd615,32'd1691,32'd-6093,32'd894,32'd-790,32'd3886,32'd-5776,32'd382,32'd-1502,32'd3305,32'd-3054,32'd-716,32'd-762,32'd-5571,32'd2976,32'd3029,32'd2634,32'd6250,32'd-4797,32'd5161,32'd877,32'd-17,32'd-30,32'd8901,32'd4372,32'd-781,32'd2121,32'd3452,32'd150,32'd638,32'd-8940,32'd709,32'd80,32'd-1564,32'd-1593,32'd5839,32'd-2050,32'd5551,32'd-2373,32'd6337,32'd-1956,32'd-4204,32'd-3291,32'd-3217,32'd2403,32'd1441,32'd-1759,32'd-1861,32'd-8959,32'd4606,32'd262,32'd2988,32'd1787,32'd-3642,32'd-4106,32'd1643,32'd1386,32'd133,32'd-2290,32'd9267,32'd4719,32'd-2313,32'd4633,32'd-2998,32'd-1241,32'd1627,32'd-2995,32'd3449,32'd3315,32'd612,32'd-2863,32'd2678,32'd-3312,32'd2800,32'd1740,32'd-1298,32'd370,32'd197,32'd3686,32'd5693,32'd-9931,32'd-3747,32'd2481,32'd8989,32'd-1667,32'd-218,32'd3894,32'd-2331,32'd-1802,32'd2182,32'd4538,32'd-2159,32'd2536,32'd-2078,32'd-396,32'd1789,32'd2253,32'd-4902,32'd3037,32'd1029,32'd1821,32'd-232,32'd721,32'd99,32'd119,32'd9296,32'd3679,32'd290,32'd-2043,32'd-2442,32'd-830,32'd-3662,32'd-3583,32'd-2355,32'd-3471,32'd-2106,32'd3190,32'd1722,32'd-6333,32'd994,32'd-2639,32'd-867,32'd2460,32'd-788,32'd-4882,32'd-4069,32'd-2420,32'd-1651,32'd-3364,32'd930,32'd-2266,32'd1895};
    Wh[42]='{32'd9575,32'd1096,32'd1463,32'd-2120,32'd-3376,32'd3620,32'd6357,32'd-5239,32'd4128,32'd622,32'd-215,32'd-3688,32'd1580,32'd875,32'd157,32'd5317,32'd-1440,32'd-970,32'd-4316,32'd-2880,32'd2274,32'd2543,32'd635,32'd419,32'd1921,32'd5800,32'd-173,32'd1295,32'd4162,32'd-2313,32'd1810,32'd1844,32'd-668,32'd-1450,32'd312,32'd-1618,32'd2242,32'd3293,32'd1616,32'd-2445,32'd-1300,32'd190,32'd-6752,32'd516,32'd-2302,32'd1163,32'd2064,32'd-1233,32'd231,32'd-2476,32'd811,32'd-3215,32'd-4782,32'd1173,32'd-3869,32'd1815,32'd2951,32'd468,32'd1173,32'd1459,32'd-1763,32'd-319,32'd-4931,32'd309,32'd3613,32'd3808,32'd1425,32'd-899,32'd66,32'd-384,32'd-516,32'd1423,32'd-3747,32'd-2807,32'd3876,32'd-3554,32'd5776,32'd-2198,32'd-2475,32'd3010,32'd-2863,32'd2409,32'd48,32'd2152,32'd266,32'd440,32'd-433,32'd941,32'd-247,32'd5395,32'd-374,32'd-2395,32'd3793,32'd4467,32'd-2475,32'd-4125,32'd-2368,32'd-1934,32'd1170,32'd2229,32'd-3630,32'd1759,32'd-961,32'd6621,32'd-3288,32'd-496,32'd-3615,32'd4697,32'd415,32'd-4799,32'd-3190,32'd3212,32'd5854,32'd-2462,32'd-623,32'd1586,32'd-3122,32'd-3774,32'd-1744,32'd-721,32'd-1904,32'd1625,32'd7602,32'd2597,32'd-3715,32'd470,32'd7539,32'd2504,32'd1828,32'd-4719,32'd-1649,32'd-1148,32'd3977,32'd-1330,32'd-2639,32'd1774,32'd9897,32'd-1121,32'd4394,32'd555,32'd4106,32'd-882,32'd-15263,32'd634,32'd-4826,32'd333,32'd1914,32'd-3789,32'd-26,32'd2768,32'd-2429,32'd2084,32'd-6376,32'd5771,32'd8281,32'd-1341,32'd-221,32'd-1953,32'd1101,32'd5356,32'd6718,32'd-2829,32'd414,32'd-807,32'd-6215,32'd-10498,32'd-807,32'd1511,32'd1174,32'd1270,32'd-6645,32'd-599,32'd-4416,32'd-4020,32'd1654,32'd-1864,32'd-1849,32'd289,32'd727,32'd6445,32'd692,32'd-1896,32'd-1336,32'd1234,32'd-3640,32'd3803,32'd4160,32'd-710,32'd-2127,32'd8159,32'd5419,32'd2061,32'd3388,32'd-1331,32'd86,32'd-1466,32'd-4221,32'd-6230,32'd2536,32'd1805,32'd-1922,32'd-2237,32'd-9589,32'd851,32'd-529,32'd-2163,32'd4941,32'd-238,32'd389,32'd4750,32'd789,32'd3076,32'd-1292,32'd1613,32'd4709,32'd2059,32'd2648,32'd-1430,32'd5908,32'd-5063,32'd535,32'd870,32'd4377,32'd1589,32'd1474,32'd4597,32'd3066,32'd1485,32'd3703,32'd209,32'd-2717,32'd1756,32'd2543,32'd4150,32'd3366,32'd548,32'd4182,32'd-1217,32'd6191,32'd2509,32'd-5820,32'd1458,32'd5561,32'd-975,32'd4055,32'd-3491,32'd7138,32'd-4360,32'd1542,32'd720,32'd4064,32'd1845,32'd3098,32'd-2504,32'd-6313,32'd-4106,32'd4882,32'd-4494,32'd-549,32'd5947,32'd-969,32'd872,32'd2156,32'd-1888,32'd3952,32'd1026,32'd1704,32'd595,32'd3471,32'd-169,32'd503,32'd6118,32'd1511,32'd2327,32'd4025,32'd1181,32'd-874,32'd6445,32'd3532,32'd-1934,32'd1524,32'd-420,32'd2810,32'd1816,32'd671,32'd808,32'd-1040,32'd-1724,32'd-1045,32'd-1801,32'd-1362,32'd3564,32'd46,32'd2580,32'd-3576,32'd2006,32'd-3564,32'd-430,32'd1584,32'd5976,32'd4077,32'd2194,32'd-2149,32'd-3305,32'd-905,32'd1148,32'd1583,32'd6250,32'd3662,32'd3559,32'd1113,32'd-993,32'd-451,32'd2800,32'd-2017,32'd3674,32'd5996,32'd3828,32'd2800,32'd38,32'd-2161,32'd1370,32'd1376,32'd2341,32'd-4670,32'd59,32'd-3576,32'd-3767,32'd1132,32'd-3540,32'd3376,32'd6093,32'd3032,32'd3615,32'd3935,32'd2661,32'd3281,32'd-8774,32'd-1345,32'd6337,32'd880,32'd1809,32'd-7680,32'd5366,32'd-2844,32'd-2375,32'd880,32'd1956,32'd-774,32'd2073,32'd-4108,32'd1339,32'd-3618,32'd2795,32'd-7939,32'd172,32'd7773,32'd3183,32'd1021,32'd3862,32'd3442,32'd1306,32'd6108,32'd596,32'd1055,32'd381,32'd-440,32'd2673,32'd1345,32'd-3972,32'd2012,32'd3266,32'd1386,32'd4189,32'd-1165,32'd5991,32'd-303,32'd3461,32'd-2719,32'd2303,32'd-1928,32'd1170,32'd-894,32'd-123,32'd-756,32'd4560,32'd5063,32'd2514,32'd4436,32'd-4975,32'd2587,32'd3723,32'd6210,32'd-4155,32'd3430,32'd1690,32'd-6723,32'd5014,32'd4604,32'd6738};
    Wh[43]='{32'd-415,32'd1292,32'd-1525,32'd2315,32'd-2136,32'd1420,32'd4206,32'd2268,32'd2641,32'd1623,32'd6967,32'd-944,32'd1684,32'd-5053,32'd-117,32'd-3937,32'd-3503,32'd5019,32'd4721,32'd-447,32'd-218,32'd-349,32'd-1012,32'd-1846,32'd2460,32'd1021,32'd-364,32'd-1663,32'd3933,32'd-2773,32'd-2454,32'd-3881,32'd5405,32'd4443,32'd448,32'd7866,32'd1188,32'd489,32'd3696,32'd-462,32'd1040,32'd-4299,32'd-595,32'd1469,32'd-878,32'd5136,32'd-2624,32'd69,32'd1915,32'd-1776,32'd-5053,32'd-88,32'd5683,32'd-985,32'd2001,32'd3574,32'd2207,32'd-3164,32'd5727,32'd-630,32'd280,32'd8056,32'd1090,32'd-3146,32'd-3369,32'd712,32'd1245,32'd-1053,32'd-2934,32'd464,32'd1084,32'd149,32'd-2313,32'd-3742,32'd-1209,32'd1385,32'd-2093,32'd-2609,32'd483,32'd2687,32'd-3242,32'd-10673,32'd-1056,32'd8295,32'd-381,32'd-4523,32'd-789,32'd11933,32'd397,32'd-7094,32'd1909,32'd-3825,32'd138,32'd-5039,32'd588,32'd1712,32'd3195,32'd297,32'd3571,32'd-896,32'd7236,32'd6000,32'd717,32'd-12500,32'd5073,32'd-238,32'd-6489,32'd3708,32'd7983,32'd1369,32'd5917,32'd-6132,32'd-3444,32'd2281,32'd1124,32'd-1892,32'd454,32'd-3889,32'd-1601,32'd-2375,32'd282,32'd-2435,32'd-14335,32'd-8906,32'd-6943,32'd-3544,32'd1910,32'd-2041,32'd4379,32'd-4213,32'd-1045,32'd-2861,32'd3200,32'd-2316,32'd1328,32'd-1258,32'd-3735,32'd-4685,32'd1313,32'd3408,32'd-440,32'd2265,32'd1118,32'd1475,32'd1123,32'd985,32'd3994,32'd1998,32'd4782,32'd2873,32'd802,32'd-235,32'd-4321,32'd-1610,32'd2,32'd-6274,32'd2983,32'd1802,32'd5336,32'd-5527,32'd2489,32'd-2200,32'd-840,32'd-2301,32'd2418,32'd-4614,32'd440,32'd-2541,32'd-4113,32'd-7304,32'd-496,32'd-2875,32'd4689,32'd-3037,32'd-15,32'd3090,32'd474,32'd130,32'd-1687,32'd-1970,32'd249,32'd-1295,32'd2427,32'd-5883,32'd1547,32'd1209,32'd386,32'd343,32'd7133,32'd-3515,32'd-254,32'd1058,32'd-5722,32'd19,32'd8110,32'd-5898,32'd205,32'd-4943,32'd850,32'd2839,32'd-1168,32'd-249,32'd-2092,32'd-9277,32'd-4084,32'd-1228,32'd4270,32'd1815,32'd-4162,32'd-1950,32'd-4736,32'd1756,32'd-972,32'd-2922,32'd165,32'd1884,32'd1174,32'd-9194,32'd2910,32'd-1326,32'd-635,32'd5253,32'd2218,32'd-1674,32'd-2183,32'd177,32'd-5908,32'd-1256,32'd1546,32'd-3684,32'd-4565,32'd670,32'd-2425,32'd690,32'd-7812,32'd-1574,32'd3269,32'd681,32'd3713,32'd-2775,32'd-8305,32'd-3532,32'd-2290,32'd-46,32'd-5698,32'd-961,32'd2824,32'd-520,32'd-5532,32'd429,32'd-1350,32'd-1528,32'd-3947,32'd-5698,32'd-1005,32'd-5273,32'd-2612,32'd6264,32'd-737,32'd-2675,32'd-4257,32'd-5673,32'd1680,32'd-1314,32'd-991,32'd-2775,32'd-5458,32'd781,32'd-3117,32'd964,32'd-2573,32'd3115,32'd1083,32'd-3908,32'd-2135,32'd1236,32'd1446,32'd5317,32'd4523,32'd3032,32'd1132,32'd5415,32'd-7739,32'd-2690,32'd879,32'd-1575,32'd-2531,32'd761,32'd-2729,32'd1949,32'd-1168,32'd2249,32'd-3342,32'd-3012,32'd3088,32'd13,32'd-3806,32'd-3842,32'd-3786,32'd424,32'd-1357,32'd-703,32'd-3237,32'd-4465,32'd-6865,32'd-7978,32'd3266,32'd5019,32'd3591,32'd866,32'd1951,32'd-2432,32'd2846,32'd6870,32'd-1628,32'd-1815,32'd8979,32'd-1827,32'd-1402,32'd3986,32'd-7080,32'd921,32'd5668,32'd-642,32'd-1067,32'd-1478,32'd-2136,32'd-1467,32'd3161,32'd-5761,32'd-2167,32'd-3840,32'd-3732,32'd2027,32'd5400,32'd-1492,32'd5683,32'd1002,32'd5517,32'd-3242,32'd-4868,32'd-6704,32'd-1719,32'd-5595,32'd-413,32'd1658,32'd380,32'd-1279,32'd-2496,32'd471,32'd-3642,32'd-113,32'd-4108,32'd-7856,32'd-401,32'd1417,32'd-2054,32'd1175,32'd-6621,32'd-155,32'd-2612,32'd-977,32'd-1125,32'd-6796,32'd-4519,32'd3691,32'd-1591,32'd-4250,32'd1030,32'd1691,32'd629,32'd-3395,32'd-2597,32'd-9106,32'd-943,32'd-1722,32'd-703,32'd-3898,32'd-1434,32'd5117,32'd144,32'd1005,32'd381,32'd899,32'd-5927,32'd-864,32'd-6904,32'd-1105,32'd1286,32'd-2194,32'd679,32'd-2171,32'd-6166,32'd6938,32'd2238,32'd-3205,32'd2749,32'd-1506,32'd7431,32'd-3557};
    Wh[44]='{32'd-3271,32'd-6044,32'd-59,32'd3796,32'd-3996,32'd-2534,32'd-3747,32'd-914,32'd-1286,32'd-2939,32'd-1497,32'd121,32'd2028,32'd376,32'd-2739,32'd-693,32'd-2614,32'd-4396,32'd-1983,32'd4414,32'd4096,32'd-1012,32'd5903,32'd655,32'd-6166,32'd2646,32'd779,32'd-1905,32'd-1635,32'd1838,32'd4206,32'd1069,32'd-3176,32'd5317,32'd-632,32'd2011,32'd-2651,32'd5917,32'd-1904,32'd186,32'd170,32'd-931,32'd-4775,32'd872,32'd1079,32'd1564,32'd2915,32'd2376,32'd-3552,32'd-10869,32'd-334,32'd2260,32'd847,32'd-934,32'd-1791,32'd-946,32'd-14,32'd6918,32'd1020,32'd-2824,32'd2817,32'd1433,32'd3210,32'd234,32'd-2651,32'd3303,32'd-1315,32'd-1479,32'd2163,32'd584,32'd-3950,32'd2448,32'd2922,32'd2109,32'd3864,32'd6142,32'd-5029,32'd2961,32'd1630,32'd730,32'd-571,32'd3432,32'd836,32'd3581,32'd-726,32'd-567,32'd418,32'd461,32'd2517,32'd-3332,32'd-429,32'd-2244,32'd7260,32'd422,32'd891,32'd-3286,32'd-5102,32'd-5419,32'd459,32'd1362,32'd2915,32'd-5839,32'd661,32'd-4775,32'd-3159,32'd2451,32'd-829,32'd2802,32'd-713,32'd6577,32'd1491,32'd-8193,32'd-15625,32'd-885,32'd4211,32'd-12,32'd4274,32'd3981,32'd-2531,32'd7324,32'd1124,32'd-2988,32'd943,32'd-6030,32'd-1855,32'd-13828,32'd1539,32'd6689,32'd8637,32'd-6308,32'd12275,32'd-9819,32'd210,32'd-2260,32'd3564,32'd-4843,32'd-4421,32'd-4523,32'd2440,32'd2668,32'd319,32'd-2270,32'd-443,32'd-5722,32'd-4372,32'd-4296,32'd318,32'd-2465,32'd7700,32'd-5190,32'd1232,32'd2819,32'd10205,32'd-3186,32'd7333,32'd-28,32'd-729,32'd577,32'd745,32'd-13457,32'd3483,32'd3710,32'd-2702,32'd-1298,32'd175,32'd-7065,32'd2641,32'd2370,32'd-557,32'd-1322,32'd8208,32'd-2023,32'd5737,32'd-3461,32'd6630,32'd3261,32'd3364,32'd567,32'd-4616,32'd2009,32'd5688,32'd-1229,32'd2587,32'd-2094,32'd2283,32'd2988,32'd9057,32'd2729,32'd6103,32'd-7519,32'd-338,32'd-2279,32'd-1492,32'd3134,32'd-4621,32'd-1018,32'd-6977,32'd-5737,32'd3164,32'd-870,32'd-3361,32'd7700,32'd-18,32'd4182,32'd-1677,32'd197,32'd4436,32'd-1013,32'd2678,32'd-1666,32'd2763,32'd4826,32'd2529,32'd-249,32'd4211,32'd9057,32'd6704,32'd-381,32'd7304,32'd3596,32'd3742,32'd4599,32'd7500,32'd-6201,32'd3828,32'd3476,32'd745,32'd2514,32'd986,32'd4599,32'd-457,32'd888,32'd3415,32'd5102,32'd-674,32'd3332,32'd2242,32'd3288,32'd6113,32'd-3557,32'd-7612,32'd1169,32'd-1227,32'd3991,32'd3486,32'd709,32'd3200,32'd-4284,32'd6293,32'd-3056,32'd-140,32'd1784,32'd1599,32'd-99,32'd-3,32'd-2198,32'd-1106,32'd-4641,32'd968,32'd-2124,32'd3298,32'd4355,32'd-6591,32'd521,32'd5859,32'd1009,32'd-4101,32'd1056,32'd836,32'd-1999,32'd3095,32'd484,32'd-607,32'd1002,32'd-1479,32'd-8901,32'd1835,32'd8012,32'd4914,32'd1829,32'd-2792,32'd3154,32'd-1538,32'd-5278,32'd3364,32'd-1083,32'd1409,32'd4323,32'd532,32'd235,32'd-2418,32'd-8242,32'd1331,32'd5053,32'd6542,32'd5419,32'd-1409,32'd2315,32'd2083,32'd-1972,32'd-1132,32'd-1712,32'd5532,32'd1812,32'd-5185,32'd-1080,32'd13007,32'd-3173,32'd1425,32'd-1078,32'd-3068,32'd3327,32'd4733,32'd-4121,32'd5791,32'd-6083,32'd655,32'd2541,32'd1347,32'd-4396,32'd-1223,32'd3676,32'd10556,32'd-6308,32'd1285,32'd4257,32'd3056,32'd3757,32'd2331,32'd1679,32'd-7031,32'd-74,32'd-670,32'd2038,32'd-2246,32'd7856,32'd6123,32'd5883,32'd2792,32'd-28,32'd-931,32'd-1189,32'd-3408,32'd-881,32'd7172,32'd-3354,32'd5556,32'd1459,32'd8090,32'd-4145,32'd-4226,32'd1013,32'd-5864,32'd-5727,32'd-5395,32'd-401,32'd1750,32'd3967,32'd-6596,32'd-2382,32'd10859,32'd7158,32'd-420,32'd-3999,32'd311,32'd748,32'd-601,32'd-2275,32'd4921,32'd4938,32'd5654,32'd2658,32'd-1079,32'd-2008,32'd1877,32'd1102,32'd5737,32'd1073,32'd1077,32'd3916,32'd2822,32'd-745,32'd4304,32'd3928,32'd-1811,32'd551,32'd4284,32'd2939,32'd1807,32'd4924,32'd-1843,32'd-1765,32'd-4589,32'd-7163,32'd-3229,32'd7099,32'd-5566,32'd-599,32'd9262,32'd411};
    Wh[45]='{32'd3789,32'd-3420,32'd2875,32'd766,32'd1806,32'd-1651,32'd2221,32'd8383,32'd7285,32'd-543,32'd-6376,32'd-52,32'd36,32'd-625,32'd3464,32'd3908,32'd-1938,32'd-3427,32'd-5097,32'd581,32'd-1123,32'd1285,32'd-1035,32'd776,32'd127,32'd-6220,32'd611,32'd533,32'd2675,32'd-1157,32'd-449,32'd3681,32'd3842,32'd3515,32'd-2344,32'd-1419,32'd-1467,32'd653,32'd3554,32'd648,32'd-4086,32'd1553,32'd1073,32'd-562,32'd7504,32'd7236,32'd548,32'd6264,32'd-804,32'd-72,32'd-5092,32'd4350,32'd4951,32'd3784,32'd6186,32'd-2666,32'd2900,32'd-3430,32'd2453,32'd-6635,32'd-365,32'd530,32'd-1730,32'd-2209,32'd-798,32'd-3449,32'd220,32'd-947,32'd160,32'd-2437,32'd2452,32'd-1019,32'd1555,32'd-3652,32'd-1800,32'd2648,32'd5883,32'd-658,32'd1842,32'd-3740,32'd-315,32'd-259,32'd1741,32'd3037,32'd3474,32'd-53,32'd-1868,32'd-87,32'd6123,32'd938,32'd-614,32'd-5039,32'd-4438,32'd5239,32'd-4855,32'd654,32'd-1056,32'd-1193,32'd2133,32'd5112,32'd-2600,32'd-2880,32'd-2442,32'd-3132,32'd2829,32'd3154,32'd8457,32'd-196,32'd204,32'd947,32'd-2585,32'd-2336,32'd4804,32'd-2551,32'd-2937,32'd-3115,32'd5864,32'd-6240,32'd6801,32'd4101,32'd-2033,32'd-643,32'd9882,32'd3881,32'd-3740,32'd49,32'd-2524,32'd4250,32'd1723,32'd1162,32'd-716,32'd6206,32'd-5087,32'd4821,32'd2507,32'd1804,32'd3500,32'd-2700,32'd6083,32'd-3044,32'd-5493,32'd5073,32'd189,32'd-2230,32'd-2507,32'd648,32'd-9672,32'd7929,32'd1397,32'd-6752,32'd748,32'd-2592,32'd1943,32'd-3337,32'd-4042,32'd6572,32'd1639,32'd3386,32'd-8261,32'd-888,32'd3652,32'd-2707,32'd582,32'd4807,32'd869,32'd7177,32'd1437,32'd1139,32'd-3427,32'd-562,32'd-1264,32'd-1959,32'd-10966,32'd6601,32'd-8867,32'd-2426,32'd3146,32'd-1512,32'd5620,32'd-2322,32'd2034,32'd7573,32'd4523,32'd-7416,32'd-638,32'd-965,32'd794,32'd-2325,32'd-8344,32'd-2785,32'd1009,32'd6855,32'd1989,32'd6669,32'd383,32'd-2802,32'd-2687,32'd-1593,32'd-4636,32'd3444,32'd-4587,32'd-968,32'd3999,32'd-1898,32'd-846,32'd-2600,32'd4125,32'd-5756,32'd5791,32'd4233,32'd2368,32'd-38,32'd106,32'd128,32'd-2912,32'd-10957,32'd3867,32'd-5004,32'd1059,32'd13,32'd-895,32'd2543,32'd-2744,32'd-2457,32'd-938,32'd231,32'd-181,32'd1036,32'd-1883,32'd5488,32'd-984,32'd1109,32'd-3796,32'd-7685,32'd-4084,32'd-3371,32'd2851,32'd2805,32'd2144,32'd-3452,32'd3503,32'd-1970,32'd1406,32'd-2377,32'd-4389,32'd4470,32'd-783,32'd1412,32'd4770,32'd69,32'd-2307,32'd-4604,32'd-2470,32'd-3239,32'd5859,32'd-1096,32'd-4565,32'd236,32'd5380,32'd136,32'd6240,32'd3579,32'd-3178,32'd-200,32'd-2587,32'd-982,32'd-63,32'd3410,32'd1489,32'd390,32'd1040,32'd747,32'd-5249,32'd-243,32'd697,32'd-2602,32'd-2116,32'd4960,32'd2336,32'd105,32'd-1779,32'd625,32'd-52,32'd-5869,32'd-5039,32'd-1846,32'd2612,32'd432,32'd2827,32'd2609,32'd-2631,32'd-1987,32'd-503,32'd-1508,32'd4104,32'd6069,32'd204,32'd728,32'd279,32'd-2590,32'd-4150,32'd-9394,32'd1701,32'd1273,32'd1145,32'd-3276,32'd5849,32'd546,32'd3134,32'd-3393,32'd-2812,32'd-1054,32'd-2347,32'd1951,32'd985,32'd-6074,32'd-8994,32'd-3432,32'd8818,32'd3967,32'd-30,32'd695,32'd-1107,32'd1613,32'd3029,32'd-1650,32'd1812,32'd1213,32'd-3088,32'd-2302,32'd2636,32'd-3999,32'd4450,32'd-2504,32'd3410,32'd1839,32'd-2614,32'd2337,32'd-1204,32'd-3542,32'd3666,32'd-1162,32'd-1728,32'd292,32'd3,32'd-5747,32'd-272,32'd-1611,32'd4174,32'd-2476,32'd-7656,32'd-627,32'd3339,32'd3903,32'd2861,32'd442,32'd1285,32'd-2687,32'd-73,32'd-148,32'd3474,32'd-5019,32'd-1071,32'd-6494,32'd-5737,32'd-1783,32'd4824,32'd-5336,32'd473,32'd-8857,32'd-2619,32'd-1500,32'd-3608,32'd-1331,32'd3278,32'd-2492,32'd74,32'd-1800,32'd-836,32'd-72,32'd2731,32'd-3581,32'd2231,32'd1851,32'd-3833,32'd1782,32'd4489,32'd-1752,32'd3986,32'd9194,32'd-3862,32'd2878,32'd-985,32'd1275,32'd-5834,32'd466,32'd487,32'd-4804,32'd2885,32'd2846};
    Wh[46]='{32'd-116,32'd-1818,32'd-5136,32'd5087,32'd-6611,32'd-1828,32'd61,32'd-3500,32'd-416,32'd2301,32'd3947,32'd42,32'd-953,32'd-4050,32'd1193,32'd4130,32'd1925,32'd-5688,32'd147,32'd1617,32'd-3986,32'd-1569,32'd-2512,32'd-2242,32'd-2344,32'd-1667,32'd-608,32'd427,32'd-1794,32'd2464,32'd2120,32'd1461,32'd579,32'd-6772,32'd-8500,32'd-2189,32'd-3698,32'd-2169,32'd-2922,32'd429,32'd-1774,32'd-810,32'd1480,32'd2070,32'd-3845,32'd-3535,32'd5473,32'd-6723,32'd4091,32'd2116,32'd150,32'd-323,32'd-10302,32'd-432,32'd4550,32'd-14804,32'd-11191,32'd-4702,32'd-16,32'd-21972,32'd2587,32'd2854,32'd-1374,32'd-3337,32'd-1895,32'd3173,32'd-6230,32'd10390,32'd-791,32'd-4963,32'd-1729,32'd4465,32'd1914,32'd3884,32'd-1231,32'd1118,32'd-2971,32'd-4819,32'd2322,32'd4047,32'd1688,32'd-189,32'd-7407,32'd2741,32'd-5078,32'd1604,32'd1049,32'd2824,32'd-2902,32'd-811,32'd-2863,32'd2897,32'd835,32'd6137,32'd1430,32'd-2486,32'd-2147,32'd6772,32'd3942,32'd-1268,32'd3859,32'd1979,32'd3601,32'd-4562,32'd-2387,32'd414,32'd110,32'd4768,32'd-1303,32'd-7690,32'd1431,32'd-7651,32'd1767,32'd-1041,32'd2263,32'd-2368,32'd-1711,32'd4545,32'd-2130,32'd625,32'd1571,32'd8320,32'd8383,32'd3581,32'd-5742,32'd-4638,32'd-10117,32'd-9760,32'd4331,32'd289,32'd10234,32'd-2415,32'd2196,32'd-960,32'd4445,32'd-1,32'd-3879,32'd-6821,32'd-2358,32'd-16,32'd6508,32'd-824,32'd-180,32'd-1157,32'd1306,32'd-1522,32'd1732,32'd-2309,32'd-8198,32'd-6743,32'd3364,32'd-54,32'd-5156,32'd-3554,32'd-545,32'd6508,32'd-1605,32'd3110,32'd1929,32'd7670,32'd-740,32'd1571,32'd-3054,32'd-5112,32'd800,32'd-3750,32'd-3132,32'd-697,32'd-1564,32'd-3254,32'd5839,32'd-2076,32'd-1535,32'd-4416,32'd-1506,32'd3215,32'd3298,32'd-1540,32'd183,32'd5029,32'd123,32'd1601,32'd-1496,32'd3464,32'd-3298,32'd-663,32'd1211,32'd8793,32'd9628,32'd-450,32'd-7099,32'd2993,32'd5751,32'd725,32'd-2973,32'd8071,32'd4787,32'd-2829,32'd-4111,32'd-7377,32'd2207,32'd6328,32'd4389,32'd5537,32'd-5258,32'd2993,32'd-2143,32'd-1545,32'd-3022,32'd-7353,32'd-949,32'd1259,32'd3933,32'd-2780,32'd219,32'd-2016,32'd5991,32'd3723,32'd-420,32'd8676,32'd-1173,32'd426,32'd-101,32'd-914,32'd6176,32'd-5927,32'd3395,32'd-4067,32'd-5048,32'd911,32'd1665,32'd-2922,32'd-1992,32'd2514,32'd-2158,32'd1054,32'd-4047,32'd3066,32'd6855,32'd1888,32'd-3825,32'd1227,32'd1359,32'd1809,32'd-2252,32'd2291,32'd-417,32'd94,32'd3381,32'd2285,32'd-3337,32'd-5571,32'd2670,32'd-1638,32'd3798,32'd9541,32'd-302,32'd-7421,32'd241,32'd-4707,32'd-580,32'd-4396,32'd6894,32'd4143,32'd-2783,32'd-671,32'd-4533,32'd-6567,32'd-4995,32'd699,32'd-1030,32'd-7143,32'd-2198,32'd-1199,32'd-255,32'd-668,32'd2314,32'd-3596,32'd1572,32'd217,32'd-6860,32'd-1143,32'd3256,32'd-8417,32'd4584,32'd-3310,32'd2340,32'd-2866,32'd-484,32'd401,32'd7368,32'd5092,32'd2360,32'd-952,32'd-383,32'd-2049,32'd3227,32'd223,32'd-7255,32'd342,32'd-2059,32'd-765,32'd-8120,32'd-4675,32'd-2746,32'd-1174,32'd-3715,32'd74,32'd-181,32'd-1928,32'd7592,32'd2028,32'd2408,32'd-7524,32'd3295,32'd-1683,32'd3911,32'd1281,32'd-1229,32'd-256,32'd-4008,32'd2563,32'd815,32'd3171,32'd1250,32'd-361,32'd1260,32'd-1192,32'd-1291,32'd967,32'd-4155,32'd-704,32'd9331,32'd-3154,32'd3134,32'd5244,32'd4987,32'd4155,32'd-794,32'd-1892,32'd-2454,32'd-858,32'd-1964,32'd-5053,32'd-2880,32'd559,32'd9375,32'd2496,32'd1602,32'd-1010,32'd-4182,32'd-4611,32'd-3237,32'd-4011,32'd8583,32'd4406,32'd2141,32'd-2829,32'd-91,32'd2010,32'd1335,32'd-107,32'd129,32'd-3637,32'd-1199,32'd4729,32'd-5249,32'd2883,32'd509,32'd-846,32'd-5073,32'd3544,32'd-7880,32'd-5615,32'd2568,32'd-1932,32'd1352,32'd-3044,32'd1157,32'd7158,32'd-932,32'd204,32'd10283,32'd-5986,32'd-4731,32'd2736,32'd-3503,32'd-6669,32'd860,32'd1262,32'd-870,32'd200,32'd-3476,32'd144,32'd-1489,32'd-233,32'd-3359,32'd-9199,32'd2119,32'd1873};
    Wh[47]='{32'd-6025,32'd5302,32'd-1981,32'd4028,32'd3371,32'd-1656,32'd8037,32'd427,32'd1095,32'd2058,32'd4055,32'd-637,32'd-678,32'd1579,32'd3942,32'd1254,32'd-426,32'd5307,32'd-3774,32'd-3225,32'd1513,32'd2324,32'd-2395,32'd3666,32'd-4282,32'd2028,32'd1259,32'd1109,32'd1333,32'd-3859,32'd-4953,32'd-699,32'd-5761,32'd2592,32'd4179,32'd2110,32'd-1347,32'd-1020,32'd2263,32'd971,32'd-244,32'd437,32'd-1634,32'd2985,32'd650,32'd600,32'd698,32'd-2319,32'd-3662,32'd-1838,32'd1213,32'd2399,32'd4589,32'd2607,32'd124,32'd398,32'd436,32'd1844,32'd1710,32'd2147,32'd44,32'd5644,32'd-1760,32'd878,32'd-1926,32'd-1502,32'd3840,32'd1070,32'd-3730,32'd-3693,32'd-690,32'd2495,32'd-2714,32'd1632,32'd121,32'd-7812,32'd-3776,32'd444,32'd-3740,32'd2561,32'd-664,32'd2932,32'd-4042,32'd-3613,32'd-1408,32'd-1253,32'd-3220,32'd1320,32'd3293,32'd3225,32'd-3850,32'd-1118,32'd-3083,32'd-2266,32'd-393,32'd3227,32'd4272,32'd5405,32'd-1417,32'd26,32'd384,32'd3618,32'd1685,32'd-3952,32'd-40,32'd944,32'd3562,32'd-3879,32'd4895,32'd-112,32'd3830,32'd4887,32'd7875,32'd4179,32'd-1749,32'd900,32'd-4987,32'd4721,32'd4348,32'd1685,32'd-1960,32'd3168,32'd-3793,32'd-1210,32'd5141,32'd-2297,32'd-670,32'd-2011,32'd-1995,32'd-2207,32'd3679,32'd2724,32'd-195,32'd-2795,32'd1057,32'd-1078,32'd9096,32'd-2102,32'd1916,32'd-5434,32'd-2919,32'd1898,32'd-6992,32'd986,32'd-268,32'd7343,32'd5253,32'd-3959,32'd-1384,32'd1687,32'd2695,32'd192,32'd4372,32'd6708,32'd585,32'd-3330,32'd-2805,32'd377,32'd-2438,32'd-2917,32'd832,32'd5727,32'd-517,32'd3513,32'd2216,32'd314,32'd-1435,32'd1538,32'd-3957,32'd573,32'd-1096,32'd892,32'd-1684,32'd1254,32'd-2619,32'd1998,32'd-1245,32'd-1472,32'd5112,32'd-7104,32'd5615,32'd-2401,32'd1507,32'd-5922,32'd5444,32'd1860,32'd-2900,32'd4777,32'd-2418,32'd-4423,32'd632,32'd753,32'd-2432,32'd-3244,32'd780,32'd5395,32'd-332,32'd-201,32'd-2106,32'd2121,32'd1173,32'd-3879,32'd396,32'd-4692,32'd-2304,32'd-2531,32'd-1298,32'd-2261,32'd4375,32'd822,32'd-964,32'd-2282,32'd-3273,32'd-747,32'd-1979,32'd5898,32'd-1718,32'd1755,32'd-6005,32'd-1137,32'd-748,32'd3491,32'd-102,32'd-339,32'd2978,32'd-766,32'd1464,32'd-590,32'd440,32'd1842,32'd-6386,32'd-2213,32'd2548,32'd-1751,32'd-2529,32'd-1678,32'd5727,32'd-4592,32'd-2081,32'd1409,32'd-3410,32'd-1680,32'd760,32'd-3283,32'd-957,32'd-1741,32'd891,32'd-11103,32'd-5180,32'd3015,32'd-777,32'd4038,32'd1729,32'd-2364,32'd1196,32'd46,32'd-3896,32'd633,32'd-825,32'd-2812,32'd5756,32'd1928,32'd-659,32'd5419,32'd4284,32'd-1516,32'd-1529,32'd-1868,32'd1468,32'd-7031,32'd1040,32'd-1253,32'd2512,32'd-980,32'd5419,32'd2137,32'd2634,32'd-1640,32'd1230,32'd1759,32'd4257,32'd-903,32'd-1018,32'd5415,32'd-4531,32'd359,32'd-4521,32'd-2568,32'd5366,32'd-3051,32'd872,32'd-3056,32'd-1728,32'd-6635,32'd-689,32'd1743,32'd-4257,32'd5634,32'd-9101,32'd-5600,32'd-4565,32'd4050,32'd-794,32'd-1207,32'd-5009,32'd-1433,32'd-4450,32'd-3989,32'd2252,32'd-4523,32'd-2321,32'd-4765,32'd3842,32'd-2403,32'd-353,32'd-339,32'd-3254,32'd-4274,32'd-3698,32'd3208,32'd-347,32'd5161,32'd-5278,32'd4714,32'd3017,32'd2354,32'd1962,32'd-249,32'd3454,32'd-64,32'd1759,32'd6323,32'd-331,32'd789,32'd-3725,32'd5092,32'd-1293,32'd-2807,32'd-1933,32'd420,32'd-2785,32'd3908,32'd1475,32'd-434,32'd-2447,32'd-2900,32'd-853,32'd-4741,32'd-4035,32'd-2026,32'd-2553,32'd-824,32'd1055,32'd2226,32'd-4770,32'd-3395,32'd-4990,32'd-5029,32'd828,32'd-2333,32'd-701,32'd-8310,32'd-5415,32'd2095,32'd-2489,32'd3088,32'd4353,32'd2993,32'd721,32'd-385,32'd-4230,32'd-62,32'd-701,32'd362,32'd9570,32'd1304,32'd4111,32'd-2205,32'd-569,32'd-1992,32'd99,32'd-1254,32'd5532,32'd1525,32'd-1194,32'd-3068,32'd-4294,32'd-6474,32'd-1578,32'd-601,32'd3776,32'd-1789,32'd-2829,32'd-1052,32'd-7338,32'd917,32'd4880,32'd-3813,32'd-839,32'd-499};
    Wh[48]='{32'd532,32'd1602,32'd1838,32'd-5200,32'd-508,32'd596,32'd-984,32'd8100,32'd-3276,32'd723,32'd-247,32'd-670,32'd3825,32'd-3142,32'd-3867,32'd2198,32'd-154,32'd-1978,32'd-35,32'd3847,32'd455,32'd-1553,32'd-399,32'd-608,32'd-1730,32'd5229,32'd-770,32'd-1015,32'd2580,32'd-2922,32'd1381,32'd2661,32'd715,32'd-1461,32'd1318,32'd-1043,32'd-4274,32'd-1600,32'd4057,32'd-548,32'd-631,32'd-6401,32'd2795,32'd2612,32'd6723,32'd2327,32'd-1473,32'd4162,32'd-247,32'd-2717,32'd-1817,32'd1461,32'd-3417,32'd2395,32'd-861,32'd3845,32'd-781,32'd-1885,32'd1691,32'd7402,32'd3427,32'd5410,32'd-2468,32'd-265,32'd-6772,32'd805,32'd1002,32'd183,32'd4797,32'd1464,32'd-1712,32'd3996,32'd1074,32'd-2714,32'd2590,32'd1838,32'd-2871,32'd842,32'd4538,32'd3227,32'd-1687,32'd-1401,32'd-1302,32'd-1765,32'd2814,32'd-852,32'd2502,32'd-3691,32'd-524,32'd3303,32'd1722,32'd7172,32'd2192,32'd-124,32'd4377,32'd-532,32'd47,32'd-1840,32'd60,32'd3383,32'd-4472,32'd2031,32'd-2648,32'd-1447,32'd2478,32'd-190,32'd-6064,32'd183,32'd-9218,32'd1754,32'd-2340,32'd-1039,32'd-8657,32'd-181,32'd-6787,32'd6552,32'd4233,32'd-13027,32'd-29,32'd-488,32'd-798,32'd-725,32'd9921,32'd-2954,32'd-1621,32'd1568,32'd755,32'd-698,32'd3857,32'd2239,32'd-3129,32'd-690,32'd-6,32'd3520,32'd2298,32'd474,32'd55,32'd2100,32'd3859,32'd2218,32'd-5424,32'd-443,32'd4079,32'd2447,32'd753,32'd-1467,32'd-3869,32'd3015,32'd-8872,32'd142,32'd-5458,32'd957,32'd-1166,32'd-3720,32'd1538,32'd-4909,32'd5493,32'd-2191,32'd5844,32'd9409,32'd-2250,32'd-1761,32'd3464,32'd-3339,32'd6352,32'd-2512,32'd-2310,32'd-401,32'd-1157,32'd2056,32'd996,32'd2976,32'd7910,32'd3024,32'd1512,32'd-2912,32'd-1040,32'd-1525,32'd3701,32'd6264,32'd2797,32'd3684,32'd-1245,32'd991,32'd5566,32'd-78,32'd1820,32'd-7861,32'd-2592,32'd-1311,32'd-1273,32'd-659,32'd4294,32'd3164,32'd2143,32'd2045,32'd-5219,32'd1329,32'd5688,32'd-2524,32'd-1246,32'd4318,32'd-1397,32'd-3872,32'd3015,32'd-368,32'd4343,32'd-5454,32'd-3608,32'd239,32'd3132,32'd1557,32'd-4565,32'd617,32'd1217,32'd-6015,32'd-1436,32'd-6191,32'd4411,32'd-76,32'd-614,32'd-1701,32'd5258,32'd-7309,32'd-3342,32'd-1329,32'd-144,32'd293,32'd-3085,32'd474,32'd-1038,32'd4387,32'd121,32'd-783,32'd2612,32'd-2322,32'd-282,32'd1403,32'd-765,32'd304,32'd-3913,32'd-799,32'd357,32'd6752,32'd1574,32'd1347,32'd-1734,32'd298,32'd2641,32'd-364,32'd5878,32'd4199,32'd-1370,32'd2185,32'd-5014,32'd-9296,32'd-320,32'd-151,32'd573,32'd-2963,32'd-58,32'd-4729,32'd-2675,32'd-790,32'd604,32'd1253,32'd-2500,32'd414,32'd2712,32'd-439,32'd-283,32'd-4284,32'd5405,32'd2209,32'd-1811,32'd-3833,32'd345,32'd2563,32'd-2308,32'd1905,32'd-4462,32'd9326,32'd-657,32'd6220,32'd1699,32'd827,32'd1221,32'd5073,32'd2319,32'd-2312,32'd-8549,32'd328,32'd-1106,32'd5815,32'd6347,32'd1779,32'd2578,32'd-3471,32'd394,32'd-49,32'd-3010,32'd-10097,32'd-4169,32'd-4006,32'd-798,32'd-4528,32'd-4826,32'd3332,32'd1541,32'd182,32'd-522,32'd-1342,32'd584,32'd3654,32'd-218,32'd-1214,32'd2274,32'd-2368,32'd3083,32'd-1372,32'd-588,32'd2329,32'd2331,32'd2602,32'd-2565,32'd6899,32'd-2390,32'd-983,32'd2239,32'd7329,32'd-2729,32'd-4741,32'd-340,32'd-1156,32'd2285,32'd-4946,32'd5039,32'd-6337,32'd5166,32'd-4023,32'd-3405,32'd-2382,32'd-621,32'd-1213,32'd-167,32'd-1912,32'd7919,32'd3310,32'd2009,32'd-953,32'd3803,32'd741,32'd-3596,32'd-224,32'd-20,32'd7846,32'd2392,32'd3110,32'd-4184,32'd-4855,32'd2145,32'd84,32'd484,32'd-2064,32'd-1705,32'd-1412,32'd-2937,32'd-123,32'd-609,32'd-5068,32'd3181,32'd366,32'd-2626,32'd-6206,32'd-6303,32'd1328,32'd-1330,32'd-2448,32'd1656,32'd1779,32'd-6718,32'd621,32'd-888,32'd2437,32'd-3376,32'd1241,32'd1674,32'd1672,32'd2199,32'd646,32'd-3513,32'd728,32'd-1170,32'd-5532,32'd-1215,32'd2043,32'd-83,32'd4995,32'd1979,32'd1546};
    Wh[49]='{32'd-2374,32'd-1043,32'd729,32'd-484,32'd1795,32'd-838,32'd-781,32'd689,32'd-1865,32'd1262,32'd5361,32'd2995,32'd2600,32'd1668,32'd2032,32'd-2971,32'd682,32'd-383,32'd-2651,32'd830,32'd1282,32'd78,32'd89,32'd-499,32'd425,32'd5659,32'd505,32'd-726,32'd50,32'd617,32'd5820,32'd1936,32'd1607,32'd2156,32'd-1079,32'd664,32'd2770,32'd1776,32'd1496,32'd4138,32'd77,32'd-1574,32'd3317,32'd1582,32'd3435,32'd-1579,32'd320,32'd1130,32'd924,32'd-2758,32'd-1669,32'd-2171,32'd-2766,32'd-4228,32'd2111,32'd-2341,32'd1970,32'd326,32'd1695,32'd848,32'd-202,32'd-1761,32'd1884,32'd-707,32'd-883,32'd-3696,32'd-481,32'd1256,32'd1069,32'd-49,32'd2282,32'd1547,32'd-302,32'd-825,32'd932,32'd-256,32'd-3261,32'd3049,32'd1389,32'd2404,32'd316,32'd2141,32'd-864,32'd1354,32'd628,32'd-270,32'd1198,32'd-181,32'd1010,32'd428,32'd1176,32'd1216,32'd4514,32'd3149,32'd4562,32'd197,32'd-142,32'd308,32'd1052,32'd2656,32'd204,32'd-1357,32'd-1416,32'd-304,32'd3142,32'd-542,32'd287,32'd-379,32'd435,32'd-3022,32'd-4458,32'd-3315,32'd4670,32'd-669,32'd325,32'd161,32'd4440,32'd-1156,32'd2932,32'd-1512,32'd-2440,32'd-1031,32'd-3515,32'd825,32'd711,32'd6791,32'd-2092,32'd1339,32'd-2585,32'd-387,32'd-252,32'd-2937,32'd-86,32'd1932,32'd579,32'd-1583,32'd-458,32'd-3076,32'd55,32'd-952,32'd1166,32'd211,32'd1390,32'd1569,32'd-3647,32'd-3437,32'd-327,32'd657,32'd-1582,32'd-6347,32'd-2203,32'd-28,32'd5200,32'd2133,32'd-1889,32'd-319,32'd2546,32'd91,32'd4138,32'd996,32'd-2238,32'd2009,32'd-588,32'd1677,32'd-703,32'd995,32'd-1372,32'd1676,32'd957,32'd3122,32'd201,32'd1107,32'd-2,32'd545,32'd-482,32'd419,32'd-555,32'd3012,32'd-3427,32'd2257,32'd-1274,32'd-1191,32'd1971,32'd-1105,32'd-276,32'd2280,32'd748,32'd3049,32'd-837,32'd-3776,32'd-490,32'd251,32'd-2873,32'd1741,32'd-3479,32'd-1074,32'd2734,32'd-1145,32'd781,32'd166,32'd-866,32'd1372,32'd1300,32'd2622,32'd5820,32'd-372,32'd612,32'd-5,32'd516,32'd572,32'd-514,32'd886,32'd31,32'd1660,32'd-2049,32'd945,32'd-1340,32'd922,32'd1545,32'd3666,32'd1083,32'd-1437,32'd945,32'd1140,32'd-2081,32'd617,32'd4025,32'd-3112,32'd4843,32'd-1290,32'd-3046,32'd1418,32'd834,32'd585,32'd2333,32'd-800,32'd1312,32'd1468,32'd3366,32'd4016,32'd-1754,32'd1354,32'd-3269,32'd1381,32'd2575,32'd1767,32'd126,32'd3256,32'd-3173,32'd-617,32'd-2154,32'd-1995,32'd-7456,32'd4570,32'd1661,32'd1046,32'd5371,32'd4272,32'd2148,32'd1459,32'd1918,32'd4113,32'd-3000,32'd1043,32'd1517,32'd51,32'd1983,32'd4101,32'd2614,32'd-112,32'd1285,32'd1322,32'd-1566,32'd-1055,32'd849,32'd38,32'd-258,32'd1154,32'd182,32'd-2700,32'd3244,32'd2993,32'd5000,32'd2355,32'd885,32'd1374,32'd288,32'd7543,32'd1343,32'd-1685,32'd-2661,32'd1003,32'd775,32'd-451,32'd1430,32'd5297,32'd657,32'd1884,32'd390,32'd-1077,32'd2384,32'd3845,32'd79,32'd3793,32'd583,32'd1173,32'd-563,32'd17,32'd3352,32'd-2386,32'd1883,32'd-1193,32'd-3186,32'd2285,32'd3933,32'd485,32'd5258,32'd-606,32'd1759,32'd997,32'd-572,32'd527,32'd-751,32'd-913,32'd-2313,32'd3032,32'd-3742,32'd3825,32'd1315,32'd2471,32'd-536,32'd3032,32'd805,32'd-2258,32'd3969,32'd2939,32'd1489,32'd1934,32'd1932,32'd328,32'd2575,32'd-892,32'd4858,32'd936,32'd-1395,32'd-53,32'd3212,32'd-663,32'd1574,32'd-2639,32'd578,32'd2836,32'd-3298,32'd3708,32'd-1782,32'd2031,32'd59,32'd-1138,32'd-3383,32'd767,32'd1508,32'd3862,32'd3083,32'd4221,32'd-3823,32'd-1971,32'd295,32'd2288,32'd2890,32'd2042,32'd-6259,32'd-585,32'd1177,32'd2091,32'd1010,32'd4028,32'd-1505,32'd-115,32'd-7519,32'd-1160,32'd4763,32'd4216,32'd248,32'd1287,32'd444,32'd817,32'd-235,32'd2390,32'd1394,32'd-1179,32'd-460,32'd3461,32'd-992,32'd253,32'd1195,32'd-648,32'd3500,32'd-1423,32'd-703,32'd1273};
    Wh[50]='{32'd-1906,32'd-2778,32'd-2529,32'd-4387,32'd1053,32'd-2426,32'd-2722,32'd-639,32'd-6098,32'd-2330,32'd-8300,32'd-4743,32'd7128,32'd-5146,32'd73,32'd-9995,32'd-4362,32'd-8105,32'd625,32'd2182,32'd-638,32'd1352,32'd-335,32'd-1049,32'd-1108,32'd772,32'd-153,32'd-1237,32'd-2351,32'd-1503,32'd-1038,32'd-1816,32'd-5561,32'd-1619,32'd-1555,32'd5458,32'd-1284,32'd982,32'd165,32'd2144,32'd3752,32'd-1070,32'd4023,32'd-82,32'd4460,32'd-2636,32'd-8422,32'd4235,32'd458,32'd2414,32'd3623,32'd-4738,32'd8652,32'd1588,32'd-6059,32'd-4895,32'd-547,32'd3002,32'd3208,32'd-2229,32'd-1702,32'd1990,32'd-4328,32'd-455,32'd-5234,32'd-3610,32'd585,32'd1492,32'd-1274,32'd-1350,32'd1405,32'd4895,32'd-167,32'd-1795,32'd-3447,32'd-3513,32'd-705,32'd-5297,32'd483,32'd-2497,32'd-4926,32'd-305,32'd-2751,32'd1697,32'd-6748,32'd-2059,32'd-675,32'd-369,32'd2558,32'd3674,32'd7163,32'd1379,32'd2797,32'd360,32'd684,32'd-1666,32'd3994,32'd2861,32'd-235,32'd-4565,32'd1416,32'd-1516,32'd-427,32'd-2514,32'd3266,32'd-1690,32'd160,32'd-526,32'd4704,32'd-1544,32'd7353,32'd-784,32'd2885,32'd2009,32'd-7416,32'd884,32'd3803,32'd3659,32'd573,32'd465,32'd2303,32'd12558,32'd830,32'd4687,32'd-4780,32'd-11601,32'd8920,32'd-3918,32'd-6743,32'd4455,32'd5390,32'd-1916,32'd-7944,32'd2220,32'd-3186,32'd3901,32'd1638,32'd1319,32'd2666,32'd1885,32'd-4194,32'd-362,32'd-11875,32'd-5688,32'd-2479,32'd4743,32'd617,32'd3725,32'd-1588,32'd-2285,32'd-5273,32'd-320,32'd1134,32'd12783,32'd-1679,32'd4072,32'd-1500,32'd-2277,32'd-5581,32'd-6000,32'd-4448,32'd-102,32'd-3137,32'd-7446,32'd1,32'd6464,32'd4357,32'd4997,32'd-2399,32'd3359,32'd2156,32'd2658,32'd2293,32'd-2137,32'd3937,32'd319,32'd2814,32'd-5917,32'd5268,32'd-7734,32'd-495,32'd2001,32'd-1296,32'd2551,32'd-1447,32'd-602,32'd-1361,32'd-44,32'd-6953,32'd-845,32'd967,32'd-1958,32'd-10361,32'd3608,32'd-5664,32'd8725,32'd2073,32'd2416,32'd8549,32'd2521,32'd778,32'd3178,32'd-4052,32'd-4450,32'd1124,32'd3012,32'd2829,32'd5312,32'd-5952,32'd-491,32'd-1431,32'd-586,32'd-4111,32'd-264,32'd-2883,32'd1445,32'd3505,32'd2524,32'd527,32'd-6269,32'd3903,32'd6250,32'd7319,32'd-2003,32'd-9702,32'd1898,32'd5009,32'd-1137,32'd-1571,32'd6728,32'd-4475,32'd8886,32'd-3491,32'd-756,32'd-3137,32'd-3293,32'd-1529,32'd1508,32'd975,32'd-12763,32'd-4333,32'd-1802,32'd-2614,32'd-1057,32'd-2817,32'd4450,32'd-4099,32'd2022,32'd-910,32'd1209,32'd4973,32'd3664,32'd2465,32'd-4982,32'd2910,32'd8842,32'd-4768,32'd-4885,32'd4985,32'd7368,32'd-3808,32'd-3923,32'd-673,32'd-2348,32'd-5292,32'd-1796,32'd3259,32'd194,32'd-2304,32'd-365,32'd-1242,32'd-4616,32'd-6440,32'd-2741,32'd-5126,32'd-3527,32'd1616,32'd-1346,32'd-399,32'd-797,32'd2883,32'd-4843,32'd2553,32'd-1173,32'd7021,32'd8818,32'd1623,32'd-1907,32'd-6181,32'd1249,32'd4455,32'd4873,32'd-533,32'd-6865,32'd450,32'd4599,32'd-299,32'd-2939,32'd123,32'd-1427,32'd-1185,32'd-2268,32'd-2580,32'd-4956,32'd-6215,32'd-600,32'd-2548,32'd-3579,32'd-5341,32'd-6201,32'd2010,32'd-2824,32'd-2008,32'd-6469,32'd2381,32'd-6259,32'd-14638,32'd-8413,32'd-1839,32'd-2194,32'd-684,32'd567,32'd3083,32'd309,32'd-5283,32'd3063,32'd5390,32'd3156,32'd-4499,32'd2766,32'd-12226,32'd-4294,32'd-271,32'd-1079,32'd-1468,32'd-9965,32'd-2844,32'd2467,32'd-238,32'd-3964,32'd1817,32'd4802,32'd1507,32'd3259,32'd991,32'd-1807,32'd1712,32'd733,32'd-7294,32'd2230,32'd1710,32'd1798,32'd2321,32'd3701,32'd-4199,32'd-147,32'd-7128,32'd-9497,32'd11298,32'd-3713,32'd-583,32'd-7465,32'd2303,32'd-6752,32'd-5214,32'd2502,32'd3139,32'd-416,32'd1772,32'd-2401,32'd3547,32'd4335,32'd1572,32'd-5429,32'd1236,32'd-7827,32'd-4409,32'd-7270,32'd-1058,32'd-423,32'd6547,32'd-7075,32'd-1354,32'd-1351,32'd4345,32'd-7968,32'd-2714,32'd5937,32'd-3232,32'd3688,32'd-283,32'd-1828,32'd-2883,32'd541,32'd-3591,32'd812,32'd985,32'd-1550,32'd3029,32'd-1761};
    Wh[51]='{32'd4392,32'd114,32'd108,32'd858,32'd111,32'd395,32'd239,32'd-3786,32'd2315,32'd3686,32'd2651,32'd328,32'd1815,32'd1423,32'd29,32'd-1796,32'd8735,32'd-5502,32'd987,32'd2971,32'd254,32'd547,32'd3134,32'd2073,32'd-184,32'd5458,32'd-1099,32'd859,32'd394,32'd3493,32'd-3500,32'd-734,32'd5356,32'd-2373,32'd4216,32'd-1898,32'd-1012,32'd-616,32'd-3320,32'd3215,32'd794,32'd-6596,32'd1660,32'd3181,32'd-299,32'd-1650,32'd2187,32'd-4436,32'd2734,32'd-1315,32'd-6250,32'd-2617,32'd918,32'd-3764,32'd-4018,32'd619,32'd-661,32'd1408,32'd-1553,32'd3388,32'd1831,32'd3901,32'd-121,32'd-147,32'd2364,32'd-2575,32'd3208,32'd-1760,32'd1960,32'd3254,32'd-4768,32'd-814,32'd7924,32'd-6225,32'd-550,32'd-187,32'd-6928,32'd-637,32'd-3173,32'd1546,32'd-2255,32'd-4763,32'd2044,32'd-9116,32'd1896,32'd-3024,32'd250,32'd-1107,32'd-2088,32'd79,32'd1339,32'd-705,32'd4453,32'd2998,32'd-6723,32'd3830,32'd-914,32'd3586,32'd-928,32'd3178,32'd-5541,32'd771,32'd2164,32'd1187,32'd3764,32'd631,32'd-2065,32'd10527,32'd5180,32'd-2347,32'd4443,32'd2763,32'd2990,32'd-5073,32'd5146,32'd5678,32'd4492,32'd7890,32'd154,32'd-2697,32'd-897,32'd-3405,32'd1292,32'd-924,32'd1776,32'd-3359,32'd7714,32'd2780,32'd-3676,32'd-6362,32'd-3208,32'd-560,32'd-2866,32'd1459,32'd2128,32'd-921,32'd8256,32'd3337,32'd11406,32'd-1274,32'd-1828,32'd709,32'd16162,32'd4504,32'd-2391,32'd3952,32'd-1705,32'd-9672,32'd3740,32'd4948,32'd-1625,32'd-4465,32'd-339,32'd134,32'd5327,32'd-3264,32'd1435,32'd1704,32'd8168,32'd-375,32'd3972,32'd1363,32'd456,32'd2434,32'd-2399,32'd-6533,32'd-217,32'd6977,32'd-763,32'd-555,32'd-6210,32'd5136,32'd15175,32'd-2919,32'd-4306,32'd-327,32'd-878,32'd-3549,32'd2758,32'd-3188,32'd-9204,32'd3125,32'd2442,32'd1536,32'd-6650,32'd3410,32'd3447,32'd3857,32'd-5576,32'd-3942,32'd1348,32'd-2695,32'd-795,32'd3623,32'd-3449,32'd8432,32'd-3562,32'd-354,32'd3046,32'd3742,32'd90,32'd72,32'd-1206,32'd1751,32'd-3134,32'd-925,32'd3334,32'd-4860,32'd-7895,32'd1212,32'd2073,32'd3852,32'd4873,32'd1282,32'd3132,32'd775,32'd2780,32'd-1500,32'd-1756,32'd-358,32'd546,32'd-3173,32'd1840,32'd12,32'd-4843,32'd-385,32'd5253,32'd2183,32'd-1082,32'd1407,32'd2802,32'd1433,32'd-4255,32'd2812,32'd101,32'd-4101,32'd227,32'd186,32'd4929,32'd3051,32'd-2337,32'd4116,32'd5532,32'd-1345,32'd-2239,32'd1347,32'd3107,32'd-8886,32'd-1042,32'd1944,32'd-224,32'd5185,32'd2709,32'd25,32'd-1090,32'd1939,32'd3383,32'd8027,32'd-2019,32'd-1812,32'd-2854,32'd-831,32'd-385,32'd-6093,32'd330,32'd-1425,32'd5478,32'd-564,32'd-604,32'd-156,32'd180,32'd2030,32'd-1362,32'd-5747,32'd-1422,32'd-447,32'd-545,32'd-3698,32'd2993,32'd-3122,32'd1851,32'd4482,32'd4367,32'd-177,32'd-305,32'd6914,32'd-1773,32'd-265,32'd-5126,32'd-2211,32'd1425,32'd5483,32'd-1192,32'd-256,32'd5947,32'd-5449,32'd-904,32'd-2008,32'd6621,32'd405,32'd1646,32'd-3139,32'd5327,32'd-8125,32'd-2692,32'd-1193,32'd-5083,32'd5473,32'd1813,32'd-1413,32'd924,32'd3723,32'd-3125,32'd-6708,32'd-4941,32'd3095,32'd2651,32'd1538,32'd-3852,32'd-3625,32'd7836,32'd446,32'd2340,32'd-1940,32'd-3603,32'd6196,32'd-1635,32'd2231,32'd-3781,32'd3027,32'd1693,32'd3244,32'd-972,32'd545,32'd1287,32'd-9013,32'd-560,32'd3217,32'd-2961,32'd-362,32'd2303,32'd3833,32'd-351,32'd-3754,32'd-78,32'd5839,32'd-14589,32'd2924,32'd-5415,32'd2124,32'd2517,32'd-131,32'd4765,32'd1783,32'd2396,32'd4245,32'd5297,32'd-8666,32'd-886,32'd8232,32'd-1301,32'd3813,32'd-704,32'd1889,32'd2354,32'd3171,32'd1596,32'd-5224,32'd-1038,32'd-4790,32'd4565,32'd4191,32'd12041,32'd-7675,32'd-596,32'd4157,32'd5703,32'd1308,32'd1079,32'd933,32'd-1146,32'd2634,32'd-2932,32'd-1739,32'd1783,32'd-2548,32'd3527,32'd-3020,32'd-2934,32'd1932,32'd-194,32'd-1979,32'd-2333,32'd5742,32'd1331,32'd-196,32'd626,32'd-3728,32'd2905,32'd-1798};
    Wh[52]='{32'd2208,32'd-1138,32'd-121,32'd-7099,32'd-1254,32'd-810,32'd-685,32'd828,32'd-1516,32'd-2388,32'd-123,32'd-1776,32'd-561,32'd-2954,32'd-1920,32'd-6562,32'd-8,32'd-5078,32'd-1811,32'd-17,32'd2192,32'd155,32'd3527,32'd-2216,32'd-926,32'd417,32'd-1374,32'd-3808,32'd-3134,32'd-569,32'd-789,32'd-372,32'd-2326,32'd-1574,32'd-755,32'd-2158,32'd396,32'd-1416,32'd-2215,32'd-3649,32'd-1604,32'd-3305,32'd1367,32'd3325,32'd3508,32'd-5415,32'd-805,32'd4528,32'd-3852,32'd5708,32'd1247,32'd-1357,32'd122,32'd641,32'd3276,32'd2932,32'd1763,32'd4807,32'd-6381,32'd1322,32'd-2113,32'd-3605,32'd-2344,32'd-1010,32'd620,32'd1773,32'd1147,32'd-3977,32'd3239,32'd-1318,32'd6,32'd-6000,32'd-3879,32'd2191,32'd-5498,32'd-2958,32'd-3850,32'd-1937,32'd1585,32'd1319,32'd1527,32'd592,32'd2078,32'd-6625,32'd-1828,32'd-1380,32'd3630,32'd-1392,32'd3247,32'd4206,32'd-1893,32'd1549,32'd1376,32'd-2587,32'd1739,32'd1334,32'd-1687,32'd-6,32'd1011,32'd4082,32'd2288,32'd-2152,32'd-4848,32'd2105,32'd-2357,32'd758,32'd-1519,32'd-1459,32'd-3193,32'd3007,32'd313,32'd5878,32'd-3173,32'd3962,32'd2944,32'd776,32'd894,32'd-376,32'd-2919,32'd793,32'd35,32'd5693,32'd-1124,32'd4152,32'd-2387,32'd1473,32'd-38,32'd445,32'd-823,32'd5961,32'd-4699,32'd-882,32'd-1408,32'd4453,32'd6079,32'd115,32'd-1206,32'd580,32'd3291,32'd-1518,32'd-2463,32'd3234,32'd-2136,32'd2966,32'd1920,32'd-5913,32'd-4511,32'd7622,32'd-623,32'd4323,32'd1417,32'd5786,32'd-11279,32'd-7045,32'd-5253,32'd235,32'd4206,32'd117,32'd3728,32'd-2452,32'd-3310,32'd2257,32'd1118,32'd171,32'd-1733,32'd5170,32'd-3820,32'd-3112,32'd-1031,32'd-370,32'd-5156,32'd-2907,32'd1218,32'd-2178,32'd68,32'd-3776,32'd-96,32'd-167,32'd-6655,32'd-1290,32'd1418,32'd1101,32'd-2437,32'd317,32'd1252,32'd538,32'd-5756,32'd-5063,32'd-2382,32'd5317,32'd112,32'd2404,32'd-25,32'd2264,32'd-1540,32'd1502,32'd-520,32'd-599,32'd6494,32'd3837,32'd-889,32'd-1953,32'd2844,32'd2214,32'd-745,32'd3220,32'd1927,32'd3251,32'd3928,32'd0,32'd3703,32'd-682,32'd-7299,32'd-2441,32'd557,32'd2258,32'd-1212,32'd957,32'd764,32'd1002,32'd2006,32'd-10,32'd-1309,32'd-3093,32'd-3645,32'd-1516,32'd453,32'd592,32'd668,32'd-610,32'd1772,32'd-1181,32'd-2546,32'd739,32'd-573,32'd900,32'd-2746,32'd848,32'd1151,32'd4421,32'd-1807,32'd-1854,32'd4650,32'd3251,32'd-491,32'd141,32'd-759,32'd3051,32'd42,32'd895,32'd-2905,32'd3103,32'd-265,32'd3483,32'd-5424,32'd3002,32'd1138,32'd2536,32'd2147,32'd-1809,32'd866,32'd211,32'd-894,32'd3647,32'd2937,32'd2027,32'd-983,32'd-417,32'd2352,32'd1925,32'd-3437,32'd3288,32'd-3691,32'd-1628,32'd-1680,32'd986,32'd1938,32'd6054,32'd-5791,32'd-1518,32'd-1813,32'd-48,32'd938,32'd2457,32'd2214,32'd-2856,32'd1948,32'd-2580,32'd1558,32'd761,32'd-5249,32'd1390,32'd6694,32'd2186,32'd1317,32'd-572,32'd3647,32'd473,32'd-2469,32'd3288,32'd-6206,32'd1746,32'd-2893,32'd2243,32'd3063,32'd-1267,32'd644,32'd-2232,32'd437,32'd654,32'd-158,32'd-647,32'd5292,32'd-2181,32'd-1739,32'd-184,32'd2120,32'd1123,32'd-606,32'd-857,32'd1678,32'd414,32'd600,32'd-3559,32'd-2575,32'd-3222,32'd-1923,32'd233,32'd3884,32'd-7495,32'd-2076,32'd-224,32'd-440,32'd-2924,32'd3532,32'd-3256,32'd-3354,32'd-1013,32'd495,32'd-209,32'd4580,32'd-841,32'd2604,32'd2993,32'd1992,32'd2587,32'd1304,32'd995,32'd302,32'd-3820,32'd4484,32'd-4858,32'd-1900,32'd253,32'd-474,32'd-1279,32'd2666,32'd-7641,32'd-2094,32'd-2028,32'd-4711,32'd2349,32'd722,32'd2697,32'd-2687,32'd-7065,32'd-1434,32'd1558,32'd2495,32'd-5156,32'd2209,32'd-1770,32'd2275,32'd628,32'd-3503,32'd1004,32'd-2014,32'd1828,32'd-339,32'd1032,32'd-1619,32'd2047,32'd1734,32'd-136,32'd-52,32'd1888,32'd1915,32'd3281,32'd-1553,32'd175,32'd-1011,32'd-1126,32'd1094,32'd131,32'd-1754,32'd7192,32'd-681,32'd1195,32'd-3156,32'd861};
    Wh[53]='{32'd-3225,32'd-412,32'd-139,32'd939,32'd2181,32'd-1264,32'd-1662,32'd-1688,32'd575,32'd-203,32'd-3784,32'd-1734,32'd-789,32'd3923,32'd3513,32'd1665,32'd-127,32'd-2597,32'd-2529,32'd-1757,32'd-1983,32'd2556,32'd722,32'd4357,32'd-885,32'd6289,32'd310,32'd2459,32'd-5322,32'd-1028,32'd-1823,32'd-561,32'd3444,32'd268,32'd-892,32'd-2233,32'd598,32'd172,32'd3200,32'd1756,32'd-4921,32'd-2880,32'd-3962,32'd1771,32'd1948,32'd-1990,32'd-1676,32'd3596,32'd2257,32'd2397,32'd-1666,32'd1638,32'd2315,32'd5449,32'd7670,32'd2631,32'd1876,32'd-3005,32'd4826,32'd-3156,32'd-2427,32'd4792,32'd4758,32'd-5346,32'd-1990,32'd-1051,32'd-1972,32'd675,32'd-1628,32'd443,32'd5546,32'd4235,32'd-2546,32'd-2419,32'd-1826,32'd-3874,32'd4025,32'd860,32'd-167,32'd3999,32'd2153,32'd2490,32'd2868,32'd-2186,32'd2800,32'd-4719,32'd1767,32'd-1328,32'd-927,32'd169,32'd-5458,32'd5195,32'd-6865,32'd1248,32'd2568,32'd4208,32'd-779,32'd415,32'd769,32'd-2327,32'd8623,32'd4016,32'd-2800,32'd-249,32'd5273,32'd2032,32'd3078,32'd1102,32'd3186,32'd-2347,32'd-3862,32'd-6982,32'd-1535,32'd2181,32'd-3320,32'd-1401,32'd-360,32'd455,32'd8579,32'd3093,32'd-3159,32'd460,32'd-3537,32'd-5473,32'd2648,32'd8237,32'd-8315,32'd2178,32'd1368,32'd-87,32'd-224,32'd-3210,32'd-875,32'd-2301,32'd-2966,32'd701,32'd-3735,32'd1777,32'd2792,32'd87,32'd-1948,32'd4255,32'd7172,32'd-1376,32'd4860,32'd2336,32'd-1380,32'd6835,32'd-2014,32'd1409,32'd63,32'd-1510,32'd428,32'd-7211,32'd-1183,32'd3251,32'd-2272,32'd-3525,32'd-875,32'd3908,32'd-2368,32'd4807,32'd-1409,32'd6860,32'd-7646,32'd-92,32'd186,32'd1833,32'd2036,32'd-2379,32'd1701,32'd-954,32'd-7412,32'd-1560,32'd-3869,32'd2788,32'd-2243,32'd7690,32'd-1112,32'd-4003,32'd-525,32'd4506,32'd3881,32'd-2397,32'd-114,32'd-2619,32'd2668,32'd545,32'd-10400,32'd-903,32'd-1877,32'd1075,32'd-1036,32'd-6752,32'd-2304,32'd339,32'd2359,32'd877,32'd-4147,32'd-115,32'd-3308,32'd-760,32'd3134,32'd8354,32'd2717,32'd-99,32'd-4218,32'd2302,32'd-899,32'd-2951,32'd1710,32'd-5312,32'd-1564,32'd-178,32'd-4628,32'd-5141,32'd578,32'd-1667,32'd-3732,32'd-954,32'd-992,32'd7338,32'd-859,32'd-2012,32'd121,32'd1849,32'd857,32'd-1589,32'd-4931,32'd-3930,32'd2988,32'd-103,32'd1527,32'd869,32'd-5454,32'd435,32'd3845,32'd-385,32'd-1671,32'd-1628,32'd3925,32'd-4992,32'd-2529,32'd-4616,32'd-4658,32'd2585,32'd-3332,32'd-439,32'd-1840,32'd1178,32'd-2176,32'd-4968,32'd245,32'd2003,32'd-610,32'd2595,32'd2277,32'd-1434,32'd345,32'd1341,32'd1011,32'd-4604,32'd-2573,32'd-3879,32'd-23,32'd1084,32'd-2425,32'd-1572,32'd-3852,32'd3737,32'd244,32'd6005,32'd-223,32'd-333,32'd389,32'd-2915,32'd-2651,32'd-1006,32'd107,32'd1582,32'd-4616,32'd1402,32'd-6899,32'd1209,32'd-1795,32'd-2406,32'd788,32'd-3864,32'd51,32'd-1043,32'd3493,32'd989,32'd-652,32'd-460,32'd-2658,32'd-673,32'd-2418,32'd-124,32'd162,32'd-3754,32'd-4313,32'd-514,32'd3076,32'd1136,32'd1172,32'd3032,32'd-1284,32'd-6352,32'd859,32'd-1633,32'd-2055,32'd4257,32'd-3066,32'd-2824,32'd3728,32'd4223,32'd-313,32'd-2177,32'd1712,32'd6528,32'd6313,32'd1961,32'd-5698,32'd1065,32'd-1361,32'd4301,32'd-828,32'd4777,32'd-1380,32'd67,32'd-342,32'd-2888,32'd-263,32'd-747,32'd-718,32'd1528,32'd1616,32'd4450,32'd1796,32'd1910,32'd3706,32'd-401,32'd1187,32'd-2198,32'd-5517,32'd-466,32'd-643,32'd-4165,32'd2220,32'd-1177,32'd-1242,32'd3901,32'd-2578,32'd5175,32'd4599,32'd-3786,32'd-1500,32'd2932,32'd-3073,32'd684,32'd745,32'd-3779,32'd-3513,32'd4604,32'd-11679,32'd6669,32'd4206,32'd-793,32'd-774,32'd6435,32'd578,32'd-1276,32'd-2963,32'd5107,32'd-1372,32'd-4177,32'd-601,32'd-3417,32'd263,32'd-127,32'd1100,32'd-2373,32'd2496,32'd-1531,32'd406,32'd-2042,32'd3764,32'd-3024,32'd2211,32'd3991,32'd-2590,32'd360,32'd1386,32'd-651,32'd-3913,32'd-1131,32'd5395,32'd-6030,32'd871,32'd256};
    Wh[54]='{32'd4870,32'd6557,32'd1606,32'd5068,32'd3947,32'd-745,32'd1873,32'd2971,32'd4062,32'd3554,32'd-578,32'd1394,32'd3671,32'd2418,32'd3173,32'd-2441,32'd733,32'd3730,32'd2758,32'd3149,32'd2042,32'd2012,32'd1040,32'd2592,32'd593,32'd-236,32'd2340,32'd-622,32'd-278,32'd6088,32'd6010,32'd1108,32'd4101,32'd4824,32'd-6323,32'd2607,32'd4506,32'd2519,32'd-1264,32'd1579,32'd7182,32'd452,32'd10351,32'd-307,32'd8315,32'd5214,32'd2724,32'd1706,32'd2113,32'd-4245,32'd781,32'd2983,32'd-2141,32'd3249,32'd1219,32'd4631,32'd4396,32'd491,32'd3020,32'd5092,32'd2629,32'd350,32'd-289,32'd4252,32'd-7832,32'd1940,32'd4538,32'd5288,32'd714,32'd-549,32'd503,32'd578,32'd4853,32'd2714,32'd4431,32'd9707,32'd9160,32'd4306,32'd416,32'd2851,32'd1667,32'd6733,32'd6254,32'd1821,32'd1268,32'd957,32'd-2188,32'd2436,32'd-7998,32'd-1539,32'd1387,32'd-520,32'd2116,32'd916,32'd1640,32'd4064,32'd-2536,32'd6967,32'd1884,32'd2509,32'd-6645,32'd3295,32'd2235,32'd14511,32'd423,32'd3730,32'd139,32'd-3691,32'd1105,32'd347,32'd2854,32'd-3945,32'd2937,32'd-822,32'd-3088,32'd7255,32'd7875,32'd11083,32'd1490,32'd2110,32'd-4123,32'd-913,32'd2415,32'd3100,32'd1118,32'd-1628,32'd1479,32'd4143,32'd-2082,32'd-7167,32'd2434,32'd2509,32'd-1436,32'd1823,32'd-501,32'd2844,32'd3374,32'd-5415,32'd1729,32'd260,32'd-1328,32'd-2912,32'd6381,32'd-4357,32'd4511,32'd-690,32'd-464,32'd-1859,32'd-3698,32'd2462,32'd2225,32'd3564,32'd-2849,32'd-5068,32'd2844,32'd6547,32'd6206,32'd2707,32'd1795,32'd11875,32'd8183,32'd1066,32'd-890,32'd-6440,32'd2985,32'd2399,32'd1917,32'd2553,32'd-100,32'd-3259,32'd1258,32'd4980,32'd-808,32'd-2058,32'd-3151,32'd-3054,32'd2746,32'd-4135,32'd2253,32'd-725,32'd-1730,32'd321,32'd-7963,32'd-504,32'd-8383,32'd563,32'd5317,32'd-4323,32'd93,32'd-6313,32'd5864,32'd-3305,32'd-3110,32'd-2546,32'd-3298,32'd-9946,32'd-6308,32'd267,32'd-5898,32'd1430,32'd-723,32'd-1237,32'd-2702,32'd-1573,32'd-1514,32'd-2187,32'd4572,32'd-276,32'd6293,32'd4333,32'd-2614,32'd3215,32'd6220,32'd118,32'd-952,32'd-577,32'd180,32'd7583,32'd3911,32'd993,32'd1392,32'd513,32'd1994,32'd1220,32'd1766,32'd1879,32'd708,32'd2054,32'd-1357,32'd2266,32'd3552,32'd-2465,32'd2181,32'd701,32'd-6806,32'd-5937,32'd3999,32'd128,32'd-310,32'd-4750,32'd762,32'd-2507,32'd-4841,32'd5776,32'd-2961,32'd1264,32'd1263,32'd-4501,32'd4753,32'd-795,32'd483,32'd-2459,32'd3933,32'd5556,32'd5058,32'd-463,32'd-888,32'd-3515,32'd6230,32'd3254,32'd3334,32'd5361,32'd-2893,32'd1057,32'd-2670,32'd-3234,32'd4553,32'd3962,32'd-1552,32'd-236,32'd2749,32'd208,32'd1737,32'd3903,32'd4028,32'd-1831,32'd-1855,32'd-2191,32'd930,32'd2231,32'd1510,32'd1529,32'd2385,32'd-1102,32'd-974,32'd6865,32'd2082,32'd1021,32'd5566,32'd-4157,32'd6801,32'd-50,32'd-724,32'd1238,32'd-1381,32'd-5278,32'd4174,32'd-7792,32'd-899,32'd3999,32'd7993,32'd-7714,32'd2836,32'd2878,32'd2242,32'd4348,32'd5419,32'd4421,32'd3564,32'd4675,32'd-37,32'd5273,32'd-1624,32'd5268,32'd575,32'd-1505,32'd-5717,32'd7592,32'd1577,32'd5898,32'd4699,32'd-664,32'd6640,32'd-1219,32'd13,32'd-2763,32'd-145,32'd2573,32'd-785,32'd4228,32'd4641,32'd1301,32'd-1578,32'd3359,32'd-1937,32'd231,32'd1391,32'd1044,32'd2954,32'd-9257,32'd3789,32'd-4335,32'd2924,32'd890,32'd5688,32'd-5551,32'd-1036,32'd4389,32'd1752,32'd2617,32'd-2418,32'd523,32'd-2480,32'd1788,32'd-1602,32'd70,32'd7412,32'd-3203,32'd2425,32'd-3620,32'd8422,32'd386,32'd364,32'd-2261,32'd1517,32'd7514,32'd7451,32'd-809,32'd-115,32'd-6386,32'd7236,32'd2536,32'd-192,32'd-4865,32'd3242,32'd-1914,32'd-472,32'd-1242,32'd2646,32'd3935,32'd4699,32'd1103,32'd3403,32'd-2846,32'd3916,32'd-4858,32'd4946,32'd3559,32'd1746,32'd315,32'd21,32'd3337,32'd4206,32'd-3574,32'd1745,32'd-7290,32'd870,32'd2407,32'd214,32'd1816};
    Wh[55]='{32'd3784,32'd5961,32'd3996,32'd-4636,32'd-2473,32'd-3364,32'd1242,32'd371,32'd-5668,32'd3200,32'd-1262,32'd-1768,32'd1109,32'd-1464,32'd3710,32'd741,32'd-58,32'd-3037,32'd1575,32'd180,32'd965,32'd159,32'd2495,32'd3090,32'd-5498,32'd3127,32'd-1227,32'd-2683,32'd-7319,32'd-1621,32'd3708,32'd502,32'd-2553,32'd4375,32'd-16660,32'd2225,32'd-10761,32'd6010,32'd3073,32'd-105,32'd9414,32'd4704,32'd2687,32'd546,32'd-797,32'd-3967,32'd-5112,32'd-2241,32'd145,32'd2457,32'd-2044,32'd1243,32'd251,32'd6328,32'd-1088,32'd-4104,32'd20,32'd2614,32'd-744,32'd-12041,32'd7705,32'd5361,32'd3684,32'd-4553,32'd-6357,32'd-875,32'd345,32'd-4733,32'd2995,32'd906,32'd-3977,32'd737,32'd2230,32'd-897,32'd2875,32'd809,32'd4658,32'd5825,32'd-2297,32'd-2003,32'd3269,32'd4975,32'd4765,32'd1896,32'd-154,32'd-2687,32'd940,32'd1480,32'd-441,32'd4230,32'd1605,32'd-635,32'd-468,32'd6357,32'd1411,32'd-797,32'd1738,32'd-1680,32'd1822,32'd1944,32'd-3383,32'd4870,32'd-2917,32'd-7797,32'd-4111,32'd3676,32'd5288,32'd2604,32'd-4509,32'd516,32'd-2663,32'd3708,32'd-2139,32'd2060,32'd-1269,32'd-3215,32'd938,32'd-3632,32'd-6083,32'd-1467,32'd-3342,32'd4895,32'd-1867,32'd-602,32'd-7207,32'd2526,32'd-616,32'd-2778,32'd-2900,32'd3645,32'd632,32'd-402,32'd5927,32'd3593,32'd15634,32'd-3957,32'd-6772,32'd6474,32'd-1669,32'd3630,32'd-6201,32'd-2277,32'd-1893,32'd1317,32'd-3256,32'd-4060,32'd-457,32'd3789,32'd5810,32'd3195,32'd-4645,32'd2407,32'd2624,32'd560,32'd-6562,32'd938,32'd1505,32'd-281,32'd2636,32'd11923,32'd-3437,32'd-543,32'd-184,32'd-4985,32'd-1916,32'd11162,32'd6811,32'd-2111,32'd206,32'd-1527,32'd-2443,32'd1130,32'd952,32'd1045,32'd1149,32'd1612,32'd4812,32'd-1195,32'd-3200,32'd-924,32'd-5,32'd-3881,32'd-3190,32'd3349,32'd-2807,32'd51,32'd1169,32'd1085,32'd-2404,32'd1179,32'd-6518,32'd-2198,32'd-3115,32'd-1287,32'd3505,32'd3684,32'd-428,32'd1019,32'd890,32'd6279,32'd1157,32'd-1308,32'd-1092,32'd-2415,32'd-4101,32'd-2006,32'd1162,32'd-264,32'd1687,32'd-5654,32'd-1749,32'd4377,32'd-5156,32'd2524,32'd-2775,32'd2127,32'd1684,32'd4328,32'd-562,32'd3132,32'd321,32'd1141,32'd-1434,32'd1457,32'd-2489,32'd2071,32'd2631,32'd-7529,32'd1539,32'd1606,32'd-2929,32'd-1125,32'd1152,32'd-2009,32'd4738,32'd-4631,32'd-4504,32'd-1386,32'd1126,32'd-4355,32'd-3242,32'd3469,32'd603,32'd5224,32'd-1634,32'd-424,32'd5249,32'd1993,32'd-1683,32'd2761,32'd4829,32'd655,32'd-2008,32'd-2746,32'd345,32'd-8276,32'd1232,32'd-3789,32'd-680,32'd5302,32'd-452,32'd-3415,32'd-4323,32'd6386,32'd265,32'd-333,32'd-5322,32'd2478,32'd2092,32'd220,32'd2229,32'd-6821,32'd2318,32'd-2114,32'd-1175,32'd-3552,32'd-2575,32'd-178,32'd-1146,32'd-2612,32'd2322,32'd-1748,32'd-5576,32'd-11806,32'd1233,32'd4548,32'd-443,32'd-7919,32'd-2841,32'd4599,32'd7172,32'd-3928,32'd3669,32'd7719,32'd-2871,32'd1842,32'd4013,32'd843,32'd354,32'd-700,32'd-1121,32'd1468,32'd7319,32'd143,32'd-3544,32'd-1383,32'd1549,32'd-3562,32'd-1483,32'd1612,32'd3559,32'd2257,32'd2110,32'd-1993,32'd-1149,32'd-8891,32'd2617,32'd7265,32'd4311,32'd-2783,32'd3217,32'd-2536,32'd3200,32'd-1550,32'd-2054,32'd4711,32'd2583,32'd2360,32'd-255,32'd-813,32'd-3686,32'd880,32'd-4565,32'd-2976,32'd983,32'd-7519,32'd-7387,32'd8344,32'd4978,32'd-722,32'd9658,32'd-1864,32'd5234,32'd961,32'd366,32'd-1606,32'd-457,32'd-4179,32'd-4489,32'd287,32'd3386,32'd-728,32'd648,32'd-3564,32'd5478,32'd-6665,32'd4208,32'd-4304,32'd2780,32'd-8095,32'd545,32'd-579,32'd2410,32'd-4753,32'd-3002,32'd-8339,32'd4809,32'd393,32'd-501,32'd1683,32'd-6162,32'd-1212,32'd-2266,32'd4204,32'd1993,32'd466,32'd3391,32'd-1590,32'd-1370,32'd5053,32'd303,32'd-8720,32'd2617,32'd512,32'd781,32'd31,32'd809,32'd1242,32'd-10576,32'd6381,32'd6342,32'd-882,32'd280,32'd-545,32'd2724,32'd3356,32'd-565,32'd481,32'd-3723,32'd-2624};
    Wh[56]='{32'd-112,32'd1662,32'd-1029,32'd-3530,32'd-2127,32'd-764,32'd1037,32'd-5024,32'd-138,32'd878,32'd-8637,32'd-1243,32'd-5083,32'd-2032,32'd3039,32'd-2331,32'd2863,32'd3283,32'd-848,32'd1407,32'd1867,32'd2279,32'd82,32'd-2902,32'd-3745,32'd1341,32'd-2514,32'd-1711,32'd343,32'd-1062,32'd-59,32'd-3649,32'd1007,32'd4240,32'd939,32'd-3925,32'd-1085,32'd-1148,32'd-327,32'd-398,32'd5668,32'd75,32'd636,32'd-2349,32'd-941,32'd2770,32'd1181,32'd-3918,32'd-803,32'd-148,32'd6464,32'd-2277,32'd-4582,32'd-3903,32'd-2534,32'd439,32'd-3166,32'd-2297,32'd999,32'd7202,32'd225,32'd-2751,32'd1756,32'd-3588,32'd-2369,32'd-2529,32'd-2225,32'd-344,32'd879,32'd403,32'd2451,32'd-4011,32'd412,32'd4167,32'd-413,32'd3664,32'd-5439,32'd138,32'd7036,32'd1001,32'd-1834,32'd8349,32'd4355,32'd-3662,32'd-575,32'd1693,32'd-1004,32'd-1056,32'd-96,32'd4082,32'd2465,32'd-3889,32'd-5087,32'd-4328,32'd-2291,32'd4594,32'd-2653,32'd-1649,32'd-2324,32'd1250,32'd1932,32'd-3164,32'd-526,32'd-949,32'd2824,32'd14,32'd-1176,32'd-11640,32'd1685,32'd-797,32'd183,32'd13867,32'd-7890,32'd791,32'd-45,32'd-2164,32'd-1706,32'd2438,32'd246,32'd-3911,32'd2963,32'd-4912,32'd5327,32'd5893,32'd-2500,32'd-5576,32'd-3125,32'd-4084,32'd6459,32'd-59,32'd4494,32'd-4489,32'd5625,32'd-245,32'd440,32'd-4580,32'd1322,32'd3439,32'd2700,32'd2119,32'd2827,32'd-3969,32'd-792,32'd-1799,32'd952,32'd527,32'd-3327,32'd-626,32'd1297,32'd-2629,32'd1636,32'd5039,32'd-4416,32'd3105,32'd0,32'd-405,32'd1446,32'd697,32'd-1182,32'd2165,32'd2946,32'd-4228,32'd-5576,32'd-898,32'd4716,32'd3835,32'd-1330,32'd370,32'd-5737,32'd2076,32'd-1990,32'd-4389,32'd-1586,32'd4289,32'd-847,32'd989,32'd736,32'd3630,32'd-971,32'd-44,32'd-2551,32'd-913,32'd-3596,32'd1467,32'd3330,32'd-2714,32'd1618,32'd7465,32'd4724,32'd2059,32'd6699,32'd-1422,32'd1994,32'd3964,32'd3640,32'd-4965,32'd-2041,32'd-2866,32'd-2335,32'd2490,32'd-1481,32'd829,32'd-1574,32'd-3776,32'd-4924,32'd-660,32'd162,32'd113,32'd-4697,32'd-93,32'd4724,32'd1431,32'd-3366,32'd5410,32'd-1788,32'd146,32'd-1962,32'd2790,32'd1211,32'd425,32'd763,32'd-4323,32'd-5864,32'd2202,32'd836,32'd1003,32'd-2749,32'd-2001,32'd-617,32'd2729,32'd-2008,32'd967,32'd106,32'd-4238,32'd2490,32'd1082,32'd-2440,32'd-255,32'd1619,32'd6552,32'd-531,32'd3701,32'd-3085,32'd3603,32'd-383,32'd690,32'd-210,32'd-375,32'd101,32'd1189,32'd-1872,32'd-841,32'd173,32'd883,32'd3903,32'd1993,32'd-2064,32'd-4128,32'd1412,32'd-2556,32'd-8081,32'd-139,32'd1584,32'd2098,32'd-463,32'd-67,32'd-4846,32'd1163,32'd2078,32'd-785,32'd-666,32'd693,32'd-2534,32'd3662,32'd-795,32'd-1739,32'd-2253,32'd295,32'd-1237,32'd-1370,32'd2086,32'd-7807,32'd1403,32'd5498,32'd-2724,32'd-459,32'd3635,32'd225,32'd-783,32'd1111,32'd-2371,32'd2065,32'd1921,32'd3061,32'd4880,32'd-2690,32'd1632,32'd1341,32'd-1178,32'd-794,32'd548,32'd4348,32'd-2095,32'd3244,32'd1274,32'd-3129,32'd-3994,32'd-3410,32'd-9316,32'd2181,32'd-1817,32'd-1633,32'd-558,32'd-1787,32'd-1483,32'd-1484,32'd4890,32'd3449,32'd-5478,32'd887,32'd-327,32'd-2912,32'd-3581,32'd-3295,32'd-3400,32'd-7348,32'd-3334,32'd-2070,32'd3898,32'd-1214,32'd-1702,32'd2261,32'd486,32'd272,32'd-177,32'd2463,32'd-2727,32'd-3937,32'd-3889,32'd981,32'd-2746,32'd-1875,32'd-220,32'd3684,32'd245,32'd729,32'd474,32'd2998,32'd-3867,32'd-2543,32'd2253,32'd133,32'd-4858,32'd-2183,32'd309,32'd-6557,32'd-806,32'd-6596,32'd7700,32'd-1211,32'd-3872,32'd1447,32'd-369,32'd-4096,32'd875,32'd-3027,32'd-1098,32'd-5405,32'd-1951,32'd-6777,32'd-410,32'd-4924,32'd-2244,32'd3723,32'd-1545,32'd-1503,32'd-1251,32'd-121,32'd139,32'd-4548,32'd786,32'd2700,32'd1636,32'd-5161,32'd2727,32'd2849,32'd947,32'd1111,32'd-2,32'd-1274,32'd4020,32'd2741,32'd6718,32'd-408,32'd952,32'd-2209,32'd860,32'd5126,32'd-1286,32'd3325};
    Wh[57]='{32'd1638,32'd5859,32'd466,32'd-5527,32'd590,32'd-2553,32'd-11728,32'd4699,32'd-2263,32'd-855,32'd2341,32'd337,32'd3852,32'd2551,32'd-4479,32'd1352,32'd-1647,32'd-2592,32'd-1580,32'd360,32'd-2058,32'd182,32'd1907,32'd-1768,32'd-121,32'd2413,32'd1865,32'd472,32'd-394,32'd-6796,32'd-4689,32'd-5659,32'd10,32'd2451,32'd-3254,32'd4191,32'd2355,32'd475,32'd-3378,32'd3789,32'd-508,32'd3459,32'd-4079,32'd5214,32'd3771,32'd-32,32'd-3117,32'd-2644,32'd-4697,32'd1225,32'd-6918,32'd2069,32'd529,32'd-945,32'd-2447,32'd-2939,32'd-712,32'd4570,32'd-1375,32'd2412,32'd-3183,32'd-7231,32'd314,32'd-1375,32'd7573,32'd-2358,32'd-2006,32'd1239,32'd-1042,32'd-1057,32'd-951,32'd126,32'd-2164,32'd-3022,32'd-246,32'd-1772,32'd-4357,32'd3610,32'd599,32'd537,32'd1560,32'd-5532,32'd5844,32'd-938,32'd141,32'd1286,32'd2937,32'd-1463,32'd-98,32'd-1350,32'd1833,32'd3786,32'd2233,32'd-484,32'd-1499,32'd1644,32'd153,32'd-164,32'd619,32'd1875,32'd-1501,32'd-707,32'd2121,32'd4057,32'd-2268,32'd2507,32'd-3132,32'd-14414,32'd-380,32'd-2403,32'd1560,32'd-596,32'd-3359,32'd-4147,32'd-5576,32'd-2253,32'd-7797,32'd-11718,32'd357,32'd-1878,32'd-3366,32'd-152,32'd1673,32'd-607,32'd4379,32'd2731,32'd-1680,32'd2702,32'd1390,32'd31406,32'd-3076,32'd309,32'd-3239,32'd2839,32'd-354,32'd2585,32'd-1488,32'd-236,32'd-3188,32'd5297,32'd-6093,32'd8359,32'd-7539,32'd-1557,32'd-849,32'd4306,32'd-1734,32'd-4306,32'd-172,32'd925,32'd-2966,32'd2644,32'd-1215,32'd-3676,32'd-739,32'd-5175,32'd-9375,32'd1907,32'd-5322,32'd7182,32'd-6801,32'd2117,32'd88,32'd-209,32'd-2932,32'd185,32'd2023,32'd-3034,32'd4323,32'd-3339,32'd4541,32'd1710,32'd1766,32'd-2053,32'd-1877,32'd-4284,32'd-4118,32'd-6796,32'd-11,32'd-155,32'd292,32'd7993,32'd-608,32'd442,32'd-2060,32'd-4853,32'd3806,32'd-5502,32'd2243,32'd-4445,32'd2795,32'd-1779,32'd989,32'd-1033,32'd-4475,32'd3593,32'd4560,32'd5727,32'd5263,32'd-947,32'd-491,32'd3725,32'd-298,32'd-696,32'd-625,32'd675,32'd-5693,32'd-8735,32'd-1622,32'd-178,32'd8007,32'd4187,32'd-242,32'd-1721,32'd4729,32'd-2325,32'd-3588,32'd-5507,32'd-1746,32'd1739,32'd-856,32'd-1403,32'd-644,32'd3723,32'd899,32'd3632,32'd397,32'd80,32'd511,32'd3049,32'd2534,32'd-5869,32'd1100,32'd775,32'd3530,32'd-4775,32'd2514,32'd593,32'd-3762,32'd-3828,32'd-1339,32'd-8408,32'd-2878,32'd1212,32'd-3273,32'd-661,32'd-2756,32'd3149,32'd-174,32'd-359,32'd-3679,32'd-3112,32'd-2687,32'd312,32'd4895,32'd-1710,32'd-4509,32'd-470,32'd-222,32'd4062,32'd5224,32'd1029,32'd3110,32'd648,32'd389,32'd-1823,32'd63,32'd1256,32'd-1480,32'd2651,32'd9443,32'd4108,32'd960,32'd-1580,32'd-1150,32'd8916,32'd4162,32'd-1296,32'd-1558,32'd103,32'd4587,32'd-619,32'd-2109,32'd-10595,32'd-1213,32'd-4819,32'd-1369,32'd1335,32'd-1837,32'd2900,32'd9814,32'd-14140,32'd-182,32'd-3962,32'd-7797,32'd6752,32'd-118,32'd-2276,32'd-1806,32'd-4567,32'd3823,32'd11542,32'd161,32'd-540,32'd642,32'd1139,32'd-3239,32'd-1866,32'd-5864,32'd1706,32'd-1287,32'd1091,32'd2990,32'd-6777,32'd-1646,32'd-805,32'd-7939,32'd-2658,32'd6308,32'd2178,32'd3623,32'd-3937,32'd-3991,32'd-34,32'd270,32'd-8,32'd-5058,32'd3132,32'd-1437,32'd-1071,32'd2248,32'd-3056,32'd1364,32'd87,32'd1752,32'd-6142,32'd1550,32'd8344,32'd5864,32'd-3161,32'd108,32'd836,32'd-2484,32'd-3574,32'd6533,32'd396,32'd-1510,32'd-5629,32'd4458,32'd-2856,32'd-2392,32'd-6108,32'd3125,32'd68,32'd7211,32'd-3259,32'd-4685,32'd16875,32'd9770,32'd3027,32'd-4772,32'd-3662,32'd-1776,32'd3178,32'd7387,32'd4440,32'd4501,32'd-603,32'd1290,32'd4882,32'd-736,32'd-4899,32'd334,32'd1174,32'd-3862,32'd-3334,32'd-7895,32'd-3410,32'd-3242,32'd-7758,32'd2626,32'd-2546,32'd-6591,32'd-4462,32'd3376,32'd3171,32'd3464,32'd7602,32'd-6337,32'd879,32'd10683,32'd-13359,32'd7626,32'd-5185,32'd-4519,32'd10410,32'd3913,32'd-2636,32'd-4392,32'd-140};
    Wh[58]='{32'd5073,32'd869,32'd-814,32'd2622,32'd548,32'd-1136,32'd4038,32'd-358,32'd-4135,32'd4047,32'd-1087,32'd2939,32'd-1368,32'd-298,32'd4274,32'd-85,32'd-241,32'd4890,32'd3530,32'd-1888,32'd-1322,32'd1915,32'd-605,32'd4731,32'd-371,32'd3801,32'd-1444,32'd170,32'd2761,32'd4375,32'd5424,32'd2242,32'd-1041,32'd4904,32'd4145,32'd3054,32'd2458,32'd2761,32'd-1100,32'd2145,32'd3005,32'd443,32'd3742,32'd-625,32'd638,32'd512,32'd5678,32'd1029,32'd-1613,32'd1342,32'd-1904,32'd-1522,32'd-2753,32'd-2185,32'd-8212,32'd-4934,32'd1436,32'd-8867,32'd3571,32'd2800,32'd-655,32'd1121,32'd-44,32'd-809,32'd-5263,32'd561,32'd-869,32'd2165,32'd4169,32'd-961,32'd-2058,32'd4448,32'd-409,32'd2106,32'd-309,32'd4135,32'd3342,32'd1475,32'd1846,32'd158,32'd1477,32'd6430,32'd-2399,32'd3378,32'd1678,32'd-1184,32'd-865,32'd-2437,32'd-2658,32'd2425,32'd4038,32'd-175,32'd2119,32'd-1436,32'd7397,32'd3725,32'd373,32'd111,32'd2307,32'd2851,32'd-5834,32'd-1840,32'd1378,32'd3171,32'd-4326,32'd1835,32'd5117,32'd5859,32'd1872,32'd983,32'd3920,32'd858,32'd-624,32'd2406,32'd2310,32'd-2805,32'd1518,32'd8754,32'd6015,32'd-5927,32'd-2751,32'd-8691,32'd-1556,32'd8051,32'd377,32'd2359,32'd2021,32'd223,32'd-3000,32'd-8041,32'd4020,32'd3405,32'd-2321,32'd-3188,32'd-6157,32'd4165,32'd5068,32'd-5966,32'd3635,32'd1450,32'd850,32'd-2819,32'd6494,32'd-2447,32'd-540,32'd-1365,32'd-2648,32'd2144,32'd4902,32'd1833,32'd-1888,32'd5097,32'd3708,32'd-5009,32'd2946,32'd-6015,32'd2880,32'd1220,32'd-2000,32'd-8803,32'd762,32'd4487,32'd-585,32'd-3554,32'd-2003,32'd-2792,32'd-671,32'd2573,32'd4704,32'd1696,32'd-2402,32'd-2509,32'd-3208,32'd3898,32'd-2961,32'd2442,32'd1916,32'd5014,32'd-5664,32'd2083,32'd2905,32'd128,32'd30,32'd2683,32'd-5063,32'd-3010,32'd696,32'd3847,32'd1250,32'd-1165,32'd-3229,32'd-2941,32'd661,32'd4592,32'd516,32'd5297,32'd-3117,32'd-2900,32'd506,32'd-3869,32'd-1429,32'd4990,32'd-4631,32'd1790,32'd4099,32'd607,32'd-1796,32'd5957,32'd472,32'd1701,32'd-3784,32'd2602,32'd9150,32'd-4294,32'd4467,32'd294,32'd-1075,32'd-415,32'd513,32'd1595,32'd4394,32'd6025,32'd2861,32'd-2462,32'd161,32'd1221,32'd3271,32'd1890,32'd1726,32'd-2683,32'd-394,32'd-1673,32'd8085,32'd-736,32'd5571,32'd-577,32'd-344,32'd-1679,32'd6723,32'd473,32'd2841,32'd-369,32'd3159,32'd-974,32'd-972,32'd392,32'd-1065,32'd-7026,32'd1788,32'd421,32'd3261,32'd952,32'd-1374,32'd-891,32'd-1932,32'd3354,32'd5283,32'd-1572,32'd4660,32'd-4001,32'd-2612,32'd7158,32'd5195,32'd3684,32'd-1773,32'd-462,32'd-153,32'd5761,32'd-364,32'd-2658,32'd-2141,32'd-5322,32'd1855,32'd-88,32'd-1574,32'd-7260,32'd2309,32'd6596,32'd-1052,32'd457,32'd-3876,32'd-609,32'd4570,32'd4287,32'd-2307,32'd-1540,32'd2442,32'd2519,32'd377,32'd-2019,32'd3500,32'd7866,32'd3825,32'd-1281,32'd1136,32'd3898,32'd1123,32'd-700,32'd5703,32'd-1832,32'd1468,32'd-6362,32'd-1557,32'd2873,32'd2081,32'd-651,32'd5761,32'd-705,32'd1309,32'd-700,32'd-2038,32'd1866,32'd3598,32'd8007,32'd4462,32'd2873,32'd3066,32'd-1822,32'd-1453,32'd6113,32'd3417,32'd5063,32'd1717,32'd-1540,32'd3852,32'd3139,32'd11650,32'd3681,32'd3950,32'd4821,32'd-994,32'd6704,32'd2756,32'd-1699,32'd-2578,32'd4489,32'd3090,32'd2961,32'd1667,32'd3774,32'd33,32'd773,32'd549,32'd2276,32'd3271,32'd-3457,32'd-5151,32'd2849,32'd14218,32'd4904,32'd-2883,32'd2253,32'd-2105,32'd-2541,32'd-1750,32'd586,32'd7553,32'd-1647,32'd60,32'd173,32'd8237,32'd7456,32'd5327,32'd1405,32'd-4626,32'd-3625,32'd-321,32'd2054,32'd513,32'd1219,32'd-1315,32'd2214,32'd-987,32'd6005,32'd391,32'd4858,32'd5522,32'd634,32'd-1934,32'd5097,32'd2651,32'd-1039,32'd-338,32'd2966,32'd-10,32'd4724,32'd3994,32'd-210,32'd663,32'd4333,32'd-1156,32'd3188,32'd-7670,32'd-435,32'd1795,32'd-7055,32'd-1502,32'd251,32'd4665,32'd1948};
    Wh[59]='{32'd-3686,32'd3286,32'd-1697,32'd-3012,32'd58,32'd-1000,32'd2261,32'd-1268,32'd2341,32'd-3596,32'd-5878,32'd-3425,32'd-2390,32'd5136,32'd-845,32'd-1210,32'd-9721,32'd157,32'd-221,32'd-784,32'd65,32'd1265,32'd1956,32'd1126,32'd-6704,32'd1113,32'd-2296,32'd445,32'd-906,32'd-2097,32'd2602,32'd-781,32'd-2792,32'd-4560,32'd-13935,32'd-4250,32'd-7080,32'd5209,32'd-1082,32'd479,32'd7612,32'd-2255,32'd1633,32'd-2619,32'd1579,32'd966,32'd8374,32'd-1351,32'd-3544,32'd718,32'd-2626,32'd-8320,32'd2021,32'd4133,32'd1718,32'd9267,32'd2502,32'd4704,32'd1745,32'd-10146,32'd5327,32'd-112,32'd3359,32'd-6904,32'd-6079,32'd123,32'd-520,32'd646,32'd-275,32'd-3977,32'd3354,32'd1291,32'd-3671,32'd1475,32'd247,32'd-825,32'd1257,32'd381,32'd5800,32'd-9687,32'd-1905,32'd3564,32'd24,32'd-579,32'd3808,32'd-4562,32'd263,32'd-543,32'd287,32'd-1203,32'd-2332,32'd-7426,32'd-366,32'd4875,32'd-572,32'd-2113,32'd-504,32'd-3510,32'd1342,32'd-1219,32'd1898,32'd444,32'd6914,32'd1146,32'd-1826,32'd-14,32'd4125,32'd2663,32'd5498,32'd-1264,32'd34,32'd-3605,32'd-2089,32'd1226,32'd307,32'd-10908,32'd-3527,32'd4777,32'd1839,32'd-12558,32'd2844,32'd905,32'd1685,32'd2065,32'd-11796,32'd-4174,32'd8881,32'd-1175,32'd3154,32'd-619,32'd1141,32'd-4431,32'd3151,32'd2751,32'd16904,32'd-1026,32'd-19208,32'd5336,32'd323,32'd-253,32'd-1311,32'd930,32'd6201,32'd-132,32'd1022,32'd-1218,32'd-1284,32'd-1813,32'd1799,32'd84,32'd-1770,32'd-48,32'd1596,32'd314,32'd-3859,32'd5048,32'd2834,32'd-1092,32'd4519,32'd-15722,32'd-5786,32'd-1850,32'd-4191,32'd-1900,32'd-5488,32'd8671,32'd1612,32'd370,32'd-6708,32'd-2435,32'd2839,32'd641,32'd191,32'd2817,32'd3701,32'd95,32'd468,32'd4401,32'd573,32'd-257,32'd-1937,32'd-7539,32'd1744,32'd1527,32'd-2426,32'd794,32'd2751,32'd-50,32'd193,32'd5205,32'd-4074,32'd-488,32'd-1651,32'd-1390,32'd834,32'd2988,32'd2170,32'd-3234,32'd-198,32'd-2125,32'd-4655,32'd4152,32'd-2344,32'd2485,32'd3642,32'd1408,32'd1848,32'd-877,32'd-2080,32'd-4401,32'd-5053,32'd1173,32'd-348,32'd515,32'd1516,32'd-5429,32'd-1326,32'd3562,32'd-3029,32'd-1468,32'd-1304,32'd-1590,32'd-2108,32'd7656,32'd4372,32'd-1668,32'd158,32'd138,32'd-2044,32'd-2783,32'd-2091,32'd-5019,32'd-1403,32'd-5229,32'd3610,32'd-1206,32'd-8388,32'd-1295,32'd3149,32'd2504,32'd-7924,32'd-1610,32'd-470,32'd4309,32'd-3710,32'd-396,32'd821,32'd-3083,32'd-3142,32'd-1904,32'd-6586,32'd-2539,32'd1589,32'd-2113,32'd-3601,32'd-7812,32'd3959,32'd3906,32'd-671,32'd1865,32'd-1671,32'd-5659,32'd2124,32'd-313,32'd-5541,32'd-5615,32'd-2280,32'd6650,32'd-2397,32'd-255,32'd-7026,32'd2360,32'd-3620,32'd-3405,32'd-8413,32'd-2490,32'd-3366,32'd-2218,32'd-4138,32'd-2236,32'd5346,32'd-7802,32'd-5771,32'd-670,32'd-718,32'd-915,32'd-451,32'd-1228,32'd-2479,32'd2724,32'd5820,32'd129,32'd-3662,32'd6079,32'd3537,32'd7827,32'd60,32'd-1330,32'd3076,32'd-371,32'd-1582,32'd-3059,32'd3771,32'd1840,32'd2237,32'd-6293,32'd-432,32'd-5917,32'd829,32'd813,32'd-3437,32'd-2646,32'd1334,32'd-721,32'd381,32'd-744,32'd-415,32'd1451,32'd-3061,32'd-3457,32'd5346,32'd-3693,32'd3808,32'd4187,32'd102,32'd2614,32'd1209,32'd-3132,32'd-37,32'd362,32'd3742,32'd-7636,32'd-8315,32'd-13681,32'd8457,32'd-4218,32'd7421,32'd7851,32'd-4294,32'd5712,32'd-1451,32'd346,32'd267,32'd314,32'd-2578,32'd-1340,32'd-7568,32'd5527,32'd7075,32'd-2014,32'd-1084,32'd-6772,32'd755,32'd-3425,32'd5922,32'd4243,32'd5722,32'd-2624,32'd-55,32'd-3286,32'd-651,32'd4794,32'd-6728,32'd-1434,32'd-5815,32'd-9394,32'd1578,32'd8857,32'd4482,32'd681,32'd-1743,32'd-938,32'd-1530,32'd-1545,32'd9018,32'd363,32'd3999,32'd-2111,32'd-611,32'd-2741,32'd2318,32'd-10449,32'd3681,32'd-5732,32'd2910,32'd2958,32'd1711,32'd2517,32'd6420,32'd-1783,32'd6347,32'd-7182,32'd758,32'd-1289,32'd30,32'd-2978,32'd2812,32'd-194,32'd3071,32'd-2880};
    Wh[60]='{32'd1503,32'd2810,32'd3540,32'd1229,32'd473,32'd-1613,32'd5205,32'd4501,32'd2318,32'd2604,32'd3964,32'd3535,32'd-3459,32'd534,32'd1879,32'd5097,32'd1049,32'd1234,32'd3281,32'd2266,32'd1500,32'd-4499,32'd-6958,32'd-185,32'd5551,32'd4797,32'd4733,32'd1027,32'd2678,32'd4428,32'd1839,32'd-761,32'd7661,32'd3271,32'd3820,32'd50,32'd3254,32'd-4194,32'd2326,32'd-711,32'd6264,32'd414,32'd2705,32'd-1782,32'd-4194,32'd1905,32'd749,32'd1312,32'd5561,32'd-9580,32'd-712,32'd4421,32'd-290,32'd4736,32'd6557,32'd-3652,32'd797,32'd3564,32'd6152,32'd-145,32'd17246,32'd2073,32'd3432,32'd3730,32'd10341,32'd3925,32'd1730,32'd144,32'd235,32'd1594,32'd4941,32'd-3605,32'd1457,32'd1602,32'd4458,32'd3850,32'd1687,32'd-5209,32'd-2932,32'd-5473,32'd1413,32'd2045,32'd341,32'd-2519,32'd7475,32'd-1357,32'd3994,32'd3452,32'd724,32'd8090,32'd3461,32'd6230,32'd4255,32'd668,32'd-880,32'd-2144,32'd2810,32'd-2609,32'd1442,32'd3708,32'd-3430,32'd1907,32'd-3623,32'd-2514,32'd-643,32'd-14,32'd-8007,32'd1614,32'd-9501,32'd3464,32'd3613,32'd2814,32'd5781,32'd-958,32'd1674,32'd2434,32'd-4965,32'd15214,32'd-4030,32'd-1361,32'd-258,32'd-2005,32'd10214,32'd34,32'd3762,32'd2053,32'd-4218,32'd-3618,32'd1372,32'd4167,32'd9291,32'd1654,32'd1539,32'd-617,32'd1667,32'd-2193,32'd-4853,32'd-1992,32'd-6162,32'd3801,32'd792,32'd-2398,32'd8115,32'd-3498,32'd-2371,32'd-4074,32'd-2049,32'd-9985,32'd-6250,32'd6455,32'd1501,32'd2556,32'd1259,32'd-2988,32'd5771,32'd4279,32'd-6235,32'd603,32'd-4445,32'd10410,32'd-3085,32'd3322,32'd2338,32'd-2482,32'd2812,32'd-1375,32'd15,32'd-4082,32'd-1882,32'd1685,32'd10546,32'd343,32'd5976,32'd-869,32'd-1130,32'd-6459,32'd-4287,32'd-8725,32'd-7133,32'd267,32'd-1878,32'd-2614,32'd-131,32'd3037,32'd1195,32'd2961,32'd-3393,32'd4406,32'd-1854,32'd1900,32'd5014,32'd2229,32'd-2924,32'd-27,32'd-283,32'd-1589,32'd-2402,32'd-1953,32'd-2563,32'd1901,32'd5859,32'd294,32'd1320,32'd2109,32'd2636,32'd151,32'd321,32'd1044,32'd7080,32'd171,32'd4968,32'd6459,32'd2359,32'd2037,32'd-995,32'd3740,32'd5239,32'd3923,32'd4011,32'd3989,32'd-107,32'd-4006,32'd3635,32'd4421,32'd3374,32'd6782,32'd1552,32'd-706,32'd6328,32'd4453,32'd6909,32'd7021,32'd-349,32'd6333,32'd7988,32'd3483,32'd274,32'd648,32'd-2006,32'd-1795,32'd2485,32'd-1420,32'd2399,32'd4294,32'd3659,32'd4504,32'd592,32'd4616,32'd-1021,32'd7597,32'd2303,32'd2800,32'd3784,32'd180,32'd9467,32'd-3569,32'd408,32'd-2005,32'd7124,32'd-2939,32'd5664,32'd9331,32'd8520,32'd-589,32'd-1828,32'd3305,32'd4113,32'd4135,32'd415,32'd3581,32'd6718,32'd1513,32'd1850,32'd2374,32'd3049,32'd942,32'd-1431,32'd3850,32'd7363,32'd4899,32'd1947,32'd-4360,32'd-1442,32'd444,32'd1862,32'd3945,32'd-132,32'd-3603,32'd-634,32'd-180,32'd853,32'd3488,32'd7626,32'd2397,32'd1348,32'd625,32'd859,32'd-3059,32'd-2253,32'd-5771,32'd764,32'd6064,32'd5830,32'd558,32'd2022,32'd1655,32'd1978,32'd2810,32'd4379,32'd4196,32'd2653,32'd6591,32'd4758,32'd2159,32'd6474,32'd4499,32'd1361,32'd3945,32'd3056,32'd-2775,32'd7412,32'd-734,32'd1839,32'd-1286,32'd1843,32'd2626,32'd1140,32'd-4108,32'd3322,32'd4062,32'd4572,32'd2316,32'd1898,32'd5585,32'd-7348,32'd-3261,32'd653,32'd-164,32'd8227,32'd1923,32'd2336,32'd2423,32'd5224,32'd-1676,32'd1492,32'd-3322,32'd2841,32'd5278,32'd733,32'd3500,32'd2614,32'd8896,32'd564,32'd960,32'd-1966,32'd-5444,32'd5097,32'd8603,32'd6596,32'd4916,32'd15361,32'd6943,32'd5629,32'd1297,32'd4470,32'd7504,32'd6513,32'd2951,32'd3032,32'd6689,32'd4741,32'd-3752,32'd941,32'd9326,32'd5141,32'd7280,32'd-336,32'd5141,32'd-7109,32'd-169,32'd8857,32'd-9248,32'd5419,32'd5107,32'd149,32'd2673,32'd4489,32'd5312,32'd-1776,32'd-1211,32'd2012,32'd4621,32'd8193,32'd-3208,32'd-5639,32'd192,32'd2126,32'd-13,32'd2058,32'd3894};
    Wh[61]='{32'd-5117,32'd-176,32'd4321,32'd-1307,32'd2056,32'd3681,32'd1080,32'd3618,32'd-699,32'd3095,32'd202,32'd-397,32'd-942,32'd1654,32'd-4248,32'd505,32'd-3051,32'd-900,32'd1015,32'd-3188,32'd2824,32'd1195,32'd-3117,32'd2556,32'd-9,32'd6870,32'd9414,32'd741,32'd6704,32'd5771,32'd2558,32'd-5014,32'd3920,32'd1524,32'd3110,32'd-2939,32'd-274,32'd-121,32'd1837,32'd1752,32'd88,32'd-3063,32'd1984,32'd2244,32'd-139,32'd-1022,32'd-915,32'd-3728,32'd3469,32'd-404,32'd-213,32'd5834,32'd-4824,32'd-1733,32'd-1977,32'd-2812,32'd153,32'd1795,32'd3249,32'd8994,32'd2376,32'd1398,32'd1209,32'd2279,32'd2199,32'd6264,32'd-3403,32'd-2758,32'd-527,32'd-4877,32'd5478,32'd4465,32'd-919,32'd5527,32'd-255,32'd102,32'd3125,32'd-1365,32'd-1728,32'd-4343,32'd714,32'd7768,32'd3107,32'd4543,32'd516,32'd1513,32'd-57,32'd-2125,32'd4370,32'd5869,32'd-2600,32'd-5317,32'd-690,32'd-1141,32'd-1170,32'd170,32'd-1505,32'd3281,32'd1805,32'd4074,32'd-2196,32'd-162,32'd-6127,32'd-1050,32'd4680,32'd-2156,32'd-3356,32'd2907,32'd-2646,32'd3217,32'd-680,32'd3715,32'd2010,32'd-1276,32'd3913,32'd-247,32'd2609,32'd1511,32'd-1401,32'd-3625,32'd521,32'd6708,32'd-1646,32'd5439,32'd4506,32'd-8925,32'd894,32'd-3615,32'd6420,32'd-653,32'd8383,32'd2858,32'd-5419,32'd4304,32'd673,32'd-4372,32'd-758,32'd1887,32'd3493,32'd4057,32'd5927,32'd2636,32'd-1658,32'd1760,32'd1233,32'd4851,32'd3498,32'd946,32'd8359,32'd-4143,32'd0,32'd-2446,32'd6518,32'd4689,32'd1889,32'd-1257,32'd-2978,32'd986,32'd1231,32'd-3557,32'd119,32'd-4870,32'd-3039,32'd4277,32'd2971,32'd-1676,32'd232,32'd772,32'd638,32'd-805,32'd4282,32'd-209,32'd-10947,32'd209,32'd6870,32'd-1215,32'd2431,32'd2258,32'd-3566,32'd4304,32'd1832,32'd-10888,32'd-1188,32'd-399,32'd-385,32'd-392,32'd2553,32'd-1226,32'd-1517,32'd242,32'd-1898,32'd40,32'd-1777,32'd-21,32'd-711,32'd2053,32'd90,32'd-4865,32'd1932,32'd-405,32'd2797,32'd3142,32'd689,32'd8164,32'd2343,32'd555,32'd2060,32'd1384,32'd4099,32'd-1721,32'd5161,32'd4523,32'd-2259,32'd2216,32'd6513,32'd3635,32'd2113,32'd-816,32'd4777,32'd-42,32'd-1014,32'd5385,32'd4091,32'd1374,32'd31,32'd6284,32'd-4011,32'd-360,32'd4086,32'd-157,32'd5590,32'd2934,32'd-4924,32'd1630,32'd3234,32'd5795,32'd2824,32'd936,32'd6953,32'd1706,32'd-2126,32'd2059,32'd180,32'd4392,32'd459,32'd34,32'd-1740,32'd-3193,32'd2888,32'd2089,32'd4785,32'd949,32'd2985,32'd1693,32'd-436,32'd2775,32'd574,32'd1547,32'd2832,32'd-2629,32'd1231,32'd977,32'd-1276,32'd2770,32'd-2939,32'd-2639,32'd2176,32'd2656,32'd709,32'd-1850,32'd2169,32'd-5454,32'd3500,32'd5517,32'd6210,32'd-2264,32'd3015,32'd-1162,32'd543,32'd-974,32'd651,32'd-3129,32'd2968,32'd4428,32'd4333,32'd1123,32'd480,32'd321,32'd-1071,32'd3435,32'd-2241,32'd11376,32'd-2071,32'd1728,32'd396,32'd2983,32'd-2233,32'd3039,32'd-1081,32'd-2602,32'd-1128,32'd-158,32'd2069,32'd2147,32'd-344,32'd5083,32'd-1397,32'd3574,32'd2998,32'd2187,32'd2648,32'd-52,32'd-2073,32'd1325,32'd-4116,32'd-861,32'd-434,32'd1435,32'd-2854,32'd-7626,32'd2622,32'd7441,32'd-3337,32'd-3488,32'd3972,32'd6376,32'd2653,32'd1119,32'd4748,32'd1986,32'd-1166,32'd-1545,32'd2362,32'd1237,32'd-4819,32'd4809,32'd-308,32'd-3664,32'd2316,32'd15,32'd-3417,32'd4799,32'd-193,32'd3903,32'd3146,32'd-1611,32'd3186,32'd-121,32'd14238,32'd586,32'd626,32'd8330,32'd-1853,32'd2653,32'd-3537,32'd-1439,32'd255,32'd7485,32'd8735,32'd255,32'd2529,32'd6210,32'd-279,32'd2878,32'd4667,32'd-1322,32'd2087,32'd-3725,32'd326,32'd-2519,32'd6728,32'd-1469,32'd-5385,32'd11894,32'd-895,32'd1644,32'd1370,32'd5727,32'd1795,32'd-4863,32'd3754,32'd5073,32'd-363,32'd-1007,32'd311,32'd4274,32'd746,32'd1787,32'd1030,32'd-1105,32'd1141,32'd-773,32'd4099,32'd-5200,32'd7031,32'd843,32'd-2944,32'd529,32'd-3635,32'd1369};
    Wh[62]='{32'd4331,32'd-600,32'd3085,32'd-458,32'd1258,32'd-980,32'd887,32'd1541,32'd4289,32'd-1032,32'd681,32'd845,32'd-650,32'd1166,32'd-2812,32'd-2666,32'd-897,32'd1160,32'd1070,32'd-2194,32'd-3645,32'd-1124,32'd1387,32'd-2208,32'd1121,32'd-3671,32'd57,32'd643,32'd324,32'd-1914,32'd-672,32'd2215,32'd-2998,32'd-3706,32'd2741,32'd5229,32'd834,32'd566,32'd-4829,32'd-1660,32'd-3869,32'd297,32'd1024,32'd1250,32'd82,32'd1199,32'd-1457,32'd9926,32'd-2583,32'd-1459,32'd2509,32'd-3674,32'd-4104,32'd-4958,32'd217,32'd-6142,32'd2937,32'd-422,32'd2983,32'd7846,32'd6582,32'd3835,32'd996,32'd3393,32'd4182,32'd1402,32'd637,32'd-1312,32'd-1212,32'd276,32'd6933,32'd-1020,32'd-100,32'd-2110,32'd553,32'd1933,32'd-2604,32'd2624,32'd-942,32'd484,32'd436,32'd-2255,32'd1767,32'd-870,32'd1707,32'd951,32'd-2946,32'd-2805,32'd4184,32'd-276,32'd-2449,32'd7075,32'd4736,32'd-808,32'd-2521,32'd5722,32'd456,32'd-1962,32'd1917,32'd749,32'd-709,32'd2697,32'd289,32'd-8325,32'd916,32'd753,32'd-4675,32'd1730,32'd897,32'd6132,32'd5620,32'd8618,32'd-3554,32'd-1750,32'd1242,32'd4672,32'd2386,32'd461,32'd-2434,32'd-6250,32'd-761,32'd-3442,32'd1320,32'd-2834,32'd1680,32'd911,32'd2294,32'd942,32'd53,32'd-3637,32'd-6884,32'd-763,32'd-1132,32'd-493,32'd1586,32'd1218,32'd-3266,32'd-3488,32'd-2500,32'd-173,32'd-3515,32'd3093,32'd3151,32'd-2534,32'd-2130,32'd-4389,32'd-870,32'd-7163,32'd2135,32'd-8374,32'd-2017,32'd726,32'd-5390,32'd1456,32'd-3791,32'd-3034,32'd-2424,32'd-1336,32'd-164,32'd14531,32'd-1138,32'd-4323,32'd-925,32'd2602,32'd3159,32'd2775,32'd3107,32'd2856,32'd484,32'd-393,32'd-1273,32'd3244,32'd943,32'd2269,32'd-116,32'd-3596,32'd2075,32'd-5473,32'd631,32'd4526,32'd625,32'd4135,32'd3425,32'd-1033,32'd-220,32'd512,32'd2113,32'd-7138,32'd6513,32'd-922,32'd757,32'd-5600,32'd-5712,32'd5024,32'd-616,32'd-3645,32'd-3945,32'd4912,32'd1045,32'd5268,32'd802,32'd2275,32'd206,32'd2229,32'd4362,32'd-232,32'd-3615,32'd5917,32'd-783,32'd3256,32'd1431,32'd3146,32'd-1810,32'd3332,32'd-400,32'd-2946,32'd-1353,32'd-2548,32'd1413,32'd699,32'd1194,32'd-1114,32'd-4575,32'd3498,32'd-1096,32'd6933,32'd2004,32'd2773,32'd1214,32'd-989,32'd5703,32'd-1111,32'd947,32'd-1950,32'd-284,32'd1229,32'd1495,32'd261,32'd-4096,32'd-2138,32'd-3103,32'd-112,32'd337,32'd-2094,32'd-1726,32'd-3703,32'd735,32'd-6137,32'd4443,32'd-629,32'd-2414,32'd101,32'd4162,32'd-231,32'd2077,32'd1746,32'd1341,32'd1304,32'd-322,32'd812,32'd-2641,32'd-408,32'd-1923,32'd-4233,32'd-825,32'd1351,32'd1284,32'd1137,32'd2421,32'd-1582,32'd631,32'd-2214,32'd4448,32'd315,32'd2592,32'd-3935,32'd-922,32'd-4118,32'd3381,32'd-578,32'd3720,32'd268,32'd-1065,32'd-5019,32'd-269,32'd-7714,32'd129,32'd3017,32'd-2145,32'd-4897,32'd-2807,32'd-28710,32'd-1674,32'd-7602,32'd5351,32'd374,32'd-6567,32'd756,32'd9238,32'd-7622,32'd2583,32'd1558,32'd886,32'd1124,32'd1475,32'd-1752,32'd5351,32'd-3298,32'd-470,32'd938,32'd4179,32'd3862,32'd-4111,32'd-1333,32'd-39,32'd-4062,32'd5937,32'd7749,32'd1268,32'd-109,32'd-491,32'd1097,32'd2344,32'd-5083,32'd-615,32'd-2890,32'd-1872,32'd645,32'd-1090,32'd1771,32'd6450,32'd-902,32'd-1005,32'd4904,32'd-1815,32'd-5332,32'd4172,32'd-154,32'd2749,32'd2504,32'd-3791,32'd970,32'd-1756,32'd-3669,32'd566,32'd4343,32'd2493,32'd1705,32'd-3291,32'd-2031,32'd3793,32'd3581,32'd1972,32'd1533,32'd760,32'd4047,32'd177,32'd-736,32'd867,32'd135,32'd5336,32'd4020,32'd-4528,32'd843,32'd181,32'd938,32'd-874,32'd2120,32'd-1024,32'd4428,32'd1326,32'd-7456,32'd-851,32'd-4111,32'd-7661,32'd-364,32'd5864,32'd2180,32'd-2322,32'd10283,32'd495,32'd-212,32'd-5087,32'd-1442,32'd-3708,32'd2365,32'd1905,32'd3557,32'd7216,32'd94,32'd4531,32'd-871,32'd7187,32'd5146,32'd8696,32'd3344,32'd-3173,32'd7700,32'd3955,32'd-814};
    Wh[63]='{32'd-4086,32'd4523,32'd-2303,32'd2131,32'd4084,32'd-577,32'd3283,32'd-2553,32'd1733,32'd-2121,32'd3740,32'd-3061,32'd1828,32'd-2988,32'd3164,32'd-5703,32'd4313,32'd-596,32'd384,32'd-18,32'd-2795,32'd2543,32'd-284,32'd4057,32'd6479,32'd8530,32'd2044,32'd2169,32'd-1798,32'd2010,32'd-2329,32'd-3208,32'd9931,32'd-389,32'd-255,32'd-377,32'd-1245,32'd1774,32'd4365,32'd2047,32'd-2534,32'd-792,32'd-7963,32'd297,32'd-209,32'd1856,32'd2197,32'd5922,32'd-702,32'd2169,32'd7543,32'd-393,32'd1488,32'd-5351,32'd-681,32'd3654,32'd4074,32'd-1494,32'd3242,32'd6962,32'd-7749,32'd1568,32'd1474,32'd12763,32'd8769,32'd-884,32'd1680,32'd2824,32'd-2037,32'd2156,32'd859,32'd2719,32'd-2069,32'd1896,32'd3005,32'd402,32'd211,32'd2369,32'd-1741,32'd-1846,32'd3151,32'd2150,32'd-795,32'd-957,32'd-1840,32'd2315,32'd-672,32'd2583,32'd7,32'd-2719,32'd171,32'd-808,32'd664,32'd-889,32'd1163,32'd1362,32'd-46,32'd3405,32'd-555,32'd-2678,32'd13496,32'd-1414,32'd2087,32'd2673,32'd-3503,32'd-828,32'd-4370,32'd213,32'd2739,32'd-4389,32'd-1627,32'd-4321,32'd6528,32'd193,32'd-657,32'd2142,32'd-725,32'd6367,32'd4975,32'd-4414,32'd-1806,32'd1008,32'd520,32'd1200,32'd5375,32'd4707,32'd-82,32'd-2344,32'd8623,32'd458,32'd3681,32'd-2045,32'd-2080,32'd5585,32'd-1755,32'd8168,32'd6586,32'd-63,32'd-1330,32'd-260,32'd-1052,32'd1385,32'd1217,32'd-7329,32'd747,32'd6591,32'd-4377,32'd-4133,32'd2736,32'd-470,32'd2438,32'd-3840,32'd1155,32'd8623,32'd-11269,32'd-5102,32'd3049,32'd2534,32'd-3217,32'd-4389,32'd-4121,32'd-1694,32'd25,32'd-685,32'd-6230,32'd-5224,32'd95,32'd5073,32'd173,32'd1810,32'd5034,32'd2507,32'd314,32'd1982,32'd-3508,32'd-4418,32'd232,32'd-2425,32'd1072,32'd-75,32'd-648,32'd-1920,32'd-2524,32'd-2470,32'd-6992,32'd1320,32'd-4528,32'd8090,32'd-16171,32'd-1367,32'd1580,32'd-803,32'd-5229,32'd4182,32'd-434,32'd2675,32'd3579,32'd-2109,32'd-1342,32'd4020,32'd-1214,32'd-4648,32'd2436,32'd595,32'd8583,32'd-855,32'd5839,32'd985,32'd3701,32'd1053,32'd-3017,32'd1270,32'd10019,32'd-895,32'd1839,32'd-772,32'd-1632,32'd761,32'd-579,32'd-5390,32'd-4672,32'd-2431,32'd-2390,32'd-3129,32'd-7387,32'd3852,32'd-3735,32'd-504,32'd6708,32'd396,32'd-2399,32'd3876,32'd-1988,32'd-406,32'd-2089,32'd2773,32'd-1859,32'd-3171,32'd-2250,32'd4243,32'd-313,32'd3891,32'd3483,32'd2091,32'd-425,32'd5214,32'd1154,32'd-1060,32'd1782,32'd-3662,32'd-1575,32'd-2312,32'd-1823,32'd-5966,32'd4082,32'd2352,32'd4145,32'd-5375,32'd2568,32'd1923,32'd-101,32'd-1160,32'd-1455,32'd447,32'd761,32'd625,32'd4313,32'd2091,32'd-1610,32'd227,32'd-5039,32'd1473,32'd4042,32'd-755,32'd1866,32'd-3520,32'd5439,32'd-1519,32'd-7324,32'd4545,32'd2912,32'd31,32'd-446,32'd-938,32'd2963,32'd-4079,32'd2000,32'd-5131,32'd-3293,32'd-1876,32'd5927,32'd6801,32'd-937,32'd1652,32'd2622,32'd2636,32'd2617,32'd138,32'd643,32'd-1428,32'd4755,32'd632,32'd3525,32'd-4812,32'd1148,32'd6904,32'd5351,32'd-3129,32'd3061,32'd-2880,32'd-2224,32'd-1235,32'd-2418,32'd2739,32'd3608,32'd-1523,32'd-1174,32'd-7041,32'd6962,32'd-3422,32'd4873,32'd-2229,32'd-3020,32'd558,32'd-2253,32'd1660,32'd495,32'd2247,32'd-539,32'd-4411,32'd-2888,32'd-2037,32'd1511,32'd827,32'd257,32'd3200,32'd-144,32'd-3303,32'd-2517,32'd-102,32'd-4838,32'd-1861,32'd-1466,32'd3164,32'd-6083,32'd-1453,32'd2045,32'd4997,32'd1248,32'd-5961,32'd2442,32'd2656,32'd-1741,32'd-3281,32'd-2128,32'd1667,32'd8510,32'd1075,32'd5283,32'd-6044,32'd-7861,32'd1102,32'd2476,32'd8750,32'd-5976,32'd5473,32'd3127,32'd-1956,32'd3693,32'd-324,32'd-1428,32'd-888,32'd2008,32'd2663,32'd-1871,32'd-722,32'd-4079,32'd-476,32'd-2851,32'd1151,32'd4694,32'd-3881,32'd8046,32'd-2736,32'd-957,32'd-754,32'd2644,32'd1082,32'd311,32'd-1343,32'd-2362,32'd1207,32'd3784,32'd-7622,32'd-1126,32'd-2178,32'd1322,32'd-2189,32'd930,32'd-4921};
    Wh[64]='{32'd-1295,32'd-3400,32'd3623,32'd-1960,32'd355,32'd277,32'd944,32'd7182,32'd-1093,32'd-3115,32'd-8554,32'd1396,32'd2082,32'd605,32'd-103,32'd-4284,32'd3852,32'd1585,32'd2316,32'd2418,32'd368,32'd-3986,32'd2622,32'd460,32'd-2539,32'd-6430,32'd1019,32'd-5000,32'd-3071,32'd3071,32'd4853,32'd-3164,32'd-9453,32'd-25,32'd114,32'd-441,32'd-3845,32'd76,32'd-11,32'd929,32'd-909,32'd-2053,32'd2873,32'd-588,32'd-2568,32'd-905,32'd2746,32'd837,32'd-2250,32'd2066,32'd1685,32'd-1163,32'd880,32'd2402,32'd582,32'd-1710,32'd-2059,32'd4113,32'd1057,32'd1572,32'd1202,32'd1322,32'd2404,32'd-2717,32'd-4528,32'd2139,32'd-5283,32'd1276,32'd4501,32'd-1479,32'd4965,32'd-892,32'd7182,32'd-955,32'd714,32'd-2751,32'd-2563,32'd-4692,32'd3095,32'd-1700,32'd2893,32'd7700,32'd-6083,32'd3554,32'd493,32'd2249,32'd-2336,32'd841,32'd5683,32'd2091,32'd1583,32'd687,32'd5122,32'd-3178,32'd-2493,32'd-4523,32'd562,32'd-574,32'd2646,32'd7514,32'd4655,32'd166,32'd-328,32'd-4094,32'd1206,32'd769,32'd1904,32'd7236,32'd-7949,32'd5649,32'd4567,32'd-410,32'd-10087,32'd-1828,32'd1809,32'd240,32'd903,32'd-4865,32'd-3559,32'd5927,32'd-2614,32'd-6127,32'd-4204,32'd-2861,32'd-12216,32'd-4316,32'd97,32'd3942,32'd254,32'd-1882,32'd212,32'd-4060,32'd285,32'd2602,32'd2602,32'd229,32'd-3593,32'd-1101,32'd-1458,32'd-889,32'd-8374,32'd5854,32'd-11181,32'd-702,32'd4729,32'd1172,32'd1616,32'd-767,32'd10595,32'd-1196,32'd-2022,32'd5185,32'd-4050,32'd-9550,32'd5317,32'd1855,32'd-3715,32'd3476,32'd-611,32'd-8178,32'd404,32'd-277,32'd2268,32'd-7656,32'd-5307,32'd12744,32'd7075,32'd-819,32'd-282,32'd-2410,32'd3767,32'd-2219,32'd606,32'd-3432,32'd473,32'd911,32'd-2259,32'd3093,32'd5952,32'd-3601,32'd693,32'd2861,32'd3869,32'd-4130,32'd4777,32'd942,32'd4851,32'd-4880,32'd3645,32'd1884,32'd-3544,32'd2885,32'd-9926,32'd2268,32'd-550,32'd-5380,32'd-1823,32'd3205,32'd1119,32'd1047,32'd-775,32'd2236,32'd4167,32'd-5722,32'd-1069,32'd1218,32'd124,32'd-5175,32'd-52,32'd-2541,32'd-2354,32'd-1021,32'd-11953,32'd-1492,32'd-622,32'd-4313,32'd-2254,32'd-6254,32'd3649,32'd1993,32'd426,32'd2331,32'd-1184,32'd104,32'd427,32'd-2431,32'd-5014,32'd-1810,32'd-6279,32'd497,32'd-2088,32'd-7373,32'd-12685,32'd-2308,32'd-1221,32'd-354,32'd3330,32'd-1025,32'd-3181,32'd-3178,32'd-1105,32'd-4528,32'd-979,32'd224,32'd-6093,32'd133,32'd789,32'd-1821,32'd1329,32'd3574,32'd-4472,32'd1993,32'd-5537,32'd-2232,32'd-383,32'd-7988,32'd-4128,32'd-5336,32'd-2727,32'd5424,32'd-672,32'd-3281,32'd2824,32'd6318,32'd1939,32'd-3371,32'd-4497,32'd4116,32'd1722,32'd-5751,32'd-2731,32'd-2279,32'd-1190,32'd-2827,32'd-6699,32'd3125,32'd-6293,32'd-4306,32'd-3007,32'd-3791,32'd-3339,32'd2612,32'd-5156,32'd1372,32'd-4291,32'd281,32'd-6655,32'd2636,32'd-1335,32'd-2670,32'd673,32'd-5693,32'd2927,32'd-554,32'd1788,32'd-2504,32'd-1988,32'd-99,32'd-355,32'd-6567,32'd732,32'd-9340,32'd3293,32'd-1567,32'd-1975,32'd3579,32'd8305,32'd-4455,32'd-5991,32'd616,32'd-3947,32'd-853,32'd-3647,32'd-6503,32'd7539,32'd-3991,32'd7504,32'd-2115,32'd6328,32'd-1695,32'd-4360,32'd733,32'd10478,32'd-3967,32'd6923,32'd700,32'd-586,32'd-4489,32'd5249,32'd8261,32'd437,32'd-200,32'd-2320,32'd-3913,32'd-639,32'd458,32'd-410,32'd6293,32'd4548,32'd-8750,32'd1719,32'd495,32'd2719,32'd-5932,32'd21,32'd-698,32'd5722,32'd-9355,32'd13427,32'd820,32'd2827,32'd-4128,32'd479,32'd-375,32'd4841,32'd-3183,32'd-3601,32'd-5776,32'd-1450,32'd2038,32'd5136,32'd2064,32'd-2412,32'd-5981,32'd-323,32'd-4582,32'd-2692,32'd-2392,32'd-2426,32'd6347,32'd4040,32'd-6030,32'd-706,32'd-2702,32'd594,32'd-6723,32'd-2531,32'd-6118,32'd-1682,32'd2205,32'd520,32'd-3583,32'd3876,32'd382,32'd-3010,32'd3869,32'd-3085,32'd1975,32'd3403,32'd5581,32'd2497,32'd-5932,32'd-1096,32'd9428,32'd-4570,32'd13476,32'd4265,32'd809,32'd-1232,32'd1148};
    Wh[65]='{32'd-583,32'd4846,32'd889,32'd-4108,32'd3791,32'd621,32'd-5937,32'd-2335,32'd-1368,32'd601,32'd-6064,32'd-4401,32'd-841,32'd2592,32'd958,32'd2349,32'd2266,32'd609,32'd-1605,32'd-2917,32'd1220,32'd-388,32'd-4770,32'd1680,32'd-2116,32'd-4592,32'd-2663,32'd3254,32'd-2651,32'd-496,32'd-1799,32'd-2866,32'd2268,32'd-1614,32'd-2797,32'd875,32'd522,32'd-1138,32'd-383,32'd-167,32'd-1936,32'd-1082,32'd7788,32'd1429,32'd-7768,32'd3662,32'd-6875,32'd-855,32'd-248,32'd631,32'd2751,32'd-1855,32'd-3110,32'd1879,32'd-4138,32'd2507,32'd1378,32'd1571,32'd-1033,32'd5268,32'd635,32'd-675,32'd-3442,32'd-1485,32'd5297,32'd-2458,32'd-1446,32'd1989,32'd1923,32'd-706,32'd-1636,32'd-4069,32'd-588,32'd145,32'd-1268,32'd-883,32'd-1076,32'd4680,32'd-1903,32'd-299,32'd-697,32'd326,32'd-5341,32'd1658,32'd-2795,32'd2281,32'd-1994,32'd-1953,32'd2827,32'd-1486,32'd-561,32'd1925,32'd1065,32'd-2451,32'd-975,32'd-1053,32'd-2961,32'd3205,32'd1192,32'd4296,32'd3664,32'd-3796,32'd2290,32'd-5483,32'd-325,32'd1074,32'd2683,32'd7485,32'd-13037,32'd3161,32'd3442,32'd-994,32'd3129,32'd-1530,32'd3271,32'd3422,32'd-1263,32'd-7353,32'd3708,32'd-2729,32'd-166,32'd-519,32'd-877,32'd-999,32'd1759,32'd-1921,32'd3747,32'd-640,32'd-880,32'd-6064,32'd2426,32'd-1342,32'd-2780,32'd-7504,32'd897,32'd-6777,32'd-6250,32'd-425,32'd-3811,32'd-1396,32'd2026,32'd-148,32'd1555,32'd2717,32'd-277,32'd-5087,32'd-2873,32'd-973,32'd-1468,32'd-3715,32'd-4943,32'd-3200,32'd-6806,32'd-4355,32'd-2780,32'd-7021,32'd-2006,32'd1464,32'd-2724,32'd5356,32'd3723,32'd1067,32'd1550,32'd4868,32'd-1770,32'd479,32'd3083,32'd110,32'd878,32'd-791,32'd10107,32'd8100,32'd-4355,32'd-818,32'd-7426,32'd-5839,32'd3061,32'd-409,32'd1988,32'd303,32'd925,32'd-6611,32'd6855,32'd-726,32'd-1206,32'd3786,32'd-1701,32'd-97,32'd-5288,32'd-196,32'd895,32'd-1429,32'd952,32'd-1722,32'd1687,32'd-4011,32'd-2917,32'd-2507,32'd-1699,32'd-5180,32'd-33,32'd5087,32'd-717,32'd-2095,32'd304,32'd-968,32'd-1641,32'd2426,32'd6987,32'd-2163,32'd4165,32'd1135,32'd2269,32'd-1005,32'd-1500,32'd-3410,32'd-2856,32'd-3310,32'd-466,32'd-484,32'd466,32'd3300,32'd3212,32'd6059,32'd319,32'd-1612,32'd821,32'd-858,32'd364,32'd2958,32'd-3586,32'd-3349,32'd1021,32'd408,32'd1644,32'd1061,32'd-199,32'd894,32'd-5107,32'd-3181,32'd659,32'd-3559,32'd4516,32'd-5053,32'd3784,32'd-198,32'd957,32'd1495,32'd1575,32'd4084,32'd2746,32'd-2496,32'd-4028,32'd-470,32'd-4675,32'd5244,32'd2479,32'd-1622,32'd-467,32'd-9677,32'd-4152,32'd3032,32'd6611,32'd519,32'd1130,32'd-894,32'd-628,32'd-7333,32'd3029,32'd-308,32'd1182,32'd-589,32'd2519,32'd818,32'd-1165,32'd-4609,32'd594,32'd809,32'd1805,32'd1074,32'd1155,32'd-5703,32'd1467,32'd-8627,32'd-633,32'd2817,32'd-2707,32'd-85,32'd7,32'd3530,32'd3374,32'd-1104,32'd1286,32'd-4697,32'd-3942,32'd-3208,32'd-256,32'd-1368,32'd5751,32'd-2006,32'd-1883,32'd-1259,32'd-2437,32'd-1391,32'd1347,32'd176,32'd-2371,32'd-1085,32'd2387,32'd925,32'd-1983,32'd-1724,32'd125,32'd-4794,32'd-6503,32'd1437,32'd120,32'd-2626,32'd572,32'd1901,32'd-2788,32'd2641,32'd1256,32'd5273,32'd-330,32'd-5917,32'd-2302,32'd-1170,32'd-138,32'd-3017,32'd-23,32'd-70,32'd-9033,32'd4006,32'd-3952,32'd6831,32'd-860,32'd340,32'd-2127,32'd-4299,32'd-5327,32'd17,32'd2761,32'd-3464,32'd-7392,32'd7758,32'd946,32'd-1082,32'd-787,32'd-1109,32'd2225,32'd-3381,32'd-2937,32'd-180,32'd-1733,32'd10029,32'd4670,32'd3259,32'd-508,32'd-3520,32'd-696,32'd-460,32'd159,32'd1824,32'd-1021,32'd-361,32'd-131,32'd99,32'd2315,32'd-364,32'd4587,32'd-326,32'd4184,32'd-4343,32'd-1181,32'd-3090,32'd-438,32'd1436,32'd-5532,32'd3703,32'd-31,32'd-4792,32'd455,32'd-4963,32'd-2222,32'd2907,32'd-1115,32'd-4931,32'd-2700,32'd1077,32'd991,32'd-5185,32'd148,32'd-6503,32'd-5351,32'd2060,32'd-2790,32'd-1427,32'd2607,32'd1395};
    Wh[66]='{32'd-1252,32'd6699,32'd4204,32'd-485,32'd1043,32'd-1062,32'd-5727,32'd-4377,32'd-2678,32'd2293,32'd2644,32'd-531,32'd-1889,32'd3344,32'd5126,32'd-8520,32'd5932,32'd2153,32'd2893,32'd-1263,32'd-647,32'd850,32'd-597,32'd1217,32'd-1994,32'd2607,32'd525,32'd-1529,32'd-1901,32'd-458,32'd2145,32'd1561,32'd1188,32'd-108,32'd-1901,32'd-1002,32'd-4538,32'd2451,32'd-2335,32'd6879,32'd-1901,32'd2197,32'd-1993,32'd2288,32'd-863,32'd-1776,32'd-5014,32'd-1574,32'd1105,32'd-1008,32'd-8681,32'd266,32'd-703,32'd1102,32'd636,32'd-3759,32'd2470,32'd-101,32'd-1295,32'd1779,32'd-913,32'd-2347,32'd2033,32'd-68,32'd-1227,32'd-411,32'd-5625,32'd6391,32'd-419,32'd-19,32'd-2692,32'd-840,32'd1987,32'd-78,32'd3120,32'd527,32'd-14,32'd3435,32'd774,32'd-3164,32'd1719,32'd2910,32'd-3559,32'd3032,32'd-1073,32'd-1121,32'd209,32'd1022,32'd-5844,32'd-1328,32'd2814,32'd2849,32'd-1408,32'd3854,32'd-1806,32'd-3500,32'd605,32'd-2192,32'd3212,32'd-2493,32'd-2785,32'd2910,32'd373,32'd6318,32'd-4804,32'd3862,32'd1900,32'd1724,32'd-1001,32'd732,32'd2072,32'd431,32'd-1995,32'd-1602,32'd5092,32'd519,32'd-4121,32'd-3071,32'd-1840,32'd-3041,32'd-2548,32'd2032,32'd-188,32'd4536,32'd-919,32'd4746,32'd-278,32'd-3537,32'd-5039,32'd-6054,32'd811,32'd-2498,32'd1303,32'd-1440,32'd-3872,32'd-628,32'd-6215,32'd3269,32'd-4543,32'd-2398,32'd-3835,32'd2331,32'd-5253,32'd3901,32'd2790,32'd-7031,32'd437,32'd-4875,32'd1591,32'd-1082,32'd-8823,32'd-20,32'd-3347,32'd4345,32'd-1430,32'd-2500,32'd-3581,32'd504,32'd-376,32'd6738,32'd-2426,32'd-3959,32'd-1953,32'd-892,32'd5888,32'd-1431,32'd2481,32'd2178,32'd-121,32'd-1149,32'd130,32'd10009,32'd687,32'd-403,32'd3073,32'd637,32'd764,32'd-258,32'd1284,32'd2281,32'd-3789,32'd-1986,32'd7207,32'd3752,32'd-5107,32'd1708,32'd-518,32'd238,32'd8300,32'd-3986,32'd-1732,32'd-89,32'd5371,32'd-1054,32'd466,32'd767,32'd474,32'd1250,32'd-185,32'd-392,32'd-52,32'd2541,32'd-1034,32'd3913,32'd2167,32'd294,32'd-15,32'd2048,32'd-1654,32'd544,32'd646,32'd897,32'd1513,32'd3762,32'd-2648,32'd828,32'd-870,32'd-4331,32'd89,32'd-4758,32'd-1353,32'd3085,32'd1892,32'd5756,32'd-3212,32'd-5712,32'd3637,32'd543,32'd-8535,32'd3405,32'd4589,32'd3999,32'd5664,32'd396,32'd9228,32'd1008,32'd-459,32'd2182,32'd1143,32'd-5361,32'd-1002,32'd-7099,32'd3684,32'd2841,32'd-3249,32'd-14,32'd1668,32'd-4592,32'd-1842,32'd3413,32'd997,32'd-1462,32'd-1981,32'd-4042,32'd1324,32'd1821,32'd-1392,32'd2551,32'd-5629,32'd-410,32'd1411,32'd1407,32'd4375,32'd4624,32'd4501,32'd-1733,32'd1702,32'd-747,32'd-1280,32'd-795,32'd-2004,32'd-2423,32'd1386,32'd2467,32'd-842,32'd-3708,32'd236,32'd1112,32'd1020,32'd816,32'd3422,32'd4533,32'd-720,32'd-6342,32'd394,32'd2810,32'd-784,32'd4809,32'd2578,32'd-358,32'd-1155,32'd-1813,32'd1169,32'd1174,32'd-3955,32'd7924,32'd-23,32'd281,32'd4233,32'd-5771,32'd-15,32'd-26,32'd2424,32'd3200,32'd-206,32'd866,32'd3522,32'd-4672,32'd838,32'd6831,32'd1771,32'd6723,32'd-1954,32'd-575,32'd-1457,32'd-4011,32'd-1461,32'd1989,32'd3388,32'd-1466,32'd-4250,32'd4384,32'd2644,32'd3884,32'd-4409,32'd-1972,32'd6367,32'd-764,32'd-6499,32'd-3471,32'd2380,32'd-2773,32'd3286,32'd3156,32'd2076,32'd1345,32'd-1374,32'd3645,32'd3991,32'd-942,32'd-5273,32'd357,32'd-975,32'd-702,32'd-6562,32'd4279,32'd-9125,32'd-3229,32'd7543,32'd-1873,32'd-3649,32'd1279,32'd-1047,32'd-3547,32'd6162,32'd3344,32'd-960,32'd7026,32'd-3322,32'd1920,32'd-1150,32'd3276,32'd-2507,32'd-1981,32'd-3144,32'd2844,32'd661,32'd-721,32'd-2937,32'd8793,32'd697,32'd5942,32'd1536,32'd-1606,32'd3464,32'd2420,32'd-963,32'd2001,32'd341,32'd251,32'd4145,32'd-2985,32'd-2861,32'd-38,32'd3383,32'd1741,32'd-132,32'd4729,32'd-4819,32'd529,32'd-1538,32'd-2949,32'd2292,32'd-1389,32'd-249,32'd1669,32'd-5141,32'd-3530,32'd-1078,32'd-1827};
    Wh[67]='{32'd4428,32'd10537,32'd-676,32'd-3161,32'd615,32'd24,32'd-3142,32'd2768,32'd6157,32'd929,32'd4082,32'd8120,32'd5058,32'd-2617,32'd5678,32'd9907,32'd3688,32'd15000,32'd7319,32'd-336,32'd4052,32'd-207,32'd-3037,32'd828,32'd1419,32'd8461,32'd1916,32'd3125,32'd-1525,32'd1733,32'd-1307,32'd-8232,32'd1806,32'd833,32'd-1999,32'd743,32'd1802,32'd5,32'd-3498,32'd78,32'd3510,32'd5190,32'd10800,32'd2556,32'd4077,32'd3410,32'd-769,32'd2413,32'd-637,32'd3920,32'd-171,32'd-4235,32'd5068,32'd-387,32'd10869,32'd4479,32'd-2055,32'd2578,32'd-5971,32'd10507,32'd-3557,32'd3261,32'd-1177,32'd2189,32'd6254,32'd-971,32'd-1035,32'd-4462,32'd-2021,32'd-592,32'd-1226,32'd3488,32'd3332,32'd451,32'd3354,32'd-2551,32'd-770,32'd7553,32'd5522,32'd1362,32'd-1827,32'd4365,32'd1503,32'd4472,32'd-3872,32'd-6899,32'd-711,32'd-2792,32'd5869,32'd3249,32'd7797,32'd-4226,32'd4060,32'd-3188,32'd-6557,32'd48,32'd379,32'd2219,32'd2597,32'd-913,32'd522,32'd4797,32'd-1730,32'd11035,32'd-2330,32'd-2202,32'd-1007,32'd5332,32'd-3708,32'd-1950,32'd-566,32'd-19677,32'd2237,32'd1721,32'd-920,32'd-5854,32'd6376,32'd-2512,32'd-2222,32'd4116,32'd-1013,32'd-2136,32'd8901,32'd6103,32'd1802,32'd2152,32'd5141,32'd5234,32'd-6499,32'd6972,32'd-3542,32'd2624,32'd276,32'd7011,32'd10273,32'd9306,32'd9296,32'd1030,32'd-3212,32'd2546,32'd-3317,32'd-1468,32'd-3251,32'd-995,32'd910,32'd-3637,32'd2303,32'd-4189,32'd1168,32'd767,32'd1345,32'd1302,32'd3112,32'd-2619,32'd-865,32'd-3342,32'd5136,32'd-4130,32'd-232,32'd17910,32'd7880,32'd-1108,32'd548,32'd-3610,32'd3120,32'd249,32'd1434,32'd108,32'd1110,32'd-113,32'd2492,32'd-224,32'd2094,32'd2685,32'd-393,32'd-1448,32'd-920,32'd-1437,32'd-445,32'd4812,32'd3520,32'd8837,32'd-5439,32'd-1040,32'd-3461,32'd-2130,32'd7045,32'd-6508,32'd-13935,32'd-2219,32'd-131,32'd-3212,32'd-3085,32'd8818,32'd3793,32'd10722,32'd1413,32'd2255,32'd4804,32'd1205,32'd-1953,32'd2100,32'd-3547,32'd-8745,32'd2973,32'd-1445,32'd-623,32'd-5039,32'd2376,32'd3696,32'd-165,32'd-867,32'd6030,32'd-8769,32'd2597,32'd-5078,32'd-3420,32'd1646,32'd-2218,32'd-3769,32'd2290,32'd1364,32'd-3400,32'd-357,32'd-4306,32'd4931,32'd-2167,32'd-1376,32'd2609,32'd1342,32'd2401,32'd2362,32'd-733,32'd-1730,32'd-6679,32'd-2379,32'd-6748,32'd5463,32'd-5502,32'd3193,32'd-1445,32'd946,32'd-6245,32'd7578,32'd-4003,32'd-647,32'd-7138,32'd-3168,32'd-255,32'd-3635,32'd-5590,32'd-2846,32'd-237,32'd-1267,32'd1003,32'd-2687,32'd-1966,32'd-2373,32'd-798,32'd-8500,32'd-2181,32'd-5673,32'd9423,32'd-1081,32'd-6713,32'd-6865,32'd-3422,32'd6909,32'd1333,32'd-3588,32'd-2626,32'd2768,32'd-986,32'd1194,32'd-2465,32'd1608,32'd3349,32'd-3522,32'd-356,32'd-4357,32'd4416,32'd-3322,32'd-1630,32'd3078,32'd-3564,32'd2180,32'd1195,32'd-4265,32'd-2705,32'd372,32'd-9863,32'd3864,32'd4990,32'd-969,32'd-2658,32'd1898,32'd-4353,32'd-5161,32'd7041,32'd-202,32'd-310,32'd2445,32'd-4460,32'd-1774,32'd1868,32'd2366,32'd1258,32'd265,32'd2976,32'd3684,32'd-2558,32'd7382,32'd-5312,32'd-603,32'd2836,32'd4741,32'd-6381,32'd-1303,32'd-2030,32'd-4836,32'd4064,32'd-6459,32'd1002,32'd-5117,32'd-4160,32'd-431,32'd3808,32'd-3181,32'd531,32'd-2661,32'd2325,32'd-6977,32'd691,32'd-5092,32'd5463,32'd5283,32'd2680,32'd1157,32'd-339,32'd-4140,32'd-5502,32'd-1589,32'd-684,32'd3896,32'd1258,32'd-1501,32'd5727,32'd2875,32'd7739,32'd509,32'd-7387,32'd-4113,32'd2607,32'd-5834,32'd-2191,32'd868,32'd6630,32'd-3884,32'd3923,32'd-2293,32'd2922,32'd3635,32'd350,32'd-824,32'd3095,32'd2551,32'd-5151,32'd-189,32'd-5234,32'd-13574,32'd-3266,32'd3972,32'd-2541,32'd-2139,32'd-7749,32'd-3403,32'd-1569,32'd6147,32'd4604,32'd2988,32'd7514,32'd4089,32'd-2758,32'd1140,32'd6093,32'd-6098,32'd-2203,32'd1331,32'd9414,32'd-3093,32'd-2352,32'd-7050,32'd3203,32'd-2770,32'd270,32'd-2763,32'd-2963,32'd8339,32'd323,32'd-2187};
    Wh[68]='{32'd-2016,32'd5141,32'd1257,32'd-3120,32'd3161,32'd-93,32'd2282,32'd-5239,32'd-661,32'd5180,32'd4987,32'd178,32'd-6069,32'd3066,32'd5517,32'd4780,32'd7778,32'd2592,32'd640,32'd-1115,32'd-957,32'd1291,32'd1105,32'd691,32'd2609,32'd-6362,32'd-2673,32'd1032,32'd-4345,32'd4287,32'd-40,32'd1673,32'd2727,32'd974,32'd-5097,32'd-2072,32'd-2531,32'd606,32'd1099,32'd852,32'd237,32'd5253,32'd-7900,32'd5307,32'd-3024,32'd-1697,32'd242,32'd2902,32'd-1469,32'd-1146,32'd-7299,32'd1386,32'd-124,32'd10185,32'd-5766,32'd-407,32'd-161,32'd-457,32'd689,32'd2253,32'd-2438,32'd886,32'd3364,32'd2692,32'd2563,32'd-2038,32'd-159,32'd1655,32'd-1127,32'd-1273,32'd-5810,32'd3127,32'd-1525,32'd6831,32'd6582,32'd-4599,32'd3251,32'd-3476,32'd-444,32'd-25,32'd-112,32'd1738,32'd-3496,32'd6816,32'd1701,32'd245,32'd106,32'd325,32'd-1491,32'd-3906,32'd258,32'd5053,32'd-154,32'd-2476,32'd2036,32'd-3105,32'd-1340,32'd5092,32'd2261,32'd5673,32'd5678,32'd-3132,32'd-2448,32'd-4406,32'd-1508,32'd3393,32'd4089,32'd3547,32'd-896,32'd607,32'd5864,32'd2656,32'd592,32'd1920,32'd4599,32'd-2639,32'd-2239,32'd-4169,32'd4580,32'd-1145,32'd-2629,32'd-4016,32'd1276,32'd3469,32'd4416,32'd985,32'd3188,32'd-653,32'd-3017,32'd-8618,32'd-2384,32'd3684,32'd1237,32'd880,32'd-6757,32'd1630,32'd358,32'd-3566,32'd-1910,32'd-2418,32'd-2314,32'd722,32'd2038,32'd-4440,32'd-1663,32'd1135,32'd-635,32'd2293,32'd-2066,32'd-5454,32'd-3569,32'd123,32'd-10673,32'd1785,32'd-684,32'd-1850,32'd-7792,32'd4233,32'd3676,32'd8569,32'd-2126,32'd-4291,32'd6889,32'd1122,32'd2020,32'd311,32'd-630,32'd5253,32'd2917,32'd-116,32'd5151,32'd6240,32'd-6547,32'd3815,32'd-67,32'd1708,32'd4360,32'd-6479,32'd8105,32'd-2653,32'd-4870,32'd-13662,32'd-1162,32'd-3015,32'd-739,32'd3457,32'd-728,32'd561,32'd-1188,32'd-3273,32'd3422,32'd3205,32'd2443,32'd-4074,32'd-2364,32'd6059,32'd-2293,32'd1949,32'd-3232,32'd2486,32'd3479,32'd-3547,32'd-1145,32'd-243,32'd382,32'd-1530,32'd681,32'd-2683,32'd983,32'd6411,32'd-4873,32'd7250,32'd3044,32'd-445,32'd1484,32'd-83,32'd-847,32'd995,32'd2609,32'd-3811,32'd2329,32'd2868,32'd-2187,32'd6845,32'd2653,32'd5893,32'd4562,32'd184,32'd3188,32'd-18,32'd7177,32'd-7680,32'd-3666,32'd-909,32'd2316,32'd3415,32'd2788,32'd-466,32'd2084,32'd238,32'd-1107,32'd-7856,32'd2568,32'd920,32'd1661,32'd-3225,32'd4460,32'd2401,32'd-3068,32'd5781,32'd-1,32'd-1822,32'd-2619,32'd3037,32'd809,32'd-1348,32'd5229,32'd-91,32'd-215,32'd-2425,32'd9506,32'd1666,32'd314,32'd527,32'd-926,32'd-4392,32'd705,32'd4929,32'd1408,32'd1473,32'd6484,32'd121,32'd5600,32'd1939,32'd4958,32'd1040,32'd2467,32'd5727,32'd-2644,32'd2156,32'd6767,32'd-3127,32'd-1628,32'd-283,32'd-1859,32'd-1286,32'd2067,32'd1427,32'd7539,32'd1041,32'd4616,32'd7558,32'd978,32'd-7373,32'd-1217,32'd-4113,32'd4160,32'd-16,32'd3164,32'd-1182,32'd-737,32'd3732,32'd3688,32'd-972,32'd-23,32'd5737,32'd2985,32'd811,32'd-1007,32'd5039,32'd-4592,32'd4711,32'd-1425,32'd4055,32'd3432,32'd1713,32'd-188,32'd-1113,32'd2788,32'd-2443,32'd8203,32'd6855,32'd26,32'd3596,32'd2360,32'd1722,32'd6318,32'd-1862,32'd-1593,32'd-6782,32'd8540,32'd5844,32'd3862,32'd4721,32'd-3205,32'd6342,32'd-1365,32'd900,32'd108,32'd-4558,32'd-3730,32'd-4855,32'd-37,32'd-1712,32'd-8710,32'd-233,32'd-2629,32'd-220,32'd6166,32'd405,32'd-4699,32'd-3964,32'd1306,32'd4538,32'd-1322,32'd-7314,32'd5751,32'd13134,32'd7270,32'd-204,32'd-1658,32'd2700,32'd3703,32'd-1143,32'd-9775,32'd1762,32'd5927,32'd-3559,32'd-3098,32'd5068,32'd1586,32'd-5224,32'd6367,32'd4377,32'd4726,32'd-1284,32'd3271,32'd-495,32'd2211,32'd-2272,32'd2702,32'd-1029,32'd301,32'd-578,32'd-1685,32'd-1231,32'd1044,32'd-3913,32'd-610,32'd-1661,32'd-3642,32'd5468,32'd4899,32'd-7358,32'd7670,32'd-1286,32'd-1684,32'd1643,32'd4306,32'd-782};
    Wh[69]='{32'd105,32'd-4511,32'd-866,32'd-2175,32'd-1981,32'd3417,32'd-1649,32'd-1097,32'd3552,32'd-4438,32'd-2354,32'd-723,32'd743,32'd-1661,32'd1154,32'd698,32'd-3835,32'd1334,32'd355,32'd-1282,32'd2868,32'd-1752,32'd-2352,32'd1120,32'd-365,32'd-891,32'd-3354,32'd2810,32'd6132,32'd2968,32'd-493,32'd1625,32'd-5000,32'd26,32'd2102,32'd1134,32'd-3759,32'd-1984,32'd-196,32'd-4394,32'd481,32'd-3649,32'd8925,32'd-3332,32'd2469,32'd-1166,32'd2770,32'd4291,32'd-102,32'd1210,32'd5219,32'd-1485,32'd-3271,32'd-4023,32'd3945,32'd-5800,32'd-2902,32'd-2324,32'd406,32'd3,32'd3439,32'd36,32'd-1036,32'd4091,32'd1976,32'd3007,32'd1658,32'd8471,32'd-2030,32'd1265,32'd1613,32'd85,32'd-2458,32'd437,32'd-2519,32'd631,32'd1646,32'd-1883,32'd-4448,32'd2053,32'd-4096,32'd3447,32'd1602,32'd-7226,32'd3073,32'd-2442,32'd102,32'd1267,32'd-1920,32'd2058,32'd-1975,32'd2172,32'd-2482,32'd-2602,32'd3317,32'd2612,32'd0,32'd-2868,32'd-5600,32'd2990,32'd-4291,32'd258,32'd-296,32'd-7358,32'd4611,32'd-1678,32'd-5976,32'd-2036,32'd-4045,32'd-5981,32'd-519,32'd413,32'd5029,32'd733,32'd-4116,32'd-4338,32'd5419,32'd8725,32'd-308,32'd7558,32'd1722,32'd-3862,32'd-1953,32'd-4643,32'd-1645,32'd3461,32'd-5522,32'd1297,32'd10039,32'd1890,32'd-3095,32'd4235,32'd2990,32'd3461,32'd-4096,32'd3464,32'd5766,32'd992,32'd1380,32'd78,32'd-1849,32'd2907,32'd-4270,32'd-1303,32'd-2058,32'd-4130,32'd8774,32'd-965,32'd6547,32'd-1921,32'd6435,32'd-5063,32'd2012,32'd-3630,32'd3918,32'd1722,32'd1807,32'd-5278,32'd-7329,32'd1068,32'd5410,32'd6870,32'd239,32'd2122,32'd-4565,32'd-875,32'd-2023,32'd2274,32'd-3317,32'd1622,32'd-968,32'd-8569,32'd-4748,32'd-2949,32'd898,32'd-1564,32'd1702,32'd7158,32'd-3173,32'd752,32'd558,32'd12480,32'd-7011,32'd5849,32'd7124,32'd-2763,32'd-3854,32'd2883,32'd-4204,32'd7080,32'd-1791,32'd3195,32'd-6796,32'd2199,32'd1334,32'd1527,32'd3479,32'd-4042,32'd-3608,32'd-937,32'd2491,32'd4714,32'd411,32'd44,32'd-3041,32'd-141,32'd-501,32'd-3342,32'd-1239,32'd-1052,32'd-772,32'd-2714,32'd3110,32'd-1212,32'd3684,32'd758,32'd-502,32'd-1519,32'd-2775,32'd5068,32'd2097,32'd-778,32'd712,32'd-286,32'd-9755,32'd-1909,32'd-177,32'd600,32'd-1341,32'd-1209,32'd2409,32'd3593,32'd8198,32'd-991,32'd-11093,32'd-1791,32'd-1571,32'd-610,32'd-854,32'd-1445,32'd79,32'd823,32'd3881,32'd1234,32'd-983,32'd-274,32'd-155,32'd282,32'd374,32'd-4758,32'd3828,32'd5737,32'd-1806,32'd-455,32'd1287,32'd1055,32'd-3557,32'd-3784,32'd742,32'd-5478,32'd-2219,32'd2626,32'd303,32'd-1817,32'd1186,32'd3989,32'd-686,32'd-3305,32'd505,32'd286,32'd-2509,32'd-5854,32'd-415,32'd-23,32'd1895,32'd-1520,32'd-4184,32'd3937,32'd-858,32'd-3073,32'd-5185,32'd-757,32'd-568,32'd2252,32'd2255,32'd-8466,32'd2414,32'd-5097,32'd213,32'd466,32'd-4323,32'd3110,32'd23,32'd-605,32'd5712,32'd-4719,32'd-2766,32'd2678,32'd2031,32'd1087,32'd-3588,32'd4003,32'd-8540,32'd-930,32'd-5083,32'd2258,32'd1115,32'd568,32'd2663,32'd-1838,32'd2319,32'd-6523,32'd4794,32'd5629,32'd7050,32'd2388,32'd-1077,32'd-832,32'd-7270,32'd1868,32'd1989,32'd-749,32'd1816,32'd837,32'd-3330,32'd-5703,32'd-253,32'd1052,32'd5947,32'd6069,32'd-3073,32'd-1674,32'd-92,32'd348,32'd-6743,32'd8232,32'd-698,32'd-3251,32'd-1326,32'd-659,32'd610,32'd-2763,32'd-235,32'd-5297,32'd3811,32'd-4934,32'd2144,32'd3295,32'd-4084,32'd332,32'd8940,32'd5576,32'd-2016,32'd1691,32'd-4760,32'd6743,32'd-4291,32'd-4370,32'd-3503,32'd1253,32'd-2824,32'd-1459,32'd1278,32'd-1102,32'd5078,32'd5322,32'd-6972,32'd-2457,32'd-3315,32'd579,32'd3276,32'd-3210,32'd-5761,32'd759,32'd-4106,32'd-2546,32'd3247,32'd-1429,32'd2495,32'd-2352,32'd-4929,32'd4926,32'd-1062,32'd2797,32'd-1481,32'd-4587,32'd-3679,32'd-3166,32'd2502,32'd-1706,32'd-3071,32'd8583,32'd-3215,32'd1351,32'd-1860,32'd-4360,32'd435,32'd778,32'd220,32'd4990};
    Wh[70]='{32'd-166,32'd2390,32'd-647,32'd2220,32'd1374,32'd2142,32'd3808,32'd2685,32'd4724,32'd3476,32'd292,32'd-1357,32'd-7021,32'd-1192,32'd4611,32'd949,32'd2919,32'd2341,32'd8681,32'd11699,32'd2951,32'd-1645,32'd1452,32'd1416,32'd3969,32'd-1818,32'd1660,32'd-1055,32'd5444,32'd1635,32'd3061,32'd-3728,32'd1307,32'd-1669,32'd1,32'd-2573,32'd-1098,32'd318,32'd-4240,32'd-102,32'd-354,32'd319,32'd-6030,32'd4770,32'd-2087,32'd1831,32'd13,32'd-2042,32'd8344,32'd-3823,32'd-3813,32'd-601,32'd6909,32'd5405,32'd-309,32'd444,32'd-4338,32'd6889,32'd4580,32'd849,32'd11435,32'd6601,32'd-5166,32'd2661,32'd-1137,32'd2536,32'd1174,32'd-2470,32'd3083,32'd-5224,32'd-520,32'd-3762,32'd-44,32'd1300,32'd4287,32'd-3144,32'd2551,32'd-1453,32'd1060,32'd-842,32'd1000,32'd337,32'd-2277,32'd-2753,32'd-1774,32'd-3261,32'd3823,32'd430,32'd209,32'd-1116,32'd6298,32'd895,32'd-3666,32'd-836,32'd-1005,32'd3229,32'd946,32'd-1071,32'd-563,32'd-1102,32'd64,32'd2675,32'd-2241,32'd1190,32'd3002,32'd-2095,32'd3654,32'd-3437,32'd-7871,32'd1292,32'd-2590,32'd-3869,32'd-2546,32'd1811,32'd1735,32'd616,32'd-191,32'd3237,32'd-12890,32'd2337,32'd-1778,32'd2073,32'd3444,32'd-1202,32'd1021,32'd5893,32'd3596,32'd-3146,32'd1864,32'd-5576,32'd7353,32'd665,32'd98,32'd-786,32'd628,32'd1784,32'd-1988,32'd-5,32'd838,32'd-548,32'd2166,32'd-2298,32'd-6054,32'd-50,32'd1319,32'd-3979,32'd-2277,32'd-9399,32'd-385,32'd3366,32'd3679,32'd-1590,32'd-7797,32'd775,32'd12832,32'd-2995,32'd-912,32'd1593,32'd-8408,32'd2944,32'd12783,32'd1881,32'd-674,32'd818,32'd-1488,32'd2580,32'd-3969,32'd-2115,32'd1496,32'd-778,32'd-4946,32'd778,32'd3005,32'd3115,32'd2524,32'd349,32'd712,32'd971,32'd4230,32'd-179,32'd2824,32'd1491,32'd-2988,32'd-2163,32'd4289,32'd2846,32'd-3173,32'd4704,32'd4934,32'd5952,32'd118,32'd2077,32'd720,32'd-2707,32'd-473,32'd-6518,32'd-2022,32'd-3647,32'd-4562,32'd1556,32'd3586,32'd102,32'd1823,32'd7031,32'd5937,32'd-1442,32'd-5434,32'd-1318,32'd71,32'd7792,32'd4960,32'd2025,32'd8134,32'd7968,32'd2932,32'd-2143,32'd963,32'd3039,32'd2115,32'd2102,32'd-1015,32'd2152,32'd2403,32'd7714,32'd4633,32'd4492,32'd-1749,32'd-2498,32'd1756,32'd4116,32'd2117,32'd1817,32'd-2819,32'd-1434,32'd3239,32'd4667,32'd387,32'd-2119,32'd856,32'd3027,32'd3815,32'd-3037,32'd9682,32'd-4670,32'd3269,32'd6967,32'd-2210,32'd-573,32'd3935,32'd-63,32'd-3061,32'd2447,32'd3845,32'd-437,32'd4582,32'd81,32'd-3293,32'd-6376,32'd5488,32'd8422,32'd625,32'd1909,32'd-6401,32'd2719,32'd-612,32'd4667,32'd3088,32'd1756,32'd1488,32'd-2094,32'd1656,32'd-1176,32'd1723,32'd1994,32'd-1069,32'd1724,32'd54,32'd-116,32'd3085,32'd2624,32'd-3886,32'd1168,32'd432,32'd-320,32'd-583,32'd-3281,32'd-1525,32'd-3229,32'd318,32'd-4223,32'd-3232,32'd4157,32'd-2727,32'd2487,32'd3195,32'd3398,32'd-124,32'd-2529,32'd-2973,32'd3703,32'd4592,32'd0,32'd-438,32'd-1868,32'd3942,32'd5161,32'd6127,32'd-611,32'd7622,32'd4616,32'd-4709,32'd2281,32'd3693,32'd7319,32'd1478,32'd3142,32'd-2102,32'd-963,32'd2456,32'd-4260,32'd-2561,32'd3803,32'd-570,32'd2211,32'd7153,32'd12753,32'd9599,32'd-5039,32'd-1629,32'd-1333,32'd980,32'd-258,32'd2749,32'd3508,32'd-257,32'd4130,32'd493,32'd2846,32'd1193,32'd701,32'd728,32'd1936,32'd-5517,32'd-350,32'd-917,32'd1093,32'd1992,32'd6196,32'd1798,32'd-178,32'd-2352,32'd5830,32'd510,32'd3942,32'd-7631,32'd-4812,32'd404,32'd-1790,32'd546,32'd786,32'd13076,32'd1140,32'd785,32'd1795,32'd1708,32'd6782,32'd2485,32'd-81,32'd-251,32'd-1178,32'd3154,32'd2175,32'd-851,32'd714,32'd7504,32'd5361,32'd-2546,32'd1588,32'd1433,32'd-1197,32'd-1708,32'd-3674,32'd-310,32'd7211,32'd-3666,32'd-1667,32'd977,32'd-1284,32'd-5180,32'd-591,32'd-9047,32'd5917,32'd9057,32'd-681,32'd-1942,32'd-7407,32'd-3762,32'd-2871,32'd2768,32'd905};
    Wh[71]='{32'd-363,32'd-1726,32'd-3273,32'd4760,32'd-168,32'd-1087,32'd2653,32'd-5747,32'd2022,32'd1372,32'd3774,32'd-248,32'd5620,32'd8486,32'd-1640,32'd2736,32'd1447,32'd-2242,32'd105,32'd1222,32'd-5830,32'd153,32'd3852,32'd709,32'd-1583,32'd-5195,32'd2158,32'd877,32'd5258,32'd3732,32'd-3139,32'd-1939,32'd5185,32'd2227,32'd-479,32'd-1746,32'd4028,32'd2546,32'd5375,32'd-1854,32'd236,32'd1113,32'd-1204,32'd4138,32'd-1547,32'd-3923,32'd4169,32'd-2912,32'd-2491,32'd-1995,32'd2580,32'd-3063,32'd1638,32'd-5415,32'd-4091,32'd5278,32'd-3984,32'd-1536,32'd-2322,32'd-3103,32'd-680,32'd-1201,32'd5717,32'd-1304,32'd-602,32'd2183,32'd-3120,32'd-5571,32'd891,32'd-4824,32'd-5517,32'd5122,32'd1162,32'd-2680,32'd-150,32'd-3349,32'd1877,32'd1244,32'd-8779,32'd-329,32'd207,32'd-721,32'd-179,32'd100,32'd328,32'd362,32'd941,32'd688,32'd967,32'd-1787,32'd-3315,32'd-3754,32'd-3752,32'd3210,32'd-2426,32'd-3952,32'd-1800,32'd-3828,32'd2325,32'd-2658,32'd2031,32'd-795,32'd6176,32'd11679,32'd236,32'd643,32'd538,32'd465,32'd-2541,32'd3615,32'd-274,32'd1826,32'd-6782,32'd-1314,32'd5346,32'd-2476,32'd-4606,32'd4731,32'd-197,32'd2575,32'd-5126,32'd-5019,32'd-3576,32'd-1470,32'd2000,32'd7778,32'd4580,32'd-2153,32'd-416,32'd-462,32'd1217,32'd-1,32'd-521,32'd-7202,32'd2875,32'd3427,32'd-3623,32'd-3854,32'd3139,32'd1763,32'd-1350,32'd1378,32'd254,32'd-2105,32'd178,32'd1262,32'd1672,32'd-1007,32'd-1549,32'd1192,32'd-2434,32'd2000,32'd-3513,32'd-2895,32'd1128,32'd-6298,32'd-5844,32'd1324,32'd4355,32'd-5629,32'd-1978,32'd-253,32'd3403,32'd7636,32'd89,32'd6718,32'd5336,32'd-3867,32'd728,32'd-562,32'd-7089,32'd-606,32'd5727,32'd820,32'd-798,32'd969,32'd1372,32'd-6948,32'd-1859,32'd298,32'd9165,32'd-6406,32'd1760,32'd-3615,32'd-2358,32'd5649,32'd1568,32'd31,32'd-1589,32'd-1701,32'd94,32'd767,32'd5732,32'd-1129,32'd1932,32'd4887,32'd-1116,32'd-195,32'd-6245,32'd3327,32'd-997,32'd-1058,32'd-3601,32'd-4401,32'd8608,32'd-1440,32'd-1093,32'd5068,32'd6469,32'd2807,32'd1723,32'd2792,32'd-1986,32'd-2578,32'd-276,32'd5961,32'd1221,32'd-579,32'd-2700,32'd-1694,32'd618,32'd2181,32'd-6923,32'd-2016,32'd4221,32'd1282,32'd459,32'd-2795,32'd3051,32'd5180,32'd-853,32'd738,32'd4401,32'd860,32'd3020,32'd7680,32'd5766,32'd-183,32'd-1323,32'd368,32'd2178,32'd-6835,32'd4091,32'd1871,32'd-61,32'd-1668,32'd-1889,32'd-5024,32'd630,32'd1342,32'd629,32'd-689,32'd1171,32'd-1043,32'd1343,32'd671,32'd146,32'd133,32'd-4245,32'd-2031,32'd2197,32'd2012,32'd1039,32'd1535,32'd5742,32'd-3410,32'd-1315,32'd1750,32'd-565,32'd-960,32'd3479,32'd1326,32'd-1782,32'd561,32'd-3132,32'd422,32'd1530,32'd963,32'd2856,32'd336,32'd2573,32'd1091,32'd1697,32'd2099,32'd-4492,32'd5590,32'd5024,32'd-1859,32'd-1811,32'd4804,32'd8725,32'd-5615,32'd1923,32'd-9677,32'd-9746,32'd22,32'd1061,32'd645,32'd2966,32'd5039,32'd1824,32'd-5683,32'd-1304,32'd6547,32'd434,32'd-1456,32'd3117,32'd-3125,32'd-1947,32'd-1431,32'd-6992,32'd-79,32'd-3459,32'd-1677,32'd-3120,32'd-5292,32'd3015,32'd29,32'd5239,32'd2342,32'd-2298,32'd4042,32'd1424,32'd-3549,32'd7412,32'd1567,32'd2226,32'd-2053,32'd2724,32'd1948,32'd5239,32'd-1079,32'd-3618,32'd5112,32'd-3518,32'd733,32'd-1358,32'd6694,32'd-4545,32'd-208,32'd-1171,32'd3376,32'd715,32'd-3186,32'd-7661,32'd3044,32'd-1083,32'd-2822,32'd-3342,32'd-3061,32'd642,32'd-3005,32'd2337,32'd-2839,32'd1909,32'd-1970,32'd2587,32'd56,32'd-2286,32'd-2331,32'd-866,32'd-3312,32'd1933,32'd2166,32'd-1967,32'd4616,32'd8696,32'd-996,32'd-945,32'd-4052,32'd1222,32'd-6928,32'd10166,32'd-8662,32'd7089,32'd1318,32'd1466,32'd104,32'd-2597,32'd4555,32'd-3293,32'd2617,32'd5576,32'd902,32'd830,32'd3225,32'd2871,32'd2631,32'd-2233,32'd7080,32'd-3579,32'd-7802,32'd-301,32'd6245,32'd3322,32'd6357,32'd1719,32'd-2215,32'd1128,32'd3891};
    Wh[72]='{32'd993,32'd-1529,32'd-1395,32'd683,32'd5786,32'd206,32'd-1035,32'd-2226,32'd-306,32'd-783,32'd-5932,32'd-2459,32'd135,32'd-4621,32'd-6220,32'd-5673,32'd433,32'd2734,32'd363,32'd2066,32'd-775,32'd-2432,32'd-689,32'd-1459,32'd5346,32'd445,32'd92,32'd-351,32'd314,32'd-580,32'd820,32'd-1328,32'd1805,32'd-1812,32'd1571,32'd-4135,32'd4123,32'd-2381,32'd-934,32'd-4641,32'd-664,32'd-1517,32'd1745,32'd-5947,32'd-524,32'd1813,32'd-826,32'd1184,32'd-2006,32'd1077,32'd0,32'd-2844,32'd796,32'd2457,32'd1696,32'd-4140,32'd-3305,32'd971,32'd2387,32'd-4941,32'd4812,32'd3828,32'd-631,32'd-1619,32'd-1064,32'd142,32'd2315,32'd-1148,32'd-24,32'd-2274,32'd3037,32'd-1232,32'd-5332,32'd-244,32'd-2170,32'd-2058,32'd124,32'd-853,32'd5087,32'd790,32'd-1826,32'd-1674,32'd-4545,32'd-4238,32'd-2056,32'd1089,32'd-188,32'd-2529,32'd-3034,32'd-1125,32'd1547,32'd-8496,32'd2683,32'd-2177,32'd-5737,32'd-2215,32'd-3569,32'd-2575,32'd770,32'd-3845,32'd-3005,32'd512,32'd3129,32'd3229,32'd7099,32'd-706,32'd2839,32'd5107,32'd-1268,32'd-2553,32'd-237,32'd-5034,32'd-228,32'd-3334,32'd-1210,32'd-8222,32'd221,32'd-1931,32'd-1433,32'd-885,32'd2144,32'd2705,32'd-4360,32'd575,32'd4025,32'd85,32'd1707,32'd-4172,32'd2337,32'd-2028,32'd335,32'd-4831,32'd68,32'd482,32'd2941,32'd3808,32'd3361,32'd-4775,32'd-4873,32'd-1981,32'd2897,32'd-3898,32'd-2565,32'd1250,32'd1215,32'd5405,32'd5151,32'd-5288,32'd-5039,32'd-838,32'd1853,32'd487,32'd3332,32'd-9858,32'd-2866,32'd4238,32'd2386,32'd-447,32'd2810,32'd-6513,32'd-4174,32'd-604,32'd-292,32'd50,32'd-3752,32'd-4484,32'd-1281,32'd5405,32'd156,32'd1278,32'd-787,32'd1674,32'd-1536,32'd-3449,32'd2448,32'd1502,32'd-528,32'd1516,32'd256,32'd-1337,32'd6909,32'd-3627,32'd4636,32'd2012,32'd-74,32'd167,32'd3742,32'd2751,32'd6660,32'd2951,32'd4,32'd1466,32'd1429,32'd4697,32'd193,32'd4943,32'd1441,32'd-2839,32'd5234,32'd1582,32'd1499,32'd4963,32'd-541,32'd3144,32'd6269,32'd342,32'd4455,32'd-16,32'd-9482,32'd-504,32'd158,32'd1877,32'd1346,32'd3518,32'd2019,32'd8837,32'd1864,32'd-209,32'd-1523,32'd13,32'd-66,32'd974,32'd-357,32'd-1280,32'd-614,32'd-791,32'd3803,32'd1474,32'd-302,32'd-2119,32'd1604,32'd-203,32'd513,32'd3273,32'd-8125,32'd1218,32'd2402,32'd3269,32'd1326,32'd1169,32'd-1855,32'd-4006,32'd-3884,32'd6113,32'd-1430,32'd3510,32'd-4572,32'd637,32'd-4428,32'd547,32'd-3308,32'd-2210,32'd2475,32'd128,32'd3393,32'd341,32'd-322,32'd4511,32'd-383,32'd-17,32'd1087,32'd-1160,32'd544,32'd-4133,32'd-359,32'd-3559,32'd505,32'd-259,32'd-682,32'd-294,32'd-3889,32'd5688,32'd-6215,32'd812,32'd-2602,32'd1621,32'd3315,32'd-660,32'd1095,32'd-1940,32'd-1270,32'd7163,32'd-3237,32'd8671,32'd4533,32'd1187,32'd-584,32'd6562,32'd3923,32'd-66,32'd-2036,32'd10781,32'd66,32'd1030,32'd3217,32'd1479,32'd3859,32'd-2941,32'd8193,32'd-1837,32'd3776,32'd2260,32'd327,32'd1121,32'd7807,32'd-3525,32'd1457,32'd-1550,32'd-4050,32'd-2651,32'd1033,32'd-471,32'd-1061,32'd-4584,32'd-1510,32'd-3288,32'd823,32'd-2182,32'd-197,32'd225,32'd-9443,32'd-183,32'd664,32'd-218,32'd3149,32'd-416,32'd-654,32'd-266,32'd8037,32'd-4270,32'd1094,32'd1816,32'd-2895,32'd6245,32'd1568,32'd-2507,32'd1945,32'd-5688,32'd3286,32'd1072,32'd-2304,32'd3051,32'd-4199,32'd-14,32'd5625,32'd1911,32'd-1112,32'd1495,32'd829,32'd-2668,32'd352,32'd1947,32'd-1787,32'd-1486,32'd4768,32'd-988,32'd-1759,32'd-3166,32'd3603,32'd-2498,32'd2015,32'd-2858,32'd1700,32'd-195,32'd2121,32'd-5776,32'd-881,32'd4482,32'd917,32'd-3159,32'd-2617,32'd5849,32'd-244,32'd-809,32'd-50,32'd5024,32'd-198,32'd915,32'd-933,32'd1464,32'd-1641,32'd4807,32'd4941,32'd-2485,32'd2514,32'd2551,32'd-3740,32'd559,32'd245,32'd-6313,32'd-741,32'd980,32'd2408,32'd-513,32'd-6523,32'd-2261,32'd-4511,32'd-2807,32'd-5327,32'd2951};
    Wh[73]='{32'd-1386,32'd-897,32'd-1396,32'd-476,32'd-40,32'd2263,32'd3083,32'd-146,32'd1929,32'd-216,32'd6855,32'd-4580,32'd497,32'd4272,32'd-375,32'd839,32'd-4892,32'd-1192,32'd-258,32'd1146,32'd-3591,32'd131,32'd1138,32'd2658,32'd611,32'd-306,32'd-61,32'd-2169,32'd2028,32'd2712,32'd6088,32'd4020,32'd7421,32'd1285,32'd-809,32'd452,32'd-948,32'd4028,32'd-3784,32'd-1611,32'd1566,32'd-3232,32'd1710,32'd751,32'd3679,32'd-2169,32'd-3054,32'd-2187,32'd2106,32'd884,32'd2124,32'd-1123,32'd266,32'd502,32'd421,32'd1093,32'd4631,32'd-3623,32'd466,32'd8012,32'd1846,32'd4272,32'd2993,32'd-3173,32'd1763,32'd591,32'd1488,32'd1130,32'd95,32'd-2136,32'd-3593,32'd397,32'd5297,32'd-2147,32'd588,32'd-2653,32'd1912,32'd-3979,32'd1531,32'd6865,32'd-1520,32'd-4357,32'd-252,32'd-1020,32'd-1888,32'd922,32'd-68,32'd2456,32'd2907,32'd880,32'd-162,32'd437,32'd3325,32'd-1711,32'd-261,32'd1199,32'd1129,32'd-406,32'd-513,32'd358,32'd3857,32'd-1251,32'd2861,32'd-5043,32'd-2844,32'd228,32'd6220,32'd-25,32'd2802,32'd-1976,32'd1738,32'd-6835,32'd7744,32'd733,32'd3317,32'd2266,32'd4099,32'd2600,32'd1800,32'd-186,32'd-1298,32'd174,32'd-4755,32'd110,32'd3886,32'd2149,32'd3168,32'd-524,32'd1370,32'd-4912,32'd-6977,32'd4819,32'd-4260,32'd-4812,32'd-7758,32'd2556,32'd7167,32'd-6318,32'd-4155,32'd1011,32'd899,32'd1072,32'd811,32'd-1011,32'd-2849,32'd4211,32'd-3305,32'd4643,32'd4641,32'd4926,32'd-1815,32'd-91,32'd-547,32'd6147,32'd-299,32'd-4704,32'd-1051,32'd-259,32'd3867,32'd-6113,32'd-5249,32'd3359,32'd4760,32'd1091,32'd3950,32'd-2841,32'd-2049,32'd1624,32'd731,32'd767,32'd-1368,32'd1093,32'd6752,32'd-2736,32'd1834,32'd184,32'd-1213,32'd595,32'd-892,32'd-953,32'd-1264,32'd3295,32'd-532,32'd366,32'd1188,32'd1177,32'd2585,32'd-391,32'd-4516,32'd1784,32'd1341,32'd293,32'd3188,32'd2066,32'd-4338,32'd-881,32'd-2491,32'd541,32'd7695,32'd-3020,32'd1435,32'd100,32'd-5395,32'd1159,32'd4277,32'd-460,32'd501,32'd181,32'd5717,32'd1629,32'd-1774,32'd7729,32'd1927,32'd-1475,32'd239,32'd-874,32'd-947,32'd-4042,32'd-2222,32'd-5566,32'd-1291,32'd6166,32'd1512,32'd-4892,32'd-474,32'd4020,32'd6157,32'd-3994,32'd515,32'd-9106,32'd-3027,32'd462,32'd4218,32'd-2292,32'd-1034,32'd6025,32'd-3867,32'd720,32'd4431,32'd5449,32'd-4338,32'd-2088,32'd1467,32'd3229,32'd-3039,32'd2211,32'd70,32'd-2822,32'd2509,32'd2890,32'd-3652,32'd-570,32'd23,32'd-3122,32'd-4733,32'd-6420,32'd1368,32'd3278,32'd4665,32'd-10019,32'd1065,32'd2805,32'd-3610,32'd2946,32'd1339,32'd-426,32'd-621,32'd1796,32'd-1107,32'd-9614,32'd2619,32'd4428,32'd1950,32'd1828,32'd-1015,32'd502,32'd-2512,32'd-2133,32'd72,32'd1036,32'd2802,32'd5361,32'd2700,32'd2702,32'd1253,32'd2885,32'd-1185,32'd488,32'd2910,32'd-722,32'd-3237,32'd1910,32'd-3205,32'd-2578,32'd-299,32'd-3413,32'd575,32'd-1015,32'd3103,32'd1594,32'd2673,32'd-4934,32'd2006,32'd-2741,32'd-4096,32'd1103,32'd-8002,32'd-2406,32'd-822,32'd-3439,32'd-2626,32'd-5366,32'd5937,32'd4470,32'd1256,32'd2687,32'd5019,32'd-6699,32'd442,32'd-6416,32'd-178,32'd3537,32'd2302,32'd-3864,32'd-1246,32'd3798,32'd3547,32'd-3325,32'd337,32'd-1462,32'd2360,32'd2712,32'd2919,32'd3671,32'd-598,32'd3505,32'd-252,32'd944,32'd491,32'd-3674,32'd280,32'd-658,32'd-637,32'd-3161,32'd-2202,32'd-2788,32'd-422,32'd2482,32'd-4787,32'd1317,32'd-1340,32'd734,32'd-257,32'd616,32'd1879,32'd-58,32'd10556,32'd4147,32'd-7714,32'd1745,32'd-2919,32'd2091,32'd399,32'd6918,32'd-853,32'd18,32'd792,32'd2004,32'd-2451,32'd-6376,32'd-747,32'd5263,32'd3715,32'd-4160,32'd1621,32'd-3212,32'd3735,32'd-1542,32'd-1111,32'd3996,32'd-1781,32'd4643,32'd-6889,32'd2673,32'd-2958,32'd-1864,32'd-3693,32'd1372,32'd-562,32'd-1805,32'd-1364,32'd105,32'd-1770,32'd182,32'd-5532,32'd-2216,32'd1843,32'd-1210,32'd-1222,32'd2136};
    Wh[74]='{32'd230,32'd-1034,32'd-1254,32'd-325,32'd-2612,32'd-1428,32'd5019,32'd-946,32'd85,32'd-961,32'd-905,32'd-686,32'd2573,32'd2744,32'd-4208,32'd-1820,32'd2,32'd3156,32'd2012,32'd2944,32'd-1407,32'd1728,32'd3576,32'd-216,32'd-2030,32'd1729,32'd-2844,32'd75,32'd2111,32'd81,32'd-870,32'd9624,32'd3513,32'd-773,32'd-326,32'd1345,32'd-854,32'd-784,32'd3867,32'd373,32'd-733,32'd-1730,32'd3017,32'd-48,32'd4787,32'd5512,32'd-3041,32'd902,32'd-1333,32'd990,32'd678,32'd-2302,32'd520,32'd2695,32'd-922,32'd-1317,32'd-1221,32'd-179,32'd-1970,32'd2609,32'd3068,32'd3767,32'd2651,32'd-1538,32'd-2014,32'd1043,32'd222,32'd294,32'd-61,32'd-115,32'd4426,32'd786,32'd-498,32'd-1820,32'd-129,32'd1972,32'd2988,32'd-1152,32'd6586,32'd-3793,32'd-2155,32'd-3969,32'd2349,32'd-3391,32'd1275,32'd170,32'd-1006,32'd-2062,32'd2668,32'd884,32'd-126,32'd-1383,32'd-939,32'd217,32'd1967,32'd-896,32'd304,32'd-1680,32'd1435,32'd2749,32'd-459,32'd2636,32'd2966,32'd707,32'd1365,32'd66,32'd1673,32'd6586,32'd4711,32'd1370,32'd-308,32'd-2307,32'd3618,32'd2186,32'd-2741,32'd-786,32'd-2739,32'd3093,32'd-5385,32'd-1165,32'd2427,32'd902,32'd-639,32'd-2023,32'd-5380,32'd-1536,32'd-2485,32'd2322,32'd7451,32'd-3078,32'd-2998,32'd-2083,32'd9028,32'd-310,32'd3688,32'd2275,32'd-3364,32'd-1893,32'd-369,32'd-3208,32'd178,32'd-764,32'd-720,32'd2575,32'd4777,32'd-567,32'd1680,32'd4270,32'd-264,32'd1512,32'd-1673,32'd-2458,32'd-1097,32'd-404,32'd-380,32'd1785,32'd3269,32'd-1312,32'd-568,32'd-5771,32'd-3232,32'd3320,32'd-839,32'd-3837,32'd-1915,32'd-509,32'd-2309,32'd-4064,32'd198,32'd153,32'd-4936,32'd-2285,32'd447,32'd-1145,32'd-42,32'd-1583,32'd-1715,32'd-520,32'd-1286,32'd255,32'd-1751,32'd-3349,32'd2108,32'd-5327,32'd-977,32'd2529,32'd1237,32'd-339,32'd3688,32'd3674,32'd-751,32'd1575,32'd-2687,32'd6025,32'd1650,32'd-4355,32'd254,32'd-5776,32'd-427,32'd2814,32'd1617,32'd718,32'd-2135,32'd-1387,32'd-3752,32'd2023,32'd-726,32'd758,32'd-717,32'd1322,32'd-2416,32'd590,32'd-760,32'd482,32'd809,32'd-7041,32'd6489,32'd56,32'd-327,32'd6083,32'd790,32'd2027,32'd-4992,32'd568,32'd2570,32'd-1777,32'd-996,32'd989,32'd3627,32'd-2385,32'd-4350,32'd3757,32'd-7036,32'd-1760,32'd-5737,32'd1179,32'd1348,32'd-521,32'd-2261,32'd4296,32'd-168,32'd4526,32'd-1578,32'd2287,32'd886,32'd1600,32'd1064,32'd1809,32'd-1201,32'd1625,32'd-30,32'd-3068,32'd3527,32'd623,32'd-913,32'd-1533,32'd-299,32'd-1800,32'd-1485,32'd-3476,32'd-4968,32'd-6860,32'd-1230,32'd-5703,32'd-4426,32'd-368,32'd-1845,32'd-5092,32'd-378,32'd969,32'd2636,32'd579,32'd-4128,32'd-284,32'd-1503,32'd-522,32'd-1794,32'd-805,32'd86,32'd-1119,32'd-3542,32'd1052,32'd1975,32'd4382,32'd426,32'd-7500,32'd264,32'd-2215,32'd-6000,32'd-1933,32'd-5576,32'd-2702,32'd-412,32'd4550,32'd-1224,32'd-4245,32'd-57,32'd-1654,32'd680,32'd-914,32'd578,32'd-3540,32'd-1386,32'd3034,32'd-1910,32'd-4987,32'd574,32'd-933,32'd1322,32'd1300,32'd1558,32'd1520,32'd-1861,32'd55,32'd1649,32'd-507,32'd7871,32'd-17,32'd-6186,32'd2327,32'd-4707,32'd1067,32'd2497,32'd1444,32'd-1405,32'd-3041,32'd-2661,32'd-1223,32'd-1053,32'd1373,32'd-5927,32'd1373,32'd3063,32'd1018,32'd2437,32'd-4555,32'd208,32'd-1810,32'd-2143,32'd155,32'd-2197,32'd-2165,32'd1126,32'd5170,32'd-53,32'd2666,32'd7490,32'd-3247,32'd-3405,32'd4074,32'd3903,32'd2587,32'd783,32'd383,32'd859,32'd577,32'd-1729,32'd-13154,32'd-3012,32'd1486,32'd1507,32'd-1761,32'd-48,32'd-2318,32'd1313,32'd2507,32'd-4633,32'd3225,32'd-3471,32'd-6230,32'd5732,32'd-3974,32'd-1818,32'd-3283,32'd-140,32'd-1381,32'd5712,32'd-620,32'd661,32'd574,32'd-4826,32'd484,32'd6826,32'd4450,32'd-3745,32'd3625,32'd614,32'd112,32'd-254,32'd1148,32'd1624,32'd6318,32'd31,32'd6323,32'd-1505,32'd-11240,32'd-1284,32'd-288,32'd367,32'd-425};
    Wh[75]='{32'd1921,32'd2963,32'd-662,32'd1229,32'd798,32'd-1553,32'd-2521,32'd-440,32'd1339,32'd-2175,32'd409,32'd-709,32'd-5751,32'd-1512,32'd-5019,32'd2324,32'd-4826,32'd968,32'd2445,32'd-1824,32'd242,32'd1423,32'd-6694,32'd-543,32'd565,32'd-212,32'd-1669,32'd-1838,32'd-6391,32'd1159,32'd2338,32'd2342,32'd-594,32'd-4099,32'd-2232,32'd-3796,32'd1346,32'd-2502,32'd-3071,32'd-5039,32'd-977,32'd-387,32'd1680,32'd-3481,32'd3132,32'd1038,32'd2597,32'd1450,32'd-4611,32'd1689,32'd-404,32'd3989,32'd-9785,32'd-1633,32'd1336,32'd-564,32'd-2480,32'd-2700,32'd1678,32'd-2210,32'd-1652,32'd29,32'd-668,32'd394,32'd-5429,32'd-117,32'd209,32'd-908,32'd3874,32'd-159,32'd2423,32'd-3637,32'd3359,32'd2302,32'd1418,32'd2502,32'd-4189,32'd2307,32'd-127,32'd1534,32'd-1248,32'd-5781,32'd505,32'd-7075,32'd3820,32'd-2731,32'd24,32'd578,32'd4492,32'd1413,32'd100,32'd-5175,32'd592,32'd-2619,32'd2739,32'd1069,32'd429,32'd-368,32'd-8627,32'd-2213,32'd-4045,32'd-704,32'd-3088,32'd-7246,32'd615,32'd-110,32'd-900,32'd670,32'd1352,32'd-2590,32'd-1992,32'd-10585,32'd-463,32'd2418,32'd2441,32'd2622,32'd3803,32'd4230,32'd-4953,32'd-659,32'd616,32'd-2479,32'd-2093,32'd-2568,32'd-5927,32'd2512,32'd529,32'd10947,32'd-1697,32'd-5380,32'd-1719,32'd359,32'd1911,32'd-938,32'd-196,32'd-3083,32'd116,32'd-1227,32'd1152,32'd-1711,32'd5859,32'd-1340,32'd-3254,32'd2064,32'd1190,32'd2666,32'd505,32'd-2792,32'd4243,32'd-4445,32'd3615,32'd2080,32'd-764,32'd4455,32'd3359,32'd-1883,32'd-1254,32'd2305,32'd500,32'd-1112,32'd3579,32'd-3593,32'd71,32'd-1583,32'd4758,32'd343,32'd-2792,32'd650,32'd-6972,32'd2196,32'd1832,32'd3088,32'd4506,32'd4016,32'd1091,32'd-479,32'd55,32'd5947,32'd-3022,32'd1549,32'd5634,32'd-2304,32'd-520,32'd350,32'd1259,32'd3193,32'd-790,32'd-2797,32'd2875,32'd803,32'd-134,32'd4448,32'd2551,32'd-4384,32'd-4082,32'd-297,32'd1385,32'd-292,32'd-2454,32'd-2250,32'd-586,32'd957,32'd5336,32'd-7666,32'd353,32'd-1301,32'd250,32'd429,32'd-4448,32'd1654,32'd-5537,32'd3041,32'd-2028,32'd-5390,32'd-2922,32'd-162,32'd-3574,32'd2459,32'd-426,32'd-13964,32'd2475,32'd997,32'd-252,32'd-2203,32'd-1031,32'd790,32'd4262,32'd-833,32'd2237,32'd-807,32'd1117,32'd476,32'd3833,32'd326,32'd-2093,32'd544,32'd-1816,32'd2207,32'd3308,32'd3627,32'd10800,32'd-1107,32'd-592,32'd2590,32'd4262,32'd-2180,32'd290,32'd-2971,32'd-3637,32'd3137,32'd-82,32'd4375,32'd-44,32'd-114,32'd2924,32'd-1268,32'd1999,32'd-2083,32'd4626,32'd-2580,32'd-1934,32'd-3405,32'd5771,32'd-1071,32'd-1635,32'd-3125,32'd-2939,32'd3845,32'd-3562,32'd3295,32'd-2113,32'd-737,32'd-1677,32'd-1763,32'd-3991,32'd-2103,32'd3625,32'd2294,32'd4201,32'd-334,32'd-1480,32'd-1771,32'd-7792,32'd-6137,32'd-3083,32'd-228,32'd413,32'd5141,32'd834,32'd1700,32'd-4748,32'd8349,32'd1247,32'd-3610,32'd-2924,32'd-7036,32'd4724,32'd1866,32'd-6948,32'd280,32'd-386,32'd-2578,32'd3837,32'd-3327,32'd4741,32'd-4086,32'd-1785,32'd-2692,32'd-1070,32'd1787,32'd-346,32'd-1741,32'd-3508,32'd12812,32'd571,32'd4926,32'd-3339,32'd89,32'd-6235,32'd-4248,32'd4956,32'd-1722,32'd-8916,32'd-5151,32'd-4155,32'd-5800,32'd4350,32'd2486,32'd-1196,32'd-4531,32'd-5903,32'd-1966,32'd-2788,32'd-1233,32'd246,32'd-5239,32'd3291,32'd-5527,32'd5122,32'd-469,32'd1796,32'd-596,32'd-728,32'd-4377,32'd-311,32'd-125,32'd-2320,32'd5058,32'd2983,32'd275,32'd-3679,32'd613,32'd2744,32'd2222,32'd3178,32'd-558,32'd2912,32'd8002,32'd6289,32'd886,32'd732,32'd428,32'd3410,32'd3305,32'd335,32'd-1719,32'd3530,32'd-5263,32'd-3098,32'd-12470,32'd-4316,32'd-3676,32'd3579,32'd-1781,32'd-5634,32'd1759,32'd222,32'd226,32'd608,32'd1004,32'd-3215,32'd1042,32'd930,32'd-801,32'd-1468,32'd1712,32'd441,32'd4372,32'd-1188,32'd-2349,32'd-7031,32'd-1104,32'd3327,32'd-3527,32'd4152,32'd-144,32'd-2275,32'd2403,32'd-314,32'd-2521};
    Wh[76]='{32'd-4970,32'd1343,32'd3413,32'd6181,32'd1835,32'd-1668,32'd49,32'd3625,32'd8696,32'd186,32'd5415,32'd2641,32'd520,32'd-2092,32'd4384,32'd1466,32'd1746,32'd2265,32'd1611,32'd1120,32'd-4047,32'd1568,32'd2463,32'd1213,32'd-4221,32'd-4013,32'd2386,32'd231,32'd2612,32'd7275,32'd2102,32'd3535,32'd3754,32'd950,32'd1,32'd615,32'd-2044,32'd-1416,32'd1494,32'd-2541,32'd-6,32'd1104,32'd536,32'd-1309,32'd-5258,32'd4592,32'd9663,32'd-1937,32'd1737,32'd2697,32'd-181,32'd-1231,32'd-2807,32'd3937,32'd1804,32'd1879,32'd3771,32'd-1055,32'd-3173,32'd4401,32'd2354,32'd-2224,32'd783,32'd4074,32'd-1350,32'd2829,32'd-3691,32'd1240,32'd3007,32'd-5019,32'd-2296,32'd-3491,32'd-447,32'd-321,32'd4157,32'd4816,32'd-6181,32'd462,32'd-1826,32'd-4936,32'd-2133,32'd1151,32'd-2546,32'd4716,32'd-3627,32'd6127,32'd820,32'd1993,32'd3505,32'd-3208,32'd2619,32'd2788,32'd-1665,32'd433,32'd-7949,32'd3771,32'd-5048,32'd822,32'd717,32'd-2352,32'd4631,32'd6166,32'd-1779,32'd2666,32'd-1314,32'd2357,32'd3542,32'd10390,32'd11962,32'd-1973,32'd5014,32'd11552,32'd4853,32'd-5532,32'd-565,32'd-3530,32'd2927,32'd17558,32'd-1445,32'd-1790,32'd-3991,32'd-6767,32'd-9555,32'd-1032,32'd3337,32'd-8750,32'd4133,32'd-187,32'd2675,32'd3923,32'd4047,32'd-7500,32'd-3342,32'd-1917,32'd1904,32'd5258,32'd-8413,32'd-575,32'd-114,32'd-1176,32'd-3884,32'd5571,32'd11992,32'd-3449,32'd3945,32'd-3583,32'd8095,32'd-9648,32'd13125,32'd1314,32'd960,32'd2875,32'd-1855,32'd5815,32'd706,32'd-9291,32'd-6752,32'd3718,32'd5883,32'd-2104,32'd-7539,32'd-5092,32'd-2470,32'd4494,32'd-3801,32'd-7871,32'd3925,32'd519,32'd4831,32'd-6284,32'd7265,32'd7475,32'd-3896,32'd2100,32'd1760,32'd-2954,32'd-1149,32'd271,32'd7441,32'd2033,32'd9672,32'd-8881,32'd6098,32'd-2785,32'd-732,32'd1541,32'd5278,32'd2978,32'd4291,32'd-7500,32'd-8574,32'd-3259,32'd-1358,32'd4528,32'd6870,32'd8222,32'd-704,32'd713,32'd2512,32'd-3847,32'd-1285,32'd3322,32'd-475,32'd2929,32'd5322,32'd-1713,32'd-708,32'd-4118,32'd3315,32'd2868,32'd-7749,32'd2303,32'd-1039,32'd7265,32'd-4851,32'd-2622,32'd2797,32'd1560,32'd3811,32'd350,32'd-2783,32'd-808,32'd2624,32'd-5966,32'd3112,32'd111,32'd682,32'd-2644,32'd-3308,32'd-3745,32'd-912,32'd-406,32'd-2822,32'd1130,32'd-4074,32'd1955,32'd-7612,32'd497,32'd4687,32'd-290,32'd183,32'd4387,32'd-621,32'd-540,32'd1405,32'd4851,32'd2810,32'd2213,32'd249,32'd-422,32'd-6157,32'd-2482,32'd5756,32'd3583,32'd2321,32'd-9067,32'd-1838,32'd-1796,32'd176,32'd-6411,32'd507,32'd889,32'd1729,32'd-7006,32'd139,32'd-1431,32'd-6801,32'd-3356,32'd-2242,32'd1484,32'd1304,32'd2709,32'd3571,32'd1557,32'd560,32'd-7441,32'd2414,32'd-3850,32'd4367,32'd-631,32'd4238,32'd4467,32'd-5380,32'd2629,32'd-6650,32'd-7978,32'd-1248,32'd2093,32'd-2900,32'd-185,32'd1033,32'd-7539,32'd-8754,32'd-1401,32'd2697,32'd218,32'd-4721,32'd-1810,32'd-5815,32'd46,32'd2800,32'd-2907,32'd7377,32'd5209,32'd2595,32'd2019,32'd5400,32'd-763,32'd2810,32'd-613,32'd4042,32'd6166,32'd-5053,32'd5327,32'd1010,32'd1026,32'd9150,32'd480,32'd6342,32'd2531,32'd8100,32'd4492,32'd3413,32'd-3874,32'd3598,32'd4265,32'd3776,32'd-4497,32'd632,32'd4626,32'd7744,32'd3276,32'd-1384,32'd1039,32'd-2314,32'd2071,32'd-2398,32'd-2373,32'd1044,32'd-5410,32'd-1656,32'd-1035,32'd415,32'd-4453,32'd-4758,32'd2539,32'd-176,32'd-1490,32'd7377,32'd-3105,32'd-2299,32'd-3886,32'd-830,32'd-924,32'd3176,32'd2441,32'd1983,32'd-2247,32'd2357,32'd4731,32'd-711,32'd2622,32'd787,32'd2800,32'd-4553,32'd4870,32'd6118,32'd6528,32'd1669,32'd-4299,32'd-1828,32'd-2988,32'd751,32'd2310,32'd9692,32'd-42,32'd1203,32'd-1398,32'd-4987,32'd2495,32'd9736,32'd3652,32'd2183,32'd2731,32'd-7475,32'd4204,32'd-3134,32'd-132,32'd7280,32'd-2814,32'd-1240,32'd-6992,32'd1067,32'd221,32'd-3244,32'd4321,32'd1442,32'd1322,32'd-1119,32'd-3503};
    Wh[77]='{32'd-3835,32'd4763,32'd-5991,32'd1262,32'd715,32'd2283,32'd-5097,32'd-2758,32'd-3027,32'd2238,32'd9311,32'd-1701,32'd964,32'd103,32'd-1616,32'd-5195,32'd4047,32'd2020,32'd581,32'd1458,32'd2849,32'd898,32'd-167,32'd108,32'd888,32'd-1012,32'd4619,32'd4538,32'd10195,32'd-2817,32'd-2452,32'd2453,32'd807,32'd-485,32'd-2282,32'd-833,32'd-3430,32'd2423,32'd-2404,32'd1066,32'd-404,32'd2709,32'd-2203,32'd653,32'd-2169,32'd-3476,32'd1788,32'd4633,32'd140,32'd279,32'd3371,32'd3710,32'd101,32'd-657,32'd-1401,32'd4094,32'd303,32'd-8232,32'd5019,32'd-6235,32'd1817,32'd-1244,32'd-2832,32'd-1770,32'd1250,32'd-213,32'd-695,32'd-7949,32'd-6059,32'd1342,32'd4411,32'd-7255,32'd-1392,32'd734,32'd-1281,32'd1311,32'd836,32'd-3491,32'd-2973,32'd924,32'd3051,32'd-3459,32'd3828,32'd680,32'd-6826,32'd-1976,32'd-1227,32'd-3769,32'd3122,32'd-3830,32'd5498,32'd110,32'd-1676,32'd-4350,32'd151,32'd-1367,32'd-41,32'd5322,32'd870,32'd5659,32'd6352,32'd-4360,32'd1193,32'd11093,32'd1513,32'd-3625,32'd-5180,32'd-1243,32'd-6372,32'd-3791,32'd-2153,32'd-519,32'd-1160,32'd-1213,32'd-2158,32'd3266,32'd-2480,32'd-6791,32'd4135,32'd4145,32'd2163,32'd3823,32'd6547,32'd-5649,32'd267,32'd4531,32'd-10791,32'd-11416,32'd409,32'd-315,32'd-1771,32'd4528,32'd6049,32'd-6035,32'd2658,32'd2181,32'd7036,32'd3483,32'd2331,32'd-3005,32'd-3564,32'd-3112,32'd886,32'd3266,32'd-135,32'd-350,32'd1375,32'd8686,32'd-192,32'd3369,32'd1707,32'd2113,32'd-1907,32'd4270,32'd-646,32'd-4187,32'd-364,32'd389,32'd1444,32'd9331,32'd-1304,32'd1126,32'd-4006,32'd5805,32'd-1705,32'd-4106,32'd2281,32'd-1658,32'd-1419,32'd1043,32'd5000,32'd1551,32'd3979,32'd-5898,32'd-4284,32'd859,32'd-4174,32'd462,32'd1246,32'd3227,32'd2353,32'd1191,32'd-2202,32'd2319,32'd-1402,32'd3359,32'd-197,32'd1536,32'd-5551,32'd3769,32'd6010,32'd1499,32'd-1525,32'd1702,32'd1284,32'd8383,32'd1291,32'd-1408,32'd-5234,32'd-249,32'd3247,32'd-1589,32'd-1666,32'd5703,32'd-413,32'd660,32'd-2651,32'd-4902,32'd-2648,32'd-1710,32'd2438,32'd-297,32'd-829,32'd3881,32'd-2430,32'd3583,32'd-406,32'd-7675,32'd-3554,32'd-1085,32'd-1263,32'd-825,32'd2785,32'd4431,32'd4902,32'd3706,32'd-1549,32'd-2741,32'd914,32'd3666,32'd5058,32'd-5532,32'd2425,32'd4013,32'd-84,32'd-1232,32'd3686,32'd103,32'd1383,32'd-1068,32'd1617,32'd-1624,32'd356,32'd-3562,32'd-1945,32'd2431,32'd-4511,32'd-3315,32'd3337,32'd-494,32'd-623,32'd2568,32'd784,32'd-5815,32'd-1027,32'd4245,32'd-3776,32'd-5747,32'd-6430,32'd394,32'd1074,32'd2346,32'd-5278,32'd-1071,32'd-3352,32'd1180,32'd2171,32'd-836,32'd-440,32'd-1078,32'd294,32'd-7119,32'd-752,32'd-2939,32'd1794,32'd-870,32'd1700,32'd-2342,32'd2795,32'd488,32'd-2243,32'd4191,32'd2203,32'd1019,32'd4550,32'd2980,32'd-2265,32'd-6625,32'd-2875,32'd-1965,32'd-2690,32'd4645,32'd2775,32'd-9047,32'd-4233,32'd4038,32'd-4953,32'd-2910,32'd-1906,32'd1145,32'd833,32'd-997,32'd-5317,32'd3127,32'd-5644,32'd-5722,32'd1561,32'd-5317,32'd-6479,32'd6645,32'd581,32'd-2070,32'd371,32'd-1447,32'd-3652,32'd2269,32'd-3874,32'd-2001,32'd5332,32'd-547,32'd-549,32'd637,32'd-6777,32'd2408,32'd3662,32'd5053,32'd6376,32'd-1724,32'd2025,32'd2125,32'd3190,32'd-1545,32'd-3508,32'd1994,32'd3747,32'd3237,32'd-496,32'd1940,32'd1424,32'd-2634,32'd657,32'd-5634,32'd-2081,32'd-327,32'd-3305,32'd1000,32'd26,32'd9707,32'd-9296,32'd-41,32'd-7319,32'd-2836,32'd-2570,32'd1966,32'd-944,32'd1485,32'd-2177,32'd-2690,32'd2543,32'd-3205,32'd240,32'd4235,32'd985,32'd2237,32'd-1068,32'd1258,32'd-1210,32'd-2585,32'd3339,32'd369,32'd-564,32'd912,32'd3315,32'd-2829,32'd-2792,32'd-1195,32'd-2346,32'd-993,32'd1436,32'd-6669,32'd-4829,32'd1182,32'd4501,32'd3225,32'd3186,32'd-6005,32'd-10,32'd-3977,32'd1756,32'd-734,32'd232,32'd1966,32'd2648,32'd-597,32'd-2812,32'd-1362,32'd-2243,32'd-508,32'd-4855,32'd1484};
    Wh[78]='{32'd-6972,32'd192,32'd-2509,32'd99,32'd-705,32'd-1370,32'd-2546,32'd-2261,32'd-268,32'd-611,32'd-5053,32'd-6162,32'd-1968,32'd623,32'd1228,32'd1181,32'd-977,32'd-3393,32'd-5053,32'd-6474,32'd-4099,32'd-1622,32'd3496,32'd-4758,32'd-2565,32'd-7231,32'd-740,32'd-1367,32'd-3540,32'd-1643,32'd-6157,32'd1534,32'd-2626,32'd-4528,32'd-2413,32'd953,32'd-2232,32'd-755,32'd-2451,32'd-3366,32'd-2019,32'd542,32'd-290,32'd-4790,32'd6938,32'd2268,32'd-673,32'd-1373,32'd-2590,32'd9716,32'd-607,32'd222,32'd3349,32'd4687,32'd-2459,32'd27,32'd2108,32'd-2447,32'd-1195,32'd802,32'd-5004,32'd-2644,32'd-2687,32'd-182,32'd8198,32'd-6992,32'd2607,32'd-1204,32'd-4707,32'd-6474,32'd-3991,32'd-4357,32'd1447,32'd2121,32'd-6562,32'd-75,32'd-1834,32'd-8466,32'd4228,32'd574,32'd-1065,32'd-3793,32'd-2026,32'd-2362,32'd922,32'd3833,32'd46,32'd-3027,32'd-307,32'd-2399,32'd-2216,32'd-2187,32'd-1943,32'd-5195,32'd-4204,32'd-2200,32'd-1037,32'd-618,32'd-3029,32'd988,32'd2320,32'd5908,32'd3891,32'd1634,32'd6718,32'd1046,32'd5410,32'd7783,32'd1527,32'd-98,32'd-982,32'd4477,32'd10390,32'd4809,32'd-709,32'd-885,32'd-734,32'd-2369,32'd6284,32'd579,32'd2048,32'd5351,32'd-10312,32'd-2255,32'd-1900,32'd-1027,32'd-2739,32'd-3144,32'd-6665,32'd7011,32'd-6835,32'd3811,32'd-3413,32'd-1795,32'd-83,32'd1018,32'd2346,32'd6054,32'd4755,32'd-5981,32'd4423,32'd-2431,32'd-392,32'd-1229,32'd1308,32'd4299,32'd1279,32'd2851,32'd1594,32'd-1025,32'd-4479,32'd-1192,32'd-24687,32'd-431,32'd-5649,32'd5156,32'd-920,32'd-3344,32'd-4748,32'd-246,32'd-9868,32'd-5229,32'd9155,32'd5756,32'd549,32'd7314,32'd-2282,32'd-3664,32'd2186,32'd-2719,32'd-3208,32'd-2966,32'd-1889,32'd-2467,32'd-487,32'd-2246,32'd3000,32'd-2658,32'd-11220,32'd855,32'd-1873,32'd2634,32'd2160,32'd-1483,32'd3452,32'd-3186,32'd-4736,32'd-2749,32'd4877,32'd1550,32'd-7158,32'd-2885,32'd-7778,32'd-1073,32'd2104,32'd931,32'd-1816,32'd-2841,32'd193,32'd-423,32'd570,32'd-3737,32'd-832,32'd-3181,32'd4453,32'd-1043,32'd-2663,32'd-2188,32'd-290,32'd-3256,32'd-3503,32'd3603,32'd-6645,32'd289,32'd-3620,32'd-8920,32'd-3815,32'd2927,32'd-5424,32'd-6445,32'd845,32'd-2666,32'd-8374,32'd1900,32'd-6254,32'd-11777,32'd-3415,32'd1067,32'd-1285,32'd-2141,32'd-3837,32'd-631,32'd-5825,32'd-726,32'd-3454,32'd1490,32'd-3847,32'd1222,32'd-5576,32'd-125,32'd-452,32'd-2932,32'd-758,32'd-3247,32'd-9692,32'd1579,32'd-2440,32'd-1934,32'd-6308,32'd-5751,32'd-5717,32'd-1359,32'd12675,32'd-7612,32'd1458,32'd607,32'd-3593,32'd7812,32'd218,32'd-2476,32'd-4675,32'd-6450,32'd2658,32'd2854,32'd-6982,32'd-8139,32'd-81,32'd-4841,32'd-1098,32'd-4892,32'd667,32'd-7124,32'd-3173,32'd-690,32'd-3583,32'd-4572,32'd833,32'd-4653,32'd-6757,32'd-242,32'd-2193,32'd-1508,32'd-6855,32'd3789,32'd1682,32'd-6606,32'd-4086,32'd-9204,32'd-3386,32'd-9692,32'd5971,32'd-381,32'd-2224,32'd-6455,32'd-4824,32'd-3620,32'd-2500,32'd-3486,32'd699,32'd-7099,32'd-6997,32'd2543,32'd-792,32'd-8325,32'd1597,32'd-1593,32'd-10693,32'd-8613,32'd1823,32'd-884,32'd-5039,32'd-9775,32'd-11503,32'd-4113,32'd-6025,32'd-1407,32'd-9677,32'd-4929,32'd-4592,32'd3483,32'd7158,32'd-3664,32'd-13994,32'd-1700,32'd4899,32'd-2526,32'd-8452,32'd-578,32'd-5327,32'd990,32'd-2685,32'd-2746,32'd-318,32'd235,32'd-5424,32'd1021,32'd-7651,32'd1052,32'd-2287,32'd-4721,32'd3417,32'd1816,32'd-5551,32'd-1871,32'd-8066,32'd-2451,32'd1611,32'd-8251,32'd-4133,32'd6459,32'd-2152,32'd-2464,32'd12548,32'd6918,32'd-5375,32'd-3713,32'd-5776,32'd-2160,32'd-2104,32'd-3398,32'd-13027,32'd-9536,32'd-4895,32'd-1028,32'd-7089,32'd-5454,32'd-4287,32'd-1660,32'd-2153,32'd2020,32'd-6567,32'd-442,32'd1893,32'd-2076,32'd-5014,32'd-6333,32'd-3415,32'd-3198,32'd7875,32'd-3820,32'd-5297,32'd123,32'd3093,32'd-2307,32'd-933,32'd-2827,32'd-9765,32'd-6948,32'd-5668,32'd4482,32'd-838,32'd-3452,32'd2529,32'd1394,32'd-5292,32'd-1263,32'd-1912,32'd-2763,32'd-9355,32'd-4768};
    Wh[79]='{32'd552,32'd424,32'd-745,32'd-1556,32'd-5131,32'd1430,32'd-2437,32'd897,32'd-2902,32'd-1431,32'd4436,32'd2006,32'd5341,32'd-947,32'd-3669,32'd1622,32'd-5117,32'd-2895,32'd-3366,32'd-331,32'd2387,32'd-4841,32'd3442,32'd82,32'd742,32'd-968,32'd-3283,32'd-2163,32'd-3063,32'd-5336,32'd214,32'd1955,32'd-5273,32'd2653,32'd-2183,32'd-5078,32'd-5556,32'd-2093,32'd3239,32'd203,32'd-1573,32'd-5688,32'd2386,32'd-946,32'd4045,32'd-1032,32'd-4291,32'd4055,32'd-2059,32'd-211,32'd4023,32'd-4794,32'd-200,32'd541,32'd-1555,32'd-97,32'd-2998,32'd2966,32'd805,32'd-2069,32'd2531,32'd-512,32'd-547,32'd2368,32'd-1522,32'd3872,32'd-1831,32'd-4990,32'd-2687,32'd-229,32'd-1850,32'd2492,32'd1132,32'd-726,32'd-352,32'd-2347,32'd1160,32'd1540,32'd5712,32'd80,32'd-791,32'd-7456,32'd-433,32'd-1872,32'd-710,32'd818,32'd-1364,32'd1424,32'd-1085,32'd1427,32'd-3129,32'd-5434,32'd3088,32'd1678,32'd6303,32'd-3305,32'd-2753,32'd-2998,32'd-1048,32'd-3066,32'd2707,32'd-945,32'd538,32'd7128,32'd-5336,32'd-12,32'd-1608,32'd1518,32'd-2719,32'd1395,32'd-6445,32'd5292,32'd-3405,32'd1104,32'd514,32'd11,32'd-150,32'd-3166,32'd4816,32'd3615,32'd2971,32'd-1271,32'd7705,32'd-5390,32'd-890,32'd-6337,32'd-3496,32'd-2763,32'd7006,32'd4177,32'd2939,32'd-2893,32'd-1785,32'd-2432,32'd-3220,32'd-2939,32'd-5214,32'd2731,32'd2322,32'd5595,32'd1379,32'd-1417,32'd3247,32'd-4001,32'd-3020,32'd-3305,32'd-1702,32'd687,32'd-3564,32'd-1931,32'd-850,32'd-1342,32'd-1434,32'd-3007,32'd5136,32'd2426,32'd-5751,32'd-2841,32'd3007,32'd-1948,32'd1971,32'd2976,32'd927,32'd-3256,32'd-229,32'd126,32'd-675,32'd-1335,32'd5292,32'd-1181,32'd-6616,32'd-4531,32'd-6250,32'd4990,32'd-133,32'd-4592,32'd140,32'd-1706,32'd-3518,32'd-1723,32'd1151,32'd-558,32'd-867,32'd-279,32'd4516,32'd2231,32'd-2080,32'd-971,32'd899,32'd-2651,32'd-809,32'd-875,32'd-2149,32'd282,32'd2648,32'd-9111,32'd-118,32'd-4851,32'd-5551,32'd205,32'd-4716,32'd2271,32'd740,32'd1855,32'd-1230,32'd370,32'd679,32'd6489,32'd-1190,32'd200,32'd-2424,32'd1646,32'd-2469,32'd-1922,32'd5673,32'd-3229,32'd6264,32'd-5214,32'd3027,32'd-1553,32'd1627,32'd3432,32'd-3549,32'd-376,32'd-4685,32'd2568,32'd-5131,32'd1496,32'd-6005,32'd624,32'd2137,32'd-3291,32'd-484,32'd-3430,32'd-9731,32'd-619,32'd-6459,32'd-364,32'd3881,32'd-1801,32'd1520,32'd2047,32'd-5595,32'd4252,32'd-4450,32'd-1531,32'd-345,32'd4238,32'd1928,32'd324,32'd692,32'd-2966,32'd-749,32'd2954,32'd496,32'd-527,32'd-2286,32'd-2117,32'd-2122,32'd745,32'd-1218,32'd2770,32'd2261,32'd802,32'd1987,32'd2521,32'd-3225,32'd-6083,32'd-1372,32'd-75,32'd-2797,32'd1517,32'd-1262,32'd4006,32'd29,32'd4511,32'd-2951,32'd-605,32'd3483,32'd-1121,32'd4602,32'd-2084,32'd-200,32'd-734,32'd-1490,32'd1621,32'd1519,32'd3251,32'd-829,32'd2697,32'd-2019,32'd-4479,32'd1372,32'd284,32'd-2722,32'd2675,32'd-4091,32'd798,32'd-5024,32'd3647,32'd433,32'd-181,32'd102,32'd967,32'd-3493,32'd-1423,32'd3635,32'd2391,32'd-3720,32'd-154,32'd4245,32'd696,32'd1739,32'd-6411,32'd-713,32'd-4226,32'd3994,32'd-2014,32'd-3781,32'd-3405,32'd-4094,32'd-567,32'd-1895,32'd-1062,32'd-1329,32'd2171,32'd-2976,32'd-4267,32'd3176,32'd-3881,32'd-3205,32'd-2780,32'd-2326,32'd564,32'd-461,32'd110,32'd-2753,32'd-2164,32'd-1046,32'd3801,32'd-2995,32'd3452,32'd-233,32'd-118,32'd186,32'd3381,32'd4240,32'd-2221,32'd613,32'd5283,32'd6401,32'd1389,32'd3981,32'd2358,32'd2656,32'd9213,32'd-1435,32'd633,32'd-4941,32'd713,32'd148,32'd4287,32'd1342,32'd4841,32'd592,32'd4638,32'd-801,32'd-582,32'd-5927,32'd-5336,32'd-148,32'd1149,32'd-3510,32'd-1177,32'd-5483,32'd-1802,32'd994,32'd-1036,32'd-1468,32'd226,32'd1217,32'd4013,32'd6674,32'd3706,32'd-1206,32'd4953,32'd-2183,32'd1704,32'd2509,32'd3166,32'd-2131,32'd420,32'd-673,32'd5415,32'd-236,32'd3339,32'd-986,32'd1065,32'd185,32'd-722};
    Wh[80]='{32'd327,32'd661,32'd-4270,32'd-3264,32'd-709,32'd2039,32'd-677,32'd-2374,32'd1418,32'd-927,32'd-5175,32'd-135,32'd2236,32'd-3266,32'd-6840,32'd195,32'd-5610,32'd-4338,32'd-221,32'd-786,32'd-1949,32'd1152,32'd3845,32'd-1958,32'd-61,32'd-3103,32'd-3420,32'd-949,32'd-2105,32'd71,32'd-2851,32'd1859,32'd498,32'd-560,32'd958,32'd-3044,32'd599,32'd-812,32'd-1078,32'd-2524,32'd2166,32'd-3007,32'd3540,32'd-6157,32'd1712,32'd-268,32'd-2780,32'd-24,32'd-1864,32'd1417,32'd-3056,32'd1331,32'd417,32'd-1409,32'd629,32'd2912,32'd-221,32'd714,32'd-3549,32'd-3208,32'd35,32'd-1613,32'd-176,32'd53,32'd-5327,32'd899,32'd489,32'd-2900,32'd-2585,32'd-885,32'd271,32'd764,32'd399,32'd-4453,32'd-375,32'd-2481,32'd-3381,32'd-3601,32'd1239,32'd81,32'd4350,32'd22,32'd-1359,32'd-3286,32'd-2031,32'd1084,32'd2539,32'd989,32'd2822,32'd284,32'd-3491,32'd-1561,32'd-570,32'd5366,32'd-474,32'd-1077,32'd-1157,32'd-5268,32'd-5761,32'd4057,32'd2658,32'd3286,32'd2807,32'd-7314,32'd-1608,32'd-3740,32'd-4531,32'd-692,32'd4904,32'd1679,32'd-2473,32'd-3657,32'd985,32'd-2192,32'd-4211,32'd265,32'd-1697,32'd-3178,32'd-202,32'd6406,32'd4116,32'd7280,32'd-316,32'd-416,32'd-1254,32'd-253,32'd-7612,32'd-791,32'd1917,32'd2302,32'd1677,32'd93,32'd-1024,32'd3366,32'd1588,32'd3791,32'd-2663,32'd1619,32'd-2480,32'd599,32'd5034,32'd1962,32'd1300,32'd4211,32'd731,32'd-3613,32'd-2075,32'd-6411,32'd1376,32'd-2409,32'd3012,32'd-1356,32'd-293,32'd-4650,32'd459,32'd5737,32'd3522,32'd2761,32'd-2425,32'd-9155,32'd1435,32'd5664,32'd-2033,32'd-4326,32'd207,32'd-2099,32'd-2227,32'd-312,32'd3994,32'd-421,32'd7490,32'd-2069,32'd-1776,32'd163,32'd648,32'd-3854,32'd-2722,32'd-1280,32'd2078,32'd776,32'd-3593,32'd-2927,32'd-1915,32'd-3420,32'd328,32'd2595,32'd-4748,32'd-2863,32'd1435,32'd3674,32'd-1264,32'd5058,32'd-6210,32'd-455,32'd-3188,32'd4511,32'd-89,32'd-3342,32'd-353,32'd1243,32'd44,32'd-930,32'd-1092,32'd-529,32'd-452,32'd1816,32'd-980,32'd-8315,32'd-6772,32'd87,32'd-1538,32'd4553,32'd-2369,32'd1113,32'd38,32'd-4526,32'd1343,32'd-2607,32'd-2128,32'd320,32'd-3269,32'd-1531,32'd7187,32'd2709,32'd1114,32'd-1972,32'd2005,32'd-3320,32'd-1398,32'd-4160,32'd712,32'd-1093,32'd-6396,32'd671,32'd-1359,32'd-1435,32'd-2065,32'd369,32'd871,32'd5180,32'd2758,32'd-2307,32'd2827,32'd-370,32'd4147,32'd614,32'd5756,32'd-227,32'd-2430,32'd-531,32'd-1195,32'd1998,32'd866,32'd320,32'd390,32'd-424,32'd-770,32'd1369,32'd-713,32'd3930,32'd595,32'd-6894,32'd4992,32'd-434,32'd-3627,32'd-150,32'd391,32'd-442,32'd-3962,32'd-1407,32'd480,32'd5991,32'd-909,32'd-2310,32'd-3364,32'd3896,32'd-2687,32'd769,32'd-2322,32'd-3388,32'd1152,32'd2030,32'd1262,32'd-704,32'd-2227,32'd-1395,32'd-1408,32'd-4758,32'd-221,32'd-1276,32'd1647,32'd1445,32'd1972,32'd2288,32'd1632,32'd-6054,32'd730,32'd-3256,32'd-1846,32'd1687,32'd2504,32'd8227,32'd50,32'd-491,32'd-469,32'd-3308,32'd-6396,32'd-2426,32'd-2968,32'd-2100,32'd77,32'd-1683,32'd-1314,32'd-4885,32'd3698,32'd-3857,32'd10781,32'd-7622,32'd-428,32'd-3527,32'd1402,32'd-1201,32'd579,32'd1535,32'd960,32'd673,32'd-4433,32'd-581,32'd1,32'd-3403,32'd-3264,32'd1359,32'd889,32'd-879,32'd-1450,32'd5053,32'd3986,32'd-8535,32'd-2047,32'd3361,32'd2536,32'd-5458,32'd2458,32'd-9028,32'd1600,32'd3701,32'd7036,32'd-2067,32'd-8017,32'd-2536,32'd836,32'd-2041,32'd-5439,32'd-3779,32'd6977,32'd3046,32'd1096,32'd8823,32'd-1693,32'd527,32'd328,32'd-3486,32'd-1599,32'd7963,32'd-1181,32'd5883,32'd-1224,32'd6738,32'd-5239,32'd-994,32'd-4270,32'd-1015,32'd-3381,32'd-3381,32'd-1262,32'd-4233,32'd5292,32'd1024,32'd-3251,32'd-3281,32'd3989,32'd4868,32'd326,32'd-1593,32'd-4101,32'd1705,32'd-1545,32'd-1580,32'd2108,32'd-487,32'd692,32'd136,32'd210,32'd-4672,32'd-1380,32'd-961,32'd7509,32'd-2856,32'd-2756,32'd343};
    Wh[81]='{32'd716,32'd-975,32'd-1533,32'd1987,32'd-2010,32'd-2902,32'd-7338,32'd4003,32'd-3723,32'd-193,32'd-4375,32'd-191,32'd-2612,32'd-1650,32'd-7094,32'd-3383,32'd-10126,32'd-3796,32'd-5517,32'd-284,32'd3293,32'd-4533,32'd-3769,32'd-1552,32'd1101,32'd674,32'd4074,32'd-1591,32'd-5869,32'd219,32'd2252,32'd3837,32'd-380,32'd989,32'd-5322,32'd3310,32'd-1079,32'd-4365,32'd48,32'd785,32'd-3254,32'd8569,32'd914,32'd298,32'd-2008,32'd-1466,32'd1354,32'd1408,32'd3959,32'd-1249,32'd-5351,32'd6821,32'd3300,32'd5219,32'd1585,32'd-9125,32'd-1751,32'd1813,32'd-1026,32'd-24648,32'd-2514,32'd-5039,32'd3317,32'd-6811,32'd-1719,32'd501,32'd-1831,32'd-7456,32'd-4536,32'd-151,32'd-2268,32'd-4082,32'd-1306,32'd-4982,32'd-3410,32'd-4167,32'd-6386,32'd-5122,32'd-3657,32'd-225,32'd592,32'd-487,32'd-3457,32'd9096,32'd-9599,32'd-5415,32'd1697,32'd1282,32'd-6489,32'd-4887,32'd3352,32'd-9423,32'd-5307,32'd3535,32'd2366,32'd-3586,32'd-2797,32'd2348,32'd1204,32'd1816,32'd11005,32'd-3728,32'd216,32'd3950,32'd-3420,32'd-390,32'd-1971,32'd-3515,32'd-8413,32'd12119,32'd2402,32'd-170,32'd823,32'd-6142,32'd-593,32'd735,32'd1949,32'd-10087,32'd-1486,32'd2575,32'd-18,32'd913,32'd-2856,32'd-5463,32'd-8496,32'd-1223,32'd-9702,32'd-7001,32'd4753,32'd-6601,32'd9179,32'd2810,32'd3342,32'd-2277,32'd2445,32'd1135,32'd6616,32'd-628,32'd-6845,32'd5400,32'd6582,32'd-538,32'd-2194,32'd1594,32'd603,32'd2304,32'd-1503,32'd3242,32'd5810,32'd-3266,32'd-3862,32'd728,32'd-6030,32'd2224,32'd-4645,32'd15625,32'd1861,32'd6430,32'd-5883,32'd-11347,32'd10966,32'd-469,32'd625,32'd730,32'd-1805,32'd-7836,32'd-5029,32'd-7192,32'd-2401,32'd-1031,32'd-5468,32'd487,32'd-795,32'd904,32'd-3457,32'd819,32'd-1214,32'd-208,32'd-1420,32'd-310,32'd2152,32'd-122,32'd-4248,32'd2709,32'd3640,32'd240,32'd534,32'd2095,32'd20175,32'd1265,32'd1517,32'd6562,32'd4553,32'd-7109,32'd-1284,32'd-1788,32'd-3913,32'd-3110,32'd-6357,32'd-2741,32'd-2489,32'd-751,32'd6870,32'd-1311,32'd-709,32'd-1128,32'd1821,32'd3442,32'd-708,32'd-7353,32'd643,32'd2484,32'd-1972,32'd3100,32'd-2226,32'd5844,32'd7207,32'd-6381,32'd2783,32'd6860,32'd1756,32'd-3535,32'd-1080,32'd-1026,32'd2685,32'd-621,32'd-531,32'd1263,32'd1821,32'd3356,32'd353,32'd-2785,32'd-3903,32'd2308,32'd-1495,32'd-3901,32'd4956,32'd3696,32'd2338,32'd-3515,32'd1604,32'd4340,32'd-1268,32'd-747,32'd3442,32'd-687,32'd-1252,32'd6489,32'd8315,32'd1479,32'd-833,32'd4699,32'd-2595,32'd-4628,32'd9443,32'd977,32'd4172,32'd-1643,32'd1663,32'd6708,32'd-951,32'd-2333,32'd9980,32'd-3833,32'd-2117,32'd3427,32'd3376,32'd-1561,32'd-2570,32'd2839,32'd-2031,32'd-1636,32'd-4794,32'd1433,32'd-2148,32'd4135,32'd-3715,32'd234,32'd499,32'd3925,32'd-7167,32'd-6772,32'd-1588,32'd3869,32'd4978,32'd3623,32'd-450,32'd-4621,32'd7890,32'd4565,32'd2080,32'd-4924,32'd2570,32'd-1711,32'd-2915,32'd-487,32'd4069,32'd-1884,32'd-503,32'd-964,32'd-6982,32'd5766,32'd2164,32'd-3371,32'd1231,32'd-8740,32'd1022,32'd-1163,32'd-3164,32'd861,32'd2727,32'd-65,32'd-1093,32'd-3898,32'd979,32'd-8588,32'd6596,32'd-2409,32'd-1512,32'd-5170,32'd-444,32'd-7050,32'd-2132,32'd8339,32'd3447,32'd2043,32'd-5800,32'd-4611,32'd-3315,32'd-1685,32'd-4687,32'd5161,32'd6777,32'd732,32'd-571,32'd6997,32'd-4853,32'd-5727,32'd1184,32'd-4431,32'd-1882,32'd-7119,32'd-4741,32'd801,32'd251,32'd-1844,32'd2819,32'd4660,32'd-6645,32'd1726,32'd-2939,32'd-4165,32'd211,32'd497,32'd359,32'd3007,32'd-2604,32'd4804,32'd-7114,32'd-8071,32'd-1442,32'd-14062,32'd1579,32'd-741,32'd682,32'd2543,32'd-1910,32'd2479,32'd-670,32'd-2529,32'd-390,32'd2282,32'd-12050,32'd-3808,32'd-1011,32'd4243,32'd1737,32'd-2758,32'd-3862,32'd-7475,32'd-3283,32'd-2854,32'd-584,32'd-820,32'd2722,32'd-5102,32'd98,32'd-1833,32'd-1018,32'd1145,32'd-2220,32'd7089,32'd-45,32'd-368,32'd-974,32'd-204,32'd771,32'd-4985,32'd-1573,32'd-982};
    Wh[82]='{32'd-112,32'd2634,32'd-2678,32'd1950,32'd-203,32'd-1629,32'd-2639,32'd-912,32'd110,32'd119,32'd-3945,32'd-1226,32'd-2534,32'd-3872,32'd-3378,32'd-645,32'd-864,32'd-1464,32'd-858,32'd2998,32'd-2247,32'd1831,32'd3281,32'd-1820,32'd-2145,32'd-1336,32'd-6303,32'd-180,32'd-3164,32'd540,32'd-568,32'd-9560,32'd709,32'd-412,32'd4111,32'd-2004,32'd3908,32'd-1436,32'd2192,32'd449,32'd-708,32'd120,32'd-944,32'd2261,32'd1857,32'd502,32'd2910,32'd-2463,32'd369,32'd-1477,32'd758,32'd1260,32'd-1550,32'd4775,32'd2355,32'd191,32'd-1944,32'd-2727,32'd-2731,32'd2761,32'd-835,32'd44,32'd731,32'd109,32'd-11259,32'd-2011,32'd-1840,32'd3569,32'd-2196,32'd2049,32'd-1796,32'd875,32'd839,32'd-3469,32'd-3259,32'd3369,32'd3139,32'd-3012,32'd-2172,32'd-7714,32'd-2180,32'd839,32'd844,32'd-4245,32'd668,32'd2602,32'd2337,32'd2587,32'd2500,32'd5766,32'd-386,32'd-661,32'd1793,32'd4489,32'd3400,32'd-611,32'd4799,32'd3293,32'd-942,32'd-194,32'd-1706,32'd-1030,32'd2819,32'd6665,32'd621,32'd3837,32'd-3999,32'd1089,32'd2597,32'd-2142,32'd-4013,32'd-206,32'd-6723,32'd-5361,32'd-1979,32'd-8725,32'd1578,32'd9501,32'd-296,32'd3400,32'd-1252,32'd-4606,32'd1069,32'd1055,32'd-1151,32'd-6162,32'd4655,32'd3791,32'd-3000,32'd2462,32'd-3391,32'd3874,32'd588,32'd-1054,32'd-6059,32'd-774,32'd-5053,32'd3552,32'd-57,32'd-3134,32'd-3291,32'd45,32'd-2856,32'd842,32'd-618,32'd2351,32'd3781,32'd5610,32'd-2785,32'd2795,32'd5058,32'd1307,32'd-674,32'd2871,32'd6430,32'd-279,32'd600,32'd-1364,32'd-1385,32'd-1621,32'd-1030,32'd3293,32'd-2770,32'd-5903,32'd-4985,32'd1696,32'd3366,32'd533,32'd460,32'd2524,32'd6210,32'd93,32'd2048,32'd-2099,32'd-2509,32'd917,32'd-2165,32'd-268,32'd-1535,32'd-4006,32'd-1235,32'd1925,32'd298,32'd-4638,32'd103,32'd-1464,32'd5317,32'd-1016,32'd-221,32'd-1150,32'd-2121,32'd-345,32'd341,32'd-2880,32'd-307,32'd96,32'd-3142,32'd-1556,32'd2109,32'd747,32'd1275,32'd2130,32'd-48,32'd-1065,32'd3984,32'd-1227,32'd3369,32'd-2739,32'd-1834,32'd1557,32'd4785,32'd3249,32'd-3547,32'd645,32'd-1068,32'd1223,32'd3068,32'd8891,32'd-276,32'd2092,32'd-2897,32'd-4035,32'd-3142,32'd-3215,32'd-1486,32'd-4091,32'd-3137,32'd186,32'd-629,32'd1925,32'd516,32'd-1348,32'd-3415,32'd2166,32'd1209,32'd-5883,32'd-3039,32'd-935,32'd-3144,32'd1796,32'd5747,32'd-790,32'd2091,32'd-1855,32'd2600,32'd2709,32'd1806,32'd-950,32'd-4675,32'd3137,32'd2932,32'd3161,32'd2384,32'd-2954,32'd663,32'd2266,32'd-3386,32'd4296,32'd-791,32'd2934,32'd1518,32'd6279,32'd-959,32'd1003,32'd-121,32'd-1518,32'd1156,32'd461,32'd-1030,32'd1883,32'd1824,32'd-190,32'd-1939,32'd-1158,32'd1466,32'd-4819,32'd10029,32'd-3786,32'd34,32'd5805,32'd-1834,32'd678,32'd5327,32'd-1339,32'd-395,32'd3457,32'd1166,32'd1154,32'd-3813,32'd175,32'd2919,32'd1828,32'd-2416,32'd275,32'd-228,32'd-2202,32'd597,32'd1329,32'd-2504,32'd-634,32'd3171,32'd-425,32'd1260,32'd1331,32'd-1387,32'd5708,32'd-2285,32'd604,32'd-848,32'd2651,32'd-1282,32'd711,32'd-4458,32'd-3642,32'd1790,32'd5615,32'd-5600,32'd-1328,32'd3234,32'd-1306,32'd-3198,32'd-5004,32'd-2946,32'd-2565,32'd1929,32'd-949,32'd-1423,32'd5219,32'd-4365,32'd-1632,32'd-1822,32'd-2019,32'd2249,32'd3671,32'd3903,32'd-7661,32'd-3576,32'd-762,32'd-3403,32'd-903,32'd-262,32'd2761,32'd939,32'd-3574,32'd2585,32'd-334,32'd-6416,32'd-3007,32'd-2427,32'd134,32'd-517,32'd3835,32'd5161,32'd6450,32'd-1018,32'd-3728,32'd-286,32'd4985,32'd3298,32'd4919,32'd2482,32'd-1654,32'd1855,32'd1246,32'd-3098,32'd3691,32'd-1966,32'd-4108,32'd2199,32'd2973,32'd-1773,32'd3864,32'd8071,32'd3308,32'd2590,32'd3149,32'd-4304,32'd-958,32'd2060,32'd2900,32'd-2296,32'd-5371,32'd5205,32'd-1034,32'd2352,32'd-1028,32'd4047,32'd3698,32'd4724,32'd3203,32'd4494,32'd-1663,32'd1871,32'd-6059,32'd-2504,32'd3535,32'd2399,32'd-4448,32'd-3039,32'd6186};
    Wh[83]='{32'd3012,32'd5683,32'd2176,32'd-2802,32'd1644,32'd697,32'd10468,32'd4553,32'd461,32'd-78,32'd5273,32'd-3449,32'd1542,32'd-7524,32'd138,32'd3447,32'd-4177,32'd3117,32'd2238,32'd-2429,32'd2034,32'd-1632,32'd1857,32'd858,32'd-1976,32'd-2277,32'd-1921,32'd1235,32'd2032,32'd1831,32'd5712,32'd-3098,32'd11132,32'd3984,32'd2054,32'd-1152,32'd2524,32'd2927,32'd3200,32'd-88,32'd4318,32'd-1047,32'd-157,32'd-2059,32'd108,32'd1228,32'd-2895,32'd-6533,32'd786,32'd-106,32'd2441,32'd-1007,32'd3833,32'd-1030,32'd919,32'd-422,32'd901,32'd-457,32'd427,32'd-1984,32'd223,32'd2502,32'd2438,32'd6689,32'd1111,32'd602,32'd7436,32'd5083,32'd2775,32'd-3710,32'd507,32'd-8300,32'd2471,32'd21,32'd2299,32'd524,32'd8437,32'd10205,32'd3469,32'd1988,32'd-4096,32'd-2014,32'd10283,32'd-6191,32'd7241,32'd282,32'd-2026,32'd-2062,32'd1779,32'd4252,32'd-3181,32'd-605,32'd3632,32'd-3332,32'd963,32'd-5971,32'd1507,32'd-8637,32'd495,32'd1722,32'd-14814,32'd416,32'd-2132,32'd2386,32'd7895,32'd-342,32'd1678,32'd11093,32'd12929,32'd5615,32'd-651,32'd16132,32'd6689,32'd2824,32'd-2087,32'd1893,32'd232,32'd1223,32'd-6088,32'd-6333,32'd5639,32'd-7363,32'd546,32'd-340,32'd9487,32'd-8237,32'd16748,32'd2401,32'd1174,32'd-335,32'd-404,32'd3000,32'd-2239,32'd706,32'd-3769,32'd-1161,32'd2944,32'd3857,32'd1802,32'd2512,32'd-9047,32'd-4645,32'd567,32'd1490,32'd1617,32'd-1104,32'd2027,32'd-2403,32'd11308,32'd2332,32'd-5688,32'd-3481,32'd3278,32'd2766,32'd7729,32'd-1774,32'd3193,32'd-2313,32'd3696,32'd8940,32'd-3835,32'd2486,32'd-4770,32'd5771,32'd3378,32'd6313,32'd-1932,32'd3874,32'd-2915,32'd-3884,32'd547,32'd-1333,32'd-2005,32'd5351,32'd2165,32'd772,32'd2445,32'd1641,32'd-1440,32'd-3627,32'd63,32'd-642,32'd-4353,32'd-4645,32'd-1176,32'd6645,32'd3393,32'd-4672,32'd-9033,32'd8334,32'd-6123,32'd-5541,32'd-3208,32'd673,32'd6040,32'd-8310,32'd-4772,32'd6748,32'd8618,32'd727,32'd1199,32'd7055,32'd-3408,32'd3364,32'd5185,32'd-2065,32'd323,32'd-3581,32'd-411,32'd10605,32'd-1518,32'd1397,32'd-8325,32'd255,32'd-5410,32'd-4643,32'd-474,32'd3063,32'd-6840,32'd-255,32'd5424,32'd168,32'd255,32'd-1610,32'd-5000,32'd-1744,32'd-707,32'd-3039,32'd-1864,32'd-711,32'd-6,32'd-1591,32'd1381,32'd-2089,32'd-3974,32'd-4328,32'd-786,32'd-5019,32'd1976,32'd4250,32'd-3134,32'd203,32'd-1138,32'd9702,32'd-2459,32'd-1909,32'd614,32'd-584,32'd499,32'd405,32'd-925,32'd3449,32'd2382,32'd-386,32'd-5708,32'd650,32'd-786,32'd-1523,32'd-236,32'd-260,32'd2829,32'd6811,32'd-6416,32'd-4379,32'd2778,32'd4406,32'd4206,32'd3618,32'd-1855,32'd-1982,32'd2413,32'd875,32'd4936,32'd2912,32'd-640,32'd4433,32'd572,32'd-381,32'd-298,32'd-1120,32'd9462,32'd3483,32'd2829,32'd-3139,32'd-2971,32'd3933,32'd-3645,32'd9399,32'd-3955,32'd-8027,32'd-3215,32'd-1419,32'd3188,32'd4377,32'd3083,32'd2636,32'd974,32'd374,32'd-696,32'd-5917,32'd6728,32'd-7646,32'd2578,32'd2707,32'd-2612,32'd4040,32'd7666,32'd3259,32'd2763,32'd-2775,32'd1282,32'd453,32'd-2954,32'd10419,32'd-2476,32'd4873,32'd2536,32'd2109,32'd2229,32'd4602,32'd9921,32'd3581,32'd1429,32'd-3525,32'd-260,32'd-4638,32'd4475,32'd770,32'd-964,32'd-394,32'd2443,32'd4355,32'd-3237,32'd-807,32'd899,32'd-4904,32'd4086,32'd-691,32'd-4685,32'd-4895,32'd2028,32'd3454,32'd-1636,32'd-5664,32'd-1590,32'd-8154,32'd-5903,32'd6083,32'd-287,32'd961,32'd398,32'd3562,32'd-1407,32'd-7646,32'd-11328,32'd-3176,32'd4394,32'd-394,32'd3876,32'd2595,32'd-3493,32'd3920,32'd-886,32'd2312,32'd3483,32'd-3095,32'd260,32'd-2983,32'd-2004,32'd-8417,32'd5258,32'd-1679,32'd3676,32'd6958,32'd839,32'd-503,32'd-4294,32'd4255,32'd4387,32'd4279,32'd-1147,32'd1754,32'd-1671,32'd-4089,32'd4245,32'd4326,32'd-2978,32'd5986,32'd-228,32'd1070,32'd1486,32'd-4580,32'd8427,32'd1175,32'd6015,32'd999,32'd1921,32'd13457,32'd-646,32'd-736};
    Wh[84]='{32'd2399,32'd-9931,32'd-1389,32'd-409,32'd-3188,32'd2797,32'd1556,32'd4177,32'd-1322,32'd-44,32'd-148,32'd-239,32'd987,32'd407,32'd5488,32'd-4260,32'd-3669,32'd2230,32'd-1452,32'd944,32'd-32,32'd-1547,32'd1750,32'd-2536,32'd-1771,32'd-1041,32'd-920,32'd-3352,32'd49,32'd-6982,32'd-1975,32'd-2296,32'd-7753,32'd628,32'd-629,32'd-3745,32'd1376,32'd-2592,32'd1011,32'd-6064,32'd908,32'd-543,32'd-1680,32'd-1351,32'd-3862,32'd-38,32'd-1068,32'd-3710,32'd-1350,32'd322,32'd-497,32'd4370,32'd2479,32'd490,32'd4165,32'd-1697,32'd-2934,32'd2607,32'd-157,32'd-9697,32'd6640,32'd-2219,32'd234,32'd-696,32'd-528,32'd-704,32'd6923,32'd-4772,32'd-1181,32'd4255,32'd2451,32'd-788,32'd-7,32'd-2861,32'd-4189,32'd-4750,32'd-2360,32'd3237,32'd3303,32'd-566,32'd-2792,32'd-9443,32'd2604,32'd-2653,32'd2861,32'd-1368,32'd-2438,32'd-96,32'd-147,32'd-247,32'd-6503,32'd-10556,32'd-5576,32'd1866,32'd-1944,32'd695,32'd-3332,32'd-100,32'd-1898,32'd-3513,32'd-3391,32'd-1551,32'd-1695,32'd-5952,32'd-1577,32'd587,32'd-3789,32'd7221,32'd3750,32'd-5883,32'd-4916,32'd5844,32'd6357,32'd-1818,32'd-4970,32'd-4301,32'd1452,32'd5078,32'd-3869,32'd908,32'd3571,32'd-1373,32'd1890,32'd662,32'd-648,32'd-3100,32'd545,32'd1826,32'd-3508,32'd7504,32'd-3012,32'd4875,32'd1702,32'd3676,32'd7338,32'd-3952,32'd2027,32'd2548,32'd3608,32'd1197,32'd-1112,32'd-498,32'd4926,32'd2526,32'd-3269,32'd-37,32'd-3710,32'd8349,32'd-6035,32'd936,32'd242,32'd-2299,32'd4636,32'd-4504,32'd1345,32'd5371,32'd-3068,32'd-4477,32'd4353,32'd-3107,32'd-2868,32'd-1529,32'd2841,32'd1047,32'd-5117,32'd-268,32'd-5375,32'd1632,32'd-1667,32'd4387,32'd-7128,32'd-2521,32'd-1716,32'd452,32'd-1574,32'd-1909,32'd-2204,32'd4184,32'd2744,32'd-2036,32'd-1038,32'd-9257,32'd-1342,32'd-419,32'd1149,32'd329,32'd350,32'd-1173,32'd-1989,32'd2043,32'd1093,32'd3588,32'd-2021,32'd2009,32'd2399,32'd-392,32'd1433,32'd-6259,32'd-3056,32'd-989,32'd-1183,32'd-1566,32'd1672,32'd3381,32'd-426,32'd1420,32'd-854,32'd-2141,32'd-2927,32'd902,32'd1154,32'd-2453,32'd-6557,32'd-3618,32'd3530,32'd2978,32'd8134,32'd2243,32'd-872,32'd-1118,32'd1815,32'd-7758,32'd-2937,32'd-989,32'd-1750,32'd-4645,32'd-9877,32'd-2005,32'd-2346,32'd496,32'd463,32'd-2092,32'd-1072,32'd-969,32'd-12177,32'd-719,32'd1627,32'd-1912,32'd1168,32'd-934,32'd-28,32'd3559,32'd-3601,32'd-2971,32'd-5356,32'd1660,32'd-3859,32'd8378,32'd-2036,32'd-5561,32'd4558,32'd-1624,32'd1001,32'd696,32'd-1376,32'd-1090,32'd-3276,32'd3762,32'd1495,32'd-3984,32'd6386,32'd2259,32'd-4921,32'd-1005,32'd4077,32'd-1405,32'd1788,32'd-2941,32'd-1268,32'd3864,32'd4506,32'd-5400,32'd-5517,32'd-77,32'd-2902,32'd3105,32'd-1224,32'd-1250,32'd-5795,32'd-1666,32'd-2607,32'd494,32'd1710,32'd3029,32'd800,32'd2792,32'd2033,32'd1668,32'd2749,32'd-1144,32'd-2590,32'd941,32'd-2398,32'd5024,32'd523,32'd3745,32'd4233,32'd-735,32'd-2727,32'd1737,32'd-3308,32'd2629,32'd-1490,32'd-887,32'd-1100,32'd-4829,32'd3991,32'd2460,32'd-18,32'd1762,32'd4160,32'd3557,32'd-42,32'd4682,32'd1481,32'd3208,32'd-5371,32'd3898,32'd-4426,32'd1582,32'd-2178,32'd-3193,32'd1077,32'd-2170,32'd-1676,32'd-765,32'd-6171,32'd-5244,32'd1514,32'd-1885,32'd-3652,32'd57,32'd5585,32'd1363,32'd1074,32'd-7241,32'd-928,32'd-219,32'd4565,32'd-1535,32'd5424,32'd1416,32'd-3530,32'd2797,32'd-4042,32'd-5239,32'd-1556,32'd752,32'd-3674,32'd-289,32'd-3518,32'd728,32'd2724,32'd2768,32'd-2514,32'd-2434,32'd-5737,32'd-8867,32'd-3894,32'd-1519,32'd907,32'd-1600,32'd358,32'd-5693,32'd-1575,32'd-4975,32'd6591,32'd2453,32'd-3435,32'd-138,32'd-2294,32'd581,32'd-4768,32'd2293,32'd-2639,32'd-621,32'd1649,32'd-703,32'd2055,32'd3498,32'd-257,32'd2070,32'd3957,32'd4902,32'd-5112,32'd-4858,32'd-1801,32'd-1784,32'd-878,32'd1372,32'd-248,32'd7055,32'd1095,32'd-567,32'd-2844,32'd-7001,32'd4916,32'd-1489,32'd-4108,32'd-945};
    Wh[85]='{32'd1375,32'd-6132,32'd-1386,32'd733,32'd2893,32'd505,32'd-3200,32'd-3154,32'd-2028,32'd334,32'd10996,32'd-1666,32'd1903,32'd4636,32'd-83,32'd-6,32'd173,32'd1171,32'd2249,32'd-148,32'd2763,32'd-1296,32'd-4689,32'd3662,32'd1804,32'd-6479,32'd6826,32'd4592,32'd2442,32'd-414,32'd1501,32'd3391,32'd1811,32'd1203,32'd235,32'd-1007,32'd-110,32'd925,32'd-1237,32'd2043,32'd-3056,32'd4042,32'd2318,32'd-4462,32'd3588,32'd4279,32'd-4902,32'd-576,32'd-4536,32'd1457,32'd-337,32'd6391,32'd1807,32'd-3293,32'd-97,32'd-2900,32'd3129,32'd2142,32'd-3684,32'd-544,32'd-1700,32'd398,32'd4421,32'd-277,32'd4465,32'd3920,32'd1099,32'd631,32'd-5634,32'd-761,32'd-5029,32'd1386,32'd-2541,32'd-120,32'd3317,32'd7285,32'd10117,32'd-2108,32'd3603,32'd-1689,32'd-1801,32'd-5766,32'd3591,32'd2983,32'd-1200,32'd4855,32'd47,32'd-891,32'd2396,32'd317,32'd1557,32'd6694,32'd575,32'd7592,32'd1155,32'd-1295,32'd390,32'd-327,32'd-1838,32'd-4675,32'd8530,32'd-4221,32'd1744,32'd-12695,32'd-4458,32'd-459,32'd2034,32'd-1898,32'd-2622,32'd1030,32'd-1870,32'd14355,32'd6635,32'd82,32'd2360,32'd-3562,32'd1654,32'd15,32'd3161,32'd2092,32'd-6196,32'd1887,32'd4697,32'd2819,32'd6601,32'd-2651,32'd-1149,32'd-4514,32'd9487,32'd4301,32'd39,32'd728,32'd2504,32'd-5952,32'd9804,32'd2568,32'd8701,32'd440,32'd3935,32'd2695,32'd-2834,32'd5053,32'd2736,32'd-4641,32'd1175,32'd-1748,32'd-4140,32'd2641,32'd-1011,32'd1129,32'd-4555,32'd-5117,32'd-4663,32'd6796,32'd7397,32'd2006,32'd-1457,32'd238,32'd-3237,32'd-600,32'd140,32'd-283,32'd1984,32'd7338,32'd2363,32'd-107,32'd-5097,32'd235,32'd4633,32'd-429,32'd-3125,32'd7304,32'd-7895,32'd1192,32'd-6767,32'd-2648,32'd5849,32'd1938,32'd509,32'd5327,32'd6318,32'd131,32'd-9809,32'd3601,32'd1912,32'd-550,32'd-4306,32'd8627,32'd-8515,32'd-930,32'd4162,32'd7729,32'd-5366,32'd2293,32'd6430,32'd-10458,32'd3369,32'd1200,32'd5156,32'd437,32'd-4501,32'd-2900,32'd-1224,32'd-7622,32'd-188,32'd-744,32'd303,32'd-4887,32'd14003,32'd-2883,32'd-6381,32'd3596,32'd220,32'd6743,32'd-6298,32'd-1340,32'd7158,32'd-343,32'd4504,32'd8041,32'd-1118,32'd6660,32'd9511,32'd6479,32'd861,32'd3281,32'd-848,32'd-2954,32'd4062,32'd-4929,32'd1229,32'd-4692,32'd2687,32'd-7592,32'd1783,32'd1140,32'd141,32'd-379,32'd440,32'd2817,32'd5410,32'd858,32'd-2382,32'd-96,32'd1549,32'd827,32'd-59,32'd-50,32'd-1207,32'd1367,32'd-3505,32'd-2239,32'd-3747,32'd-1739,32'd-2220,32'd-1406,32'd-6733,32'd127,32'd2050,32'd-6586,32'd3454,32'd-476,32'd-5532,32'd-3806,32'd1424,32'd-651,32'd-3940,32'd-1513,32'd-2556,32'd-1047,32'd-629,32'd-2695,32'd3735,32'd-775,32'd-584,32'd437,32'd-2467,32'd-3461,32'd-2077,32'd2053,32'd4067,32'd-902,32'd-4506,32'd-8232,32'd-1697,32'd-1511,32'd2607,32'd-6401,32'd15312,32'd-908,32'd5751,32'd8198,32'd-957,32'd624,32'd2442,32'd-5649,32'd-632,32'd3701,32'd-2766,32'd-1070,32'd-615,32'd1572,32'd-719,32'd5800,32'd3249,32'd4089,32'd-4687,32'd-2207,32'd426,32'd-5029,32'd9291,32'd229,32'd-3764,32'd1339,32'd-2556,32'd-3088,32'd1644,32'd5888,32'd1784,32'd3981,32'd4514,32'd6586,32'd7065,32'd-2583,32'd1895,32'd1185,32'd-2360,32'd-485,32'd-853,32'd631,32'd100,32'd-1462,32'd-690,32'd-2612,32'd1563,32'd6069,32'd-553,32'd-2609,32'd5766,32'd138,32'd672,32'd-4121,32'd6,32'd-670,32'd2648,32'd3454,32'd-404,32'd-3959,32'd-4599,32'd1078,32'd-853,32'd-3266,32'd1304,32'd-1176,32'd4401,32'd-529,32'd2832,32'd-2414,32'd-110,32'd575,32'd-5991,32'd776,32'd-1160,32'd1300,32'd-4257,32'd994,32'd1668,32'd-692,32'd1435,32'd880,32'd39,32'd-4702,32'd431,32'd8647,32'd1159,32'd-2445,32'd3986,32'd4831,32'd982,32'd-7392,32'd14638,32'd-287,32'd402,32'd9682,32'd-3361,32'd3635,32'd2000,32'd-3942,32'd-151,32'd-6000,32'd-1270,32'd1611,32'd-66,32'd-8002,32'd-491,32'd-714,32'd3256,32'd-7651,32'd-271,32'd-4079};
    Wh[86]='{32'd-1676,32'd323,32'd-372,32'd3269,32'd1354,32'd-699,32'd-3623,32'd-2602,32'd3518,32'd1628,32'd3620,32'd1069,32'd1308,32'd-4399,32'd-5434,32'd1981,32'd-163,32'd-609,32'd-4685,32'd2780,32'd-1608,32'd1560,32'd6860,32'd-784,32'd-1556,32'd-4511,32'd776,32'd-428,32'd-297,32'd2015,32'd1069,32'd1275,32'd-697,32'd250,32'd-12,32'd-458,32'd-1535,32'd-166,32'd-1086,32'd342,32'd2729,32'd1931,32'd-2355,32'd-1081,32'd222,32'd-3225,32'd1503,32'd3974,32'd-33,32'd-2335,32'd-3879,32'd1423,32'd-2851,32'd-1205,32'd-2653,32'd-4812,32'd3171,32'd-3889,32'd3449,32'd2229,32'd3137,32'd3710,32'd-4003,32'd-6562,32'd-8461,32'd4147,32'd258,32'd4394,32'd2454,32'd-1768,32'd668,32'd2036,32'd3330,32'd7,32'd1002,32'd2338,32'd5727,32'd5249,32'd83,32'd-1015,32'd-2724,32'd2432,32'd-7084,32'd458,32'd601,32'd-4094,32'd-703,32'd-2761,32'd-503,32'd2709,32'd1434,32'd-886,32'd2458,32'd-1500,32'd2697,32'd1975,32'd872,32'd-667,32'd2922,32'd299,32'd-3867,32'd-2291,32'd2934,32'd1431,32'd-894,32'd-1267,32'd87,32'd-792,32'd1334,32'd-1278,32'd1979,32'd2174,32'd-5166,32'd-390,32'd624,32'd-200,32'd-1658,32'd1690,32'd5288,32'd185,32'd-1425,32'd-2868,32'd7988,32'd-592,32'd3291,32'd-220,32'd4257,32'd-388,32'd1633,32'd-4211,32'd7260,32'd-535,32'd1384,32'd-2702,32'd-3464,32'd749,32'd-1151,32'd-4550,32'd-3688,32'd246,32'd284,32'd-1768,32'd-2998,32'd-7285,32'd-1379,32'd-1337,32'd-688,32'd-370,32'd2978,32'd-5991,32'd1666,32'd-3039,32'd-3308,32'd2150,32'd876,32'd-294,32'd-1971,32'd1923,32'd5073,32'd-5175,32'd2722,32'd3251,32'd-1462,32'd-3278,32'd2028,32'd-4113,32'd2807,32'd4492,32'd1341,32'd-139,32'd3010,32'd3454,32'd1882,32'd969,32'd-84,32'd877,32'd-792,32'd2249,32'd-2117,32'd-418,32'd-551,32'd-579,32'd5278,32'd2951,32'd114,32'd7211,32'd2279,32'd2968,32'd1052,32'd-921,32'd4343,32'd2258,32'd-3129,32'd-1556,32'd-5781,32'd696,32'd-1751,32'd982,32'd679,32'd-3889,32'd-627,32'd2558,32'd-778,32'd2880,32'd2135,32'd-1719,32'd1246,32'd2119,32'd-442,32'd-676,32'd1569,32'd3740,32'd5742,32'd2702,32'd2210,32'd2460,32'd2189,32'd3071,32'd4155,32'd-2291,32'd-673,32'd210,32'd-3579,32'd762,32'd-1188,32'd5737,32'd1909,32'd1427,32'd3608,32'd4038,32'd1840,32'd910,32'd-304,32'd2183,32'd5615,32'd-2156,32'd3430,32'd2048,32'd5000,32'd1211,32'd2003,32'd-6376,32'd82,32'd-3352,32'd-822,32'd-266,32'd3020,32'd-8100,32'd-2362,32'd-164,32'd-2386,32'd620,32'd-2988,32'd3994,32'd-3117,32'd4572,32'd-957,32'd-1026,32'd52,32'd3442,32'd-2661,32'd-58,32'd5458,32'd-1208,32'd584,32'd784,32'd-389,32'd-2531,32'd29,32'd-1424,32'd-2362,32'd4536,32'd-371,32'd-2138,32'd-2529,32'd1785,32'd1871,32'd3256,32'd676,32'd-643,32'd-725,32'd-1011,32'd-141,32'd1994,32'd-449,32'd1155,32'd1951,32'd-11,32'd4147,32'd2270,32'd2749,32'd2785,32'd-4865,32'd-1978,32'd600,32'd-1984,32'd-2631,32'd3339,32'd6596,32'd3200,32'd-179,32'd-712,32'd512,32'd2856,32'd1763,32'd706,32'd-3515,32'd-2196,32'd1340,32'd-1718,32'd554,32'd4016,32'd2707,32'd-5878,32'd1340,32'd-1406,32'd-5146,32'd-797,32'd4072,32'd-3022,32'd-4079,32'd3532,32'd1901,32'd-56,32'd-916,32'd1718,32'd4653,32'd910,32'd296,32'd1735,32'd-102,32'd2575,32'd-5161,32'd480,32'd3286,32'd508,32'd2763,32'd-1940,32'd-3920,32'd377,32'd766,32'd-3339,32'd-3195,32'd-2335,32'd-3266,32'd312,32'd-3110,32'd419,32'd3129,32'd1048,32'd-2142,32'd-4055,32'd-1458,32'd-451,32'd-1826,32'd-6430,32'd-1085,32'd4340,32'd2517,32'd-3884,32'd-3100,32'd-293,32'd1386,32'd-1960,32'd-456,32'd-1943,32'd-770,32'd2812,32'd-3161,32'd1759,32'd961,32'd2639,32'd3845,32'd-3713,32'd-531,32'd717,32'd-3928,32'd-485,32'd5146,32'd6259,32'd-1474,32'd-4960,32'd1607,32'd-8432,32'd-525,32'd-1304,32'd4213,32'd878,32'd-861,32'd-1877,32'd1025,32'd590,32'd-5854,32'd-2653,32'd668,32'd2700,32'd-2973,32'd-4133,32'd2780,32'd3559};
    Wh[87]='{32'd1759,32'd967,32'd1506,32'd-2121,32'd-711,32'd4704,32'd-4001,32'd-3125,32'd1734,32'd-2788,32'd798,32'd-363,32'd-2093,32'd1651,32'd3420,32'd911,32'd-4794,32'd-5664,32'd2258,32'd-336,32'd1018,32'd559,32'd-5708,32'd-823,32'd-451,32'd7133,32'd3388,32'd614,32'd4267,32'd81,32'd-622,32'd1060,32'd-1571,32'd-899,32'd4299,32'd-1584,32'd2536,32'd1397,32'd-482,32'd-3496,32'd852,32'd-581,32'd4919,32'd-3212,32'd4873,32'd3032,32'd563,32'd68,32'd2937,32'd-836,32'd1804,32'd-3227,32'd-4313,32'd-698,32'd-723,32'd-1998,32'd-2067,32'd316,32'd-691,32'd7617,32'd-5644,32'd582,32'd-3334,32'd531,32'd3762,32'd4667,32'd3842,32'd-576,32'd-1184,32'd877,32'd-2695,32'd-4067,32'd-230,32'd5869,32'd-545,32'd-3786,32'd163,32'd5297,32'd3137,32'd286,32'd-634,32'd-4560,32'd6352,32'd-1712,32'd983,32'd-381,32'd-1296,32'd-2141,32'd-1335,32'd2785,32'd6054,32'd-756,32'd-1,32'd-3059,32'd-2446,32'd-2152,32'd-1578,32'd3068,32'd-2746,32'd1233,32'd3554,32'd1738,32'd494,32'd-288,32'd469,32'd-4665,32'd-6025,32'd-657,32'd-4409,32'd-3500,32'd2469,32'd-2634,32'd1229,32'd-2800,32'd2514,32'd4580,32'd2009,32'd-1779,32'd-5131,32'd444,32'd911,32'd8037,32'd7553,32'd-1063,32'd-5493,32'd-6215,32'd3303,32'd-789,32'd-992,32'd1578,32'd910,32'd834,32'd2215,32'd-1690,32'd1711,32'd4440,32'd419,32'd2731,32'd-1818,32'd1662,32'd-1958,32'd1560,32'd310,32'd1528,32'd163,32'd3686,32'd6040,32'd-3491,32'd-2030,32'd-1083,32'd2229,32'd1872,32'd2390,32'd5415,32'd2253,32'd1319,32'd1519,32'd-3513,32'd-2265,32'd10947,32'd-3784,32'd6367,32'd-1352,32'd-2465,32'd2556,32'd-2191,32'd1301,32'd-2407,32'd-867,32'd6684,32'd3305,32'd7475,32'd-2415,32'd-3322,32'd3803,32'd-2124,32'd2023,32'd-240,32'd-2253,32'd-1662,32'd-2343,32'd-1513,32'd-3005,32'd-426,32'd5209,32'd2890,32'd1423,32'd-3369,32'd2700,32'd231,32'd2683,32'd-1862,32'd664,32'd-2218,32'd-2731,32'd4929,32'd391,32'd289,32'd-5961,32'd1687,32'd3085,32'd-1027,32'd-1320,32'd-3046,32'd-938,32'd-966,32'd528,32'd1939,32'd548,32'd-345,32'd-1479,32'd-695,32'd-1398,32'd-3967,32'd-480,32'd-5493,32'd1625,32'd5312,32'd1336,32'd503,32'd650,32'd-1754,32'd-586,32'd1118,32'd-4775,32'd-1302,32'd2048,32'd95,32'd486,32'd1572,32'd4072,32'd379,32'd3635,32'd485,32'd-3688,32'd1347,32'd-2810,32'd3015,32'd-4226,32'd-908,32'd-3627,32'd-3623,32'd2196,32'd3969,32'd-2237,32'd-1500,32'd5781,32'd1602,32'd-33,32'd2042,32'd-1911,32'd-917,32'd-1422,32'd-7426,32'd-508,32'd-3354,32'd-2396,32'd-6850,32'd-597,32'd-4338,32'd7949,32'd-1857,32'd4157,32'd2165,32'd-218,32'd-148,32'd189,32'd-65,32'd2385,32'd1151,32'd-1419,32'd-939,32'd3959,32'd-1685,32'd4707,32'd2619,32'd4628,32'd-258,32'd2890,32'd6064,32'd281,32'd2445,32'd4436,32'd-2822,32'd3205,32'd3618,32'd-848,32'd4582,32'd3342,32'd-3828,32'd-2449,32'd-1802,32'd131,32'd-1868,32'd1716,32'd-183,32'd3359,32'd2644,32'd-3657,32'd2746,32'd186,32'd5786,32'd102,32'd4409,32'd-1258,32'd4245,32'd3405,32'd-4396,32'd510,32'd3676,32'd-2839,32'd1779,32'd-4465,32'd1660,32'd4760,32'd-2239,32'd5839,32'd178,32'd6083,32'd-2622,32'd-2158,32'd-890,32'd-1994,32'd-1894,32'd-5576,32'd3217,32'd-6113,32'd-1781,32'd5327,32'd3225,32'd3315,32'd3732,32'd4414,32'd2998,32'd-3977,32'd128,32'd-422,32'd-1264,32'd1062,32'd-2739,32'd1594,32'd6162,32'd1730,32'd-719,32'd5141,32'd-4802,32'd5112,32'd-369,32'd5937,32'd-3356,32'd6816,32'd2805,32'd-2841,32'd1927,32'd-4138,32'd-2575,32'd3061,32'd5498,32'd10214,32'd2939,32'd-407,32'd-487,32'd-211,32'd-4868,32'd-205,32'd672,32'd-563,32'd4572,32'd-1928,32'd-1254,32'd-3776,32'd3508,32'd430,32'd3090,32'd1018,32'd2924,32'd-246,32'd-2260,32'd2401,32'd-1862,32'd1968,32'd1978,32'd2949,32'd1911,32'd-3901,32'd4958,32'd-176,32'd2158,32'd-3813,32'd-2468,32'd1268,32'd110,32'd-7919,32'd-5224,32'd-4682,32'd92,32'd-1018,32'd114,32'd-1534,32'd-97};
    Wh[88]='{32'd2714,32'd353,32'd152,32'd-3442,32'd466,32'd2019,32'd1462,32'd-1127,32'd-2683,32'd-1217,32'd1236,32'd1879,32'd-7158,32'd1915,32'd2702,32'd847,32'd1658,32'd1121,32'd-346,32'd1049,32'd-587,32'd1889,32'd-2462,32'd1575,32'd-351,32'd-673,32'd-1755,32'd944,32'd-2385,32'd-2670,32'd-593,32'd1772,32'd2644,32'd4567,32'd-4038,32'd-1336,32'd-1287,32'd-4050,32'd977,32'd-1162,32'd-397,32'd568,32'd3786,32'd-3139,32'd519,32'd-1589,32'd-5083,32'd185,32'd-735,32'd4416,32'd-2333,32'd2917,32'd-1148,32'd3234,32'd-241,32'd-1282,32'd167,32'd4826,32'd-227,32'd456,32'd2011,32'd4299,32'd-1625,32'd-2113,32'd-3493,32'd-4936,32'd1076,32'd667,32'd-1804,32'd-1033,32'd6674,32'd-1623,32'd532,32'd1635,32'd-239,32'd-3044,32'd-92,32'd3679,32'd2729,32'd-1495,32'd-750,32'd3,32'd-6337,32'd1774,32'd2702,32'd1735,32'd2512,32'd-1485,32'd7919,32'd1345,32'd-679,32'd4909,32'd332,32'd368,32'd3566,32'd-2310,32'd892,32'd2491,32'd-207,32'd1528,32'd-1855,32'd1612,32'd1185,32'd-2208,32'd329,32'd141,32'd-1926,32'd-1674,32'd2983,32'd2364,32'd-2438,32'd-1591,32'd-5283,32'd-2443,32'd1241,32'd7163,32'd1594,32'd-3339,32'd3820,32'd-5727,32'd356,32'd-8017,32'd1444,32'd806,32'd-2340,32'd4262,32'd71,32'd4201,32'd-89,32'd-2316,32'd1262,32'd566,32'd-2478,32'd-2084,32'd7153,32'd-531,32'd5371,32'd-5927,32'd-1129,32'd2214,32'd298,32'd-254,32'd385,32'd-2197,32'd2486,32'd-3215,32'd767,32'd1180,32'd-603,32'd-1811,32'd1466,32'd2011,32'd-2705,32'd-5581,32'd-2656,32'd4479,32'd-4870,32'd-297,32'd-715,32'd12343,32'd-3615,32'd-2939,32'd1062,32'd-5537,32'd725,32'd-2937,32'd-2185,32'd1671,32'd1754,32'd2130,32'd4328,32'd1922,32'd3886,32'd589,32'd-302,32'd416,32'd-537,32'd618,32'd-2288,32'd2739,32'd-1196,32'd3093,32'd3088,32'd2827,32'd-4057,32'd1004,32'd-390,32'd1995,32'd-4448,32'd-4240,32'd1499,32'd640,32'd2900,32'd-1413,32'd-2015,32'd568,32'd-3864,32'd1290,32'd145,32'd-242,32'd-1172,32'd5034,32'd-684,32'd2800,32'd-869,32'd2912,32'd-1522,32'd5200,32'd2305,32'd502,32'd-947,32'd2062,32'd2612,32'd-2958,32'd3144,32'd2937,32'd3312,32'd-646,32'd-2478,32'd2753,32'd3244,32'd876,32'd587,32'd-2626,32'd3413,32'd1676,32'd3430,32'd-188,32'd269,32'd2897,32'd6660,32'd-3395,32'd1894,32'd1444,32'd-1013,32'd1384,32'd599,32'd526,32'd-1973,32'd-415,32'd3254,32'd-1156,32'd-2966,32'd-1469,32'd-1372,32'd-2264,32'd1229,32'd1298,32'd-1518,32'd5,32'd2152,32'd-2968,32'd-1166,32'd4624,32'd-1411,32'd-1280,32'd1459,32'd2636,32'd3608,32'd-4438,32'd322,32'd-2331,32'd1744,32'd-2465,32'd-1336,32'd-47,32'd5429,32'd1683,32'd-620,32'd-3527,32'd-3864,32'd-2351,32'd-1138,32'd1361,32'd774,32'd4604,32'd-930,32'd552,32'd-1767,32'd-2427,32'd74,32'd-2075,32'd54,32'd-3156,32'd-1884,32'd1153,32'd-1474,32'd532,32'd2015,32'd822,32'd-2288,32'd1091,32'd2208,32'd-2531,32'd4118,32'd2199,32'd-188,32'd-2148,32'd3850,32'd-1295,32'd1132,32'd3378,32'd556,32'd1608,32'd-631,32'd2258,32'd-3305,32'd2912,32'd-240,32'd5258,32'd117,32'd3923,32'd1078,32'd2337,32'd-2114,32'd-2507,32'd-7275,32'd1927,32'd3459,32'd-2707,32'd-1422,32'd-1232,32'd-3405,32'd-4577,32'd3127,32'd-228,32'd-1437,32'd2390,32'd-8125,32'd-1671,32'd3679,32'd1984,32'd4201,32'd455,32'd5083,32'd383,32'd1488,32'd-1953,32'd118,32'd-1798,32'd-1091,32'd-1346,32'd-1787,32'd-312,32'd2093,32'd-1372,32'd19,32'd-2700,32'd1093,32'd385,32'd-3674,32'd2009,32'd1821,32'd-795,32'd1702,32'd2482,32'd1315,32'd-517,32'd1059,32'd4541,32'd4802,32'd2429,32'd3303,32'd2322,32'd-3764,32'd-785,32'd-739,32'd1630,32'd-192,32'd1337,32'd4975,32'd2047,32'd-304,32'd-3168,32'd3386,32'd3894,32'd795,32'd-197,32'd-1148,32'd2663,32'd-3903,32'd5942,32'd1250,32'd3398,32'd4091,32'd-3808,32'd-4089,32'd1265,32'd6132,32'd-5253,32'd233,32'd-226,32'd-465,32'd-769,32'd-1271,32'd1697,32'd2817,32'd-2498,32'd1622,32'd-380};
    Wh[89]='{32'd4338,32'd1990,32'd-2924,32'd1013,32'd-909,32'd2098,32'd-4758,32'd-4350,32'd-2093,32'd-2531,32'd913,32'd-1522,32'd439,32'd-1662,32'd-1683,32'd-3833,32'd-446,32'd3691,32'd-591,32'd-949,32'd1524,32'd-1132,32'd-4865,32'd-1513,32'd-3359,32'd1212,32'd834,32'd257,32'd900,32'd2414,32'd903,32'd7919,32'd-6386,32'd-1710,32'd3420,32'd-1041,32'd-303,32'd1041,32'd4060,32'd-3498,32'd-1657,32'd-1993,32'd10683,32'd-1798,32'd-3757,32'd-2220,32'd-3818,32'd4082,32'd526,32'd3103,32'd-3117,32'd-3281,32'd4558,32'd3049,32'd3549,32'd8007,32'd-29,32'd5434,32'd1621,32'd4279,32'd1383,32'd196,32'd671,32'd458,32'd3100,32'd740,32'd-3217,32'd-4621,32'd-339,32'd1900,32'd3193,32'd3105,32'd-1004,32'd-3083,32'd-3605,32'd575,32'd-4924,32'd-3103,32'd4533,32'd-377,32'd-1353,32'd-1069,32'd-2294,32'd399,32'd-486,32'd-1853,32'd-2797,32'd-1212,32'd-3095,32'd-2531,32'd-1735,32'd-3312,32'd-2132,32'd-2666,32'd-3676,32'd-571,32'd-7211,32'd2878,32'd-1260,32'd-4177,32'd-728,32'd-7480,32'd-6416,32'd6186,32'd-1805,32'd-2778,32'd3837,32'd4985,32'd-6342,32'd1446,32'd99,32'd-6000,32'd2875,32'd1837,32'd-1427,32'd4511,32'd119,32'd9072,32'd2438,32'd-1842,32'd3952,32'd-206,32'd-2254,32'd1940,32'd-5053,32'd-1569,32'd-7290,32'd-1350,32'd-566,32'd-14589,32'd-700,32'd1647,32'd446,32'd2802,32'd2941,32'd1959,32'd5078,32'd1346,32'd5947,32'd-2019,32'd4416,32'd-3364,32'd8300,32'd-1282,32'd316,32'd-895,32'd-6059,32'd7792,32'd-368,32'd-749,32'd3283,32'd-1391,32'd3457,32'd562,32'd-3112,32'd14121,32'd4633,32'd-6499,32'd1072,32'd965,32'd3212,32'd-30,32'd3403,32'd-4726,32'd1569,32'd-2541,32'd-2573,32'd-2832,32'd-5161,32'd6225,32'd-1939,32'd-3469,32'd-1135,32'd-1004,32'd-673,32'd1579,32'd-3867,32'd70,32'd-4638,32'd3747,32'd-4277,32'd8779,32'd-5717,32'd3354,32'd8388,32'd999,32'd-7709,32'd1505,32'd1407,32'd1110,32'd6708,32'd9687,32'd-3549,32'd1278,32'd-3613,32'd-1101,32'd-1198,32'd-1639,32'd-1733,32'd-325,32'd-1293,32'd-2512,32'd-401,32'd476,32'd-1843,32'd-157,32'd1663,32'd9711,32'd2297,32'd-3076,32'd-2629,32'd-3120,32'd-2115,32'd1451,32'd-2083,32'd-109,32'd-4777,32'd-8857,32'd-1250,32'd-1335,32'd2219,32'd-3869,32'd-1334,32'd523,32'd-4287,32'd983,32'd1563,32'd1939,32'd-2022,32'd2849,32'd-1451,32'd1604,32'd-221,32'd-1339,32'd-1095,32'd435,32'd-5693,32'd1734,32'd5268,32'd-800,32'd6445,32'd4843,32'd1707,32'd4792,32'd3962,32'd-698,32'd2875,32'd988,32'd4995,32'd-3981,32'd6337,32'd342,32'd-3259,32'd4182,32'd2463,32'd6816,32'd2763,32'd1453,32'd-725,32'd-3017,32'd-9106,32'd-946,32'd9409,32'd221,32'd-2558,32'd2783,32'd1473,32'd-192,32'd1892,32'd1475,32'd-335,32'd2958,32'd-3425,32'd3320,32'd-3063,32'd-4479,32'd-2426,32'd-502,32'd-4645,32'd2502,32'd-4709,32'd-1604,32'd202,32'd182,32'd-1132,32'd-537,32'd4331,32'd-2707,32'd-1309,32'd3115,32'd-10791,32'd6777,32'd7182,32'd-3662,32'd-8281,32'd331,32'd1445,32'd-3991,32'd7729,32'd-3361,32'd-6176,32'd-441,32'd-9980,32'd1856,32'd2700,32'd-7348,32'd682,32'd-531,32'd1098,32'd-2849,32'd1558,32'd-8071,32'd1115,32'd430,32'd-3576,32'd-2261,32'd4592,32'd1079,32'd-10068,32'd1259,32'd-6582,32'd-1707,32'd2822,32'd-1268,32'd-2656,32'd4960,32'd-1256,32'd-971,32'd716,32'd432,32'd-7021,32'd3696,32'd2753,32'd2678,32'd-5214,32'd3811,32'd-7172,32'd2648,32'd3955,32'd-163,32'd239,32'd4821,32'd4448,32'd5532,32'd757,32'd3151,32'd-4084,32'd-1216,32'd3391,32'd718,32'd4555,32'd3891,32'd-529,32'd2309,32'd-1072,32'd-1834,32'd-2639,32'd-9936,32'd-8525,32'd-856,32'd2910,32'd3437,32'd3862,32'd-2199,32'd-1987,32'd3273,32'd-997,32'd-4667,32'd-3417,32'd-1614,32'd7646,32'd-467,32'd-2348,32'd-3793,32'd-3205,32'd1798,32'd4145,32'd3247,32'd-4079,32'd951,32'd2424,32'd-1773,32'd5336,32'd4333,32'd-3391,32'd-322,32'd756,32'd-4118,32'd-3640,32'd9501,32'd-10742,32'd3706,32'd-293,32'd-3681,32'd-1918,32'd-5839,32'd-3271,32'd3251,32'd2385,32'd-3017};
    Wh[90]='{32'd-1010,32'd466,32'd-256,32'd3769,32'd-1439,32'd-1043,32'd3210,32'd-1049,32'd-1068,32'd1256,32'd4567,32'd1824,32'd1064,32'd2915,32'd-995,32'd5244,32'd4912,32'd4150,32'd2612,32'd-3146,32'd1838,32'd-2055,32'd-295,32'd1541,32'd-2366,32'd4924,32'd1259,32'd57,32'd144,32'd6474,32'd-20,32'd4780,32'd2990,32'd1656,32'd3891,32'd1239,32'd1655,32'd-118,32'd208,32'd3955,32'd11,32'd5000,32'd-1596,32'd1655,32'd2045,32'd2573,32'd960,32'd-3588,32'd-102,32'd-3957,32'd693,32'd1040,32'd-2183,32'd2326,32'd-2912,32'd5737,32'd2462,32'd-2885,32'd4016,32'd8247,32'd-1274,32'd3474,32'd-2110,32'd-1683,32'd278,32'd1065,32'd3039,32'd9096,32'd1726,32'd2675,32'd1066,32'd3662,32'd4543,32'd157,32'd1095,32'd-2741,32'd4748,32'd-955,32'd-2363,32'd1528,32'd581,32'd386,32'd8222,32'd3427,32'd177,32'd-120,32'd166,32'd5034,32'd1342,32'd4050,32'd-416,32'd-117,32'd2661,32'd-3867,32'd5258,32'd5541,32'd-1205,32'd7749,32'd3503,32'd1718,32'd-3283,32'd-3928,32'd-1820,32'd7045,32'd-6748,32'd-787,32'd806,32'd6025,32'd1224,32'd5263,32'd405,32'd3276,32'd2038,32'd-1025,32'd-839,32'd1815,32'd1717,32'd-5771,32'd1818,32'd-3718,32'd-4265,32'd-5537,32'd-3203,32'd2009,32'd-606,32'd-392,32'd2177,32'd-2083,32'd-3105,32'd-12324,32'd-1894,32'd1997,32'd3310,32'd-3188,32'd-4899,32'd2668,32'd1475,32'd-2604,32'd3408,32'd1840,32'd-828,32'd2473,32'd-3146,32'd-1586,32'd49,32'd-1726,32'd-3740,32'd2407,32'd6445,32'd-820,32'd-4663,32'd839,32'd-642,32'd408,32'd2196,32'd3984,32'd-552,32'd-1046,32'd6030,32'd8974,32'd554,32'd-737,32'd396,32'd791,32'd-1132,32'd3325,32'd-2512,32'd2854,32'd1161,32'd-516,32'd-168,32'd1499,32'd-1347,32'd-1245,32'd-394,32'd1148,32'd-7646,32'd4196,32'd-2612,32'd2827,32'd-2016,32'd2656,32'd-1945,32'd556,32'd3762,32'd-1899,32'd2003,32'd-1337,32'd-6572,32'd1877,32'd-1207,32'd-4755,32'd4479,32'd-190,32'd2729,32'd-2145,32'd-3857,32'd787,32'd-5883,32'd-2215,32'd3881,32'd3986,32'd-1069,32'd-2209,32'd-1943,32'd-1431,32'd2077,32'd3837,32'd-4890,32'd5605,32'd4245,32'd1160,32'd4689,32'd-4453,32'd760,32'd2408,32'd-3830,32'd2261,32'd2729,32'd-3039,32'd-635,32'd1148,32'd108,32'd-1850,32'd-2471,32'd4548,32'd1802,32'd2358,32'd-1206,32'd-3134,32'd-1727,32'd-942,32'd474,32'd-4555,32'd-1263,32'd-970,32'd24,32'd1251,32'd4118,32'd1318,32'd-357,32'd4694,32'd-908,32'd-2,32'd84,32'd-1212,32'd-7338,32'd-111,32'd5537,32'd-1535,32'd4206,32'd1384,32'd1517,32'd231,32'd-3425,32'd2602,32'd-21,32'd3286,32'd1490,32'd-6762,32'd-6215,32'd5961,32'd2371,32'd6777,32'd-2844,32'd2070,32'd3349,32'd290,32'd3483,32'd-40,32'd800,32'd-9716,32'd3769,32'd4628,32'd6835,32'd-3142,32'd1398,32'd-248,32'd3840,32'd5888,32'd-111,32'd-878,32'd4516,32'd9008,32'd-1351,32'd-13,32'd338,32'd1564,32'd584,32'd-690,32'd-399,32'd-179,32'd3300,32'd-2322,32'd-4650,32'd3784,32'd4772,32'd298,32'd4257,32'd-2629,32'd2861,32'd-6538,32'd-1087,32'd588,32'd-3308,32'd10166,32'd2722,32'd207,32'd-1828,32'd1992,32'd812,32'd5209,32'd2257,32'd-807,32'd-3298,32'd-197,32'd-2360,32'd2988,32'd-605,32'd4785,32'd374,32'd1638,32'd3015,32'd222,32'd-1223,32'd1741,32'd5327,32'd2971,32'd3732,32'd7480,32'd1177,32'd-2369,32'd2192,32'd1982,32'd-1057,32'd2145,32'd-150,32'd6035,32'd530,32'd-2565,32'd301,32'd3771,32'd2844,32'd4938,32'd2995,32'd285,32'd-5478,32'd2145,32'd7192,32'd1624,32'd92,32'd-253,32'd770,32'd-2247,32'd397,32'd-3479,32'd6215,32'd-689,32'd-2392,32'd-117,32'd4145,32'd4807,32'd-1206,32'd311,32'd-2036,32'd4978,32'd-484,32'd-2790,32'd4511,32'd2121,32'd5566,32'd-567,32'd2397,32'd1903,32'd3544,32'd1520,32'd-1761,32'd-601,32'd3715,32'd1409,32'd2039,32'd7905,32'd4333,32'd-771,32'd5585,32'd6,32'd897,32'd3903,32'd1566,32'd7138,32'd-7114,32'd-3044,32'd2626,32'd906,32'd4326,32'd-1684,32'd-2907,32'd194,32'd6430,32'd-3427};
    Wh[91]='{32'd-1303,32'd-4248,32'd3586,32'd-3193,32'd326,32'd1168,32'd-5185,32'd2680,32'd-2597,32'd1248,32'd-2939,32'd-1071,32'd-1551,32'd681,32'd635,32'd-96,32'd166,32'd-5253,32'd-230,32'd-5312,32'd3334,32'd-1647,32'd1322,32'd-663,32'd2032,32'd-1106,32'd-480,32'd135,32'd-13906,32'd-1311,32'd6362,32'd-7685,32'd932,32'd-588,32'd4418,32'd1258,32'd1463,32'd669,32'd-176,32'd10791,32'd-1557,32'd-8945,32'd-3635,32'd684,32'd-2216,32'd-177,32'd2924,32'd867,32'd-504,32'd1055,32'd-2106,32'd-17,32'd5078,32'd4260,32'd-4738,32'd1557,32'd-2086,32'd5961,32'd1105,32'd-7041,32'd737,32'd5668,32'd2272,32'd-3737,32'd2235,32'd-1915,32'd573,32'd2092,32'd2149,32'd4868,32'd-872,32'd-2775,32'd5009,32'd-2976,32'd7221,32'd3698,32'd1120,32'd5541,32'd1333,32'd-4645,32'd-54,32'd5419,32'd-1204,32'd-557,32'd1166,32'd-4291,32'd153,32'd1028,32'd-547,32'd-1353,32'd-6958,32'd-1470,32'd2504,32'd2254,32'd-1099,32'd-525,32'd439,32'd-9340,32'd-4746,32'd2176,32'd-1019,32'd-4460,32'd-2481,32'd7509,32'd-2026,32'd-1934,32'd-3381,32'd2639,32'd-10380,32'd11406,32'd-2464,32'd3325,32'd1380,32'd3986,32'd23,32'd6328,32'd-9218,32'd-14091,32'd-13525,32'd-18105,32'd698,32'd7402,32'd997,32'd-4506,32'd-7631,32'd-991,32'd7607,32'd3330,32'd-1435,32'd-3435,32'd772,32'd707,32'd-1956,32'd7382,32'd-2783,32'd-3527,32'd-5693,32'd-508,32'd40,32'd-2067,32'd-6352,32'd-553,32'd-6508,32'd30,32'd-4580,32'd1103,32'd-5273,32'd771,32'd-6904,32'd67,32'd-1853,32'd-3806,32'd2019,32'd-1655,32'd4121,32'd3857,32'd-4501,32'd-785,32'd297,32'd14707,32'd-8579,32'd-4199,32'd261,32'd-1365,32'd-1826,32'd7656,32'd1972,32'd885,32'd2023,32'd-548,32'd994,32'd2854,32'd6918,32'd5561,32'd1193,32'd-2841,32'd281,32'd-1214,32'd-158,32'd1306,32'd392,32'd-3962,32'd5698,32'd-1542,32'd115,32'd-3164,32'd-1706,32'd-3090,32'd-6782,32'd-3867,32'd-1649,32'd-5927,32'd520,32'd2055,32'd1909,32'd-13906,32'd-9575,32'd1518,32'd389,32'd-936,32'd-3452,32'd3750,32'd1364,32'd6123,32'd4113,32'd1987,32'd4248,32'd1245,32'd-495,32'd-884,32'd10341,32'd2783,32'd7041,32'd286,32'd712,32'd3850,32'd-831,32'd1467,32'd2257,32'd1257,32'd2905,32'd-6547,32'd-5385,32'd2985,32'd-988,32'd-3686,32'd-4543,32'd3422,32'd543,32'd6523,32'd531,32'd1705,32'd471,32'd-3806,32'd5009,32'd6772,32'd754,32'd2027,32'd-1238,32'd-1839,32'd-6337,32'd4667,32'd3181,32'd3562,32'd-175,32'd-2932,32'd-2188,32'd6494,32'd3295,32'd-1486,32'd6914,32'd69,32'd246,32'd-4130,32'd4011,32'd-583,32'd6816,32'd3107,32'd3447,32'd13525,32'd5371,32'd491,32'd-1287,32'd762,32'd1354,32'd4711,32'd5766,32'd4758,32'd1904,32'd321,32'd-2854,32'd-5458,32'd-505,32'd2124,32'd3937,32'd4133,32'd-547,32'd3303,32'd1524,32'd3388,32'd382,32'd-454,32'd3347,32'd-5590,32'd3605,32'd-3310,32'd4326,32'd955,32'd-12089,32'd-5869,32'd-9746,32'd-8056,32'd550,32'd5380,32'd-12,32'd8081,32'd-1143,32'd4394,32'd3876,32'd-1801,32'd3825,32'd-88,32'd5458,32'd-95,32'd4187,32'd8535,32'd3259,32'd341,32'd844,32'd3615,32'd535,32'd935,32'd1295,32'd2448,32'd-4167,32'd838,32'd-2888,32'd-366,32'd5688,32'd-6567,32'd-9663,32'd-1791,32'd-4772,32'd565,32'd-2276,32'd-2578,32'd-4440,32'd-1383,32'd3684,32'd-1763,32'd-1345,32'd337,32'd-2846,32'd511,32'd-747,32'd-3110,32'd-3437,32'd4792,32'd-3581,32'd3491,32'd-2423,32'd-2294,32'd1125,32'd725,32'd29,32'd-2690,32'd-3002,32'd948,32'd-9926,32'd-568,32'd1209,32'd-4768,32'd316,32'd1313,32'd-7119,32'd-3466,32'd516,32'd9355,32'd1109,32'd-3408,32'd4628,32'd1850,32'd3007,32'd-5229,32'd2756,32'd-5322,32'd-907,32'd-4379,32'd-1542,32'd2222,32'd560,32'd-3017,32'd-2028,32'd-1607,32'd374,32'd321,32'd-8823,32'd1596,32'd-1899,32'd-493,32'd-3239,32'd-7607,32'd-429,32'd1149,32'd-561,32'd4150,32'd7480,32'd2985,32'd-3427,32'd-2218,32'd-3276,32'd3085,32'd4272,32'd-1489,32'd9096,32'd5278,32'd549,32'd2956,32'd2512,32'd831};
    Wh[92]='{32'd-1851,32'd1235,32'd-203,32'd2871,32'd-133,32'd1516,32'd-491,32'd-3330,32'd-1760,32'd-2517,32'd1693,32'd-155,32'd388,32'd1352,32'd2222,32'd871,32'd4396,32'd-867,32'd2941,32'd229,32'd419,32'd2196,32'd-4333,32'd-133,32'd1331,32'd1446,32'd1362,32'd1029,32'd5434,32'd111,32'd-1329,32'd1285,32'd4536,32'd1450,32'd1193,32'd836,32'd-775,32'd1877,32'd-1143,32'd1057,32'd-1455,32'd1467,32'd-1005,32'd6054,32'd-1361,32'd3427,32'd1606,32'd-597,32'd5537,32'd965,32'd8203,32'd-782,32'd-2379,32'd1816,32'd6743,32'd-5146,32'd-472,32'd-5019,32'd-1575,32'd-2332,32'd-747,32'd4484,32'd842,32'd2766,32'd4597,32'd-2661,32'd1218,32'd4545,32'd-4023,32'd-2983,32'd1001,32'd-4345,32'd-977,32'd567,32'd1489,32'd7094,32'd7504,32'd3994,32'd-1683,32'd-266,32'd1065,32'd2502,32'd-632,32'd2382,32'd-2432,32'd3051,32'd-265,32'd-4628,32'd2834,32'd-2160,32'd-822,32'd-2570,32'd-850,32'd2800,32'd-817,32'd-570,32'd-1307,32'd-662,32'd2844,32'd-1810,32'd2727,32'd-4299,32'd615,32'd-742,32'd-580,32'd-1845,32'd4980,32'd3315,32'd17265,32'd1176,32'd194,32'd-2376,32'd3041,32'd-1545,32'd-4785,32'd-1550,32'd-654,32'd4921,32'd-4265,32'd3291,32'd-206,32'd489,32'd3295,32'd-2702,32'd6494,32'd-4140,32'd-4162,32'd2937,32'd1849,32'd2937,32'd-3505,32'd1619,32'd-3354,32'd-1654,32'd-2897,32'd-1235,32'd-227,32'd1431,32'd-474,32'd-4055,32'd695,32'd-3281,32'd-459,32'd1574,32'd-2697,32'd-2138,32'd103,32'd3984,32'd-56,32'd1440,32'd-433,32'd-3161,32'd-444,32'd173,32'd-3557,32'd2432,32'd5341,32'd-2344,32'd-138,32'd-41,32'd-5385,32'd-1210,32'd5263,32'd8515,32'd-5561,32'd-260,32'd3000,32'd1518,32'd-3398,32'd780,32'd1708,32'd-2343,32'd6577,32'd-5097,32'd-2612,32'd5478,32'd-1868,32'd-5322,32'd-1374,32'd2851,32'd-1088,32'd3244,32'd57,32'd-709,32'd-1490,32'd-278,32'd832,32'd-3063,32'd4677,32'd-3535,32'd-3586,32'd3632,32'd-1564,32'd-2819,32'd-3984,32'd850,32'd-1912,32'd-473,32'd-5180,32'd-6845,32'd1188,32'd-1165,32'd-3066,32'd4890,32'd2426,32'd808,32'd-2338,32'd-5244,32'd-1579,32'd-1206,32'd933,32'd-3461,32'd3852,32'd-552,32'd-1419,32'd-2846,32'd300,32'd3967,32'd-2990,32'd-665,32'd1468,32'd-1590,32'd-4262,32'd-7553,32'd6137,32'd6206,32'd2834,32'd2384,32'd-656,32'd3532,32'd747,32'd-508,32'd2199,32'd-3249,32'd-6552,32'd-3476,32'd1501,32'd-592,32'd-3103,32'd1292,32'd6645,32'd2551,32'd608,32'd-5815,32'd2661,32'd4731,32'd2731,32'd622,32'd-655,32'd-1406,32'd768,32'd-7290,32'd-1240,32'd-3417,32'd-599,32'd1859,32'd-2227,32'd1765,32'd4257,32'd685,32'd3806,32'd1364,32'd-10292,32'd-855,32'd-4401,32'd-2526,32'd61,32'd182,32'd-7265,32'd2413,32'd-1206,32'd5000,32'd4831,32'd723,32'd-4394,32'd-2008,32'd-1923,32'd-1423,32'd-639,32'd1638,32'd-1923,32'd2237,32'd2810,32'd-3415,32'd1180,32'd424,32'd313,32'd27,32'd-2341,32'd2343,32'd-4909,32'd-4177,32'd3903,32'd1248,32'd654,32'd5083,32'd-1610,32'd156,32'd1828,32'd988,32'd-4309,32'd290,32'd-3520,32'd2880,32'd1597,32'd943,32'd1844,32'd-3894,32'd1226,32'd-3381,32'd-2258,32'd6064,32'd-1536,32'd1601,32'd1564,32'd5395,32'd1352,32'd-847,32'd2332,32'd5268,32'd1292,32'd-2487,32'd-1628,32'd961,32'd746,32'd4069,32'd-1026,32'd4248,32'd-4396,32'd-1157,32'd5131,32'd2410,32'd-1284,32'd572,32'd2319,32'd1205,32'd-59,32'd1037,32'd-3647,32'd3669,32'd802,32'd3027,32'd-1101,32'd-3874,32'd-795,32'd-1478,32'd-4091,32'd-478,32'd5854,32'd1555,32'd-2585,32'd5336,32'd3513,32'd1524,32'd1735,32'd-1691,32'd1340,32'd8540,32'd-8676,32'd5263,32'd-3393,32'd8032,32'd2868,32'd7231,32'd-7631,32'd2346,32'd-897,32'd1110,32'd-4921,32'd-4855,32'd707,32'd-281,32'd4533,32'd-3095,32'd738,32'd1936,32'd-960,32'd2871,32'd-3310,32'd1599,32'd-4458,32'd1636,32'd3889,32'd-2519,32'd-3361,32'd-4731,32'd819,32'd-4794,32'd4575,32'd-3554,32'd-2277,32'd-3552,32'd-2785,32'd3464,32'd-874,32'd4643,32'd830,32'd-4260,32'd3134,32'd-899};
    Wh[93]='{32'd-1640,32'd-1614,32'd-1881,32'd-128,32'd-4182,32'd3315,32'd-5834,32'd922,32'd-2595,32'd-3334,32'd-5390,32'd5180,32'd2844,32'd-152,32'd-3691,32'd5048,32'd-12382,32'd-974,32'd-3076,32'd-3374,32'd-2714,32'd-3725,32'd352,32'd-4680,32'd-3688,32'd-4650,32'd-575,32'd-2293,32'd-8666,32'd-4309,32'd-4621,32'd-9980,32'd-12812,32'd-3061,32'd8789,32'd-1188,32'd-3134,32'd-4536,32'd5156,32'd-331,32'd2452,32'd807,32'd38,32'd4536,32'd-6484,32'd-8681,32'd-848,32'd-4980,32'd-4028,32'd6381,32'd1811,32'd-10078,32'd-1834,32'd-2863,32'd-5278,32'd-3168,32'd-3752,32'd6269,32'd-6411,32'd18183,32'd3867,32'd920,32'd-4523,32'd-3483,32'd-5698,32'd-4631,32'd-1693,32'd-4577,32'd476,32'd1884,32'd6118,32'd2308,32'd-3012,32'd-9311,32'd-5600,32'd-3764,32'd5957,32'd-5590,32'd2087,32'd-2521,32'd-101,32'd-7373,32'd-5166,32'd-1337,32'd534,32'd-2403,32'd648,32'd-3239,32'd1721,32'd3842,32'd-2834,32'd-11542,32'd-6328,32'd-5541,32'd-5336,32'd-892,32'd2897,32'd-6381,32'd-5336,32'd-3229,32'd-6191,32'd-3881,32'd-5766,32'd5244,32'd-1424,32'd-4169,32'd-3151,32'd-10126,32'd848,32'd-4379,32'd-2927,32'd-3027,32'd3105,32'd2846,32'd-4091,32'd5141,32'd-7607,32'd-1674,32'd243,32'd3703,32'd5219,32'd4907,32'd1712,32'd-2298,32'd-1931,32'd625,32'd-8291,32'd5947,32'd4326,32'd9892,32'd3017,32'd2832,32'd-824,32'd3625,32'd-3200,32'd-194,32'd-7856,32'd-826,32'd-748,32'd2,32'd-1256,32'd3376,32'd-6513,32'd-2386,32'd-352,32'd-4167,32'd-3999,32'd-509,32'd-11503,32'd851,32'd2232,32'd1552,32'd2929,32'd-1849,32'd-1768,32'd-7441,32'd-10839,32'd-3452,32'd-8476,32'd-31289,32'd4555,32'd2963,32'd5371,32'd-921,32'd1527,32'd-681,32'd197,32'd2413,32'd-5327,32'd2182,32'd-2423,32'd-2866,32'd4060,32'd2556,32'd3591,32'd1976,32'd-1220,32'd-3718,32'd-89,32'd870,32'd8549,32'd10859,32'd4494,32'd4765,32'd6972,32'd-567,32'd6469,32'd2790,32'd902,32'd2188,32'd-2575,32'd345,32'd-2985,32'd-232,32'd5390,32'd4233,32'd6767,32'd-3144,32'd-5083,32'd272,32'd-2371,32'd3168,32'd3400,32'd7968,32'd-3435,32'd3120,32'd5244,32'd5004,32'd-5590,32'd-6982,32'd4609,32'd-10878,32'd-7216,32'd-4001,32'd-1064,32'd4177,32'd2910,32'd-2121,32'd-5239,32'd1319,32'd452,32'd-10117,32'd-643,32'd-6069,32'd-4843,32'd-9785,32'd-3645,32'd-2988,32'd4665,32'd3161,32'd-3811,32'd9389,32'd334,32'd1896,32'd4831,32'd-986,32'd-3630,32'd-3630,32'd-2517,32'd2073,32'd3469,32'd7832,32'd1971,32'd-7539,32'd1666,32'd1868,32'd-4704,32'd-988,32'd-1840,32'd-3447,32'd-2612,32'd-3281,32'd388,32'd992,32'd293,32'd4899,32'd-989,32'd894,32'd-1712,32'd-6376,32'd-6987,32'd-451,32'd4904,32'd-164,32'd-2152,32'd1865,32'd2196,32'd-2993,32'd1429,32'd1191,32'd-1105,32'd7695,32'd-9355,32'd-183,32'd-3029,32'd1428,32'd-8500,32'd2150,32'd-841,32'd2927,32'd-2644,32'd2329,32'd5883,32'd9223,32'd817,32'd-3181,32'd-897,32'd3815,32'd-7260,32'd2866,32'd-2724,32'd12021,32'd-3908,32'd5385,32'd-2976,32'd698,32'd-2697,32'd1506,32'd-2048,32'd11132,32'd-9296,32'd6596,32'd-9521,32'd-2587,32'd-751,32'd-5043,32'd4189,32'd-901,32'd-5537,32'd-3796,32'd-8081,32'd-7441,32'd-1012,32'd-1949,32'd988,32'd7661,32'd9404,32'd-2714,32'd-12714,32'd-10224,32'd-10234,32'd-11660,32'd-2663,32'd-406,32'd-215,32'd331,32'd-2998,32'd-2104,32'd875,32'd-586,32'd-6801,32'd3605,32'd-1147,32'd-597,32'd-8549,32'd5380,32'd-1035,32'd-8349,32'd-2885,32'd7548,32'd1124,32'd5395,32'd2166,32'd13554,32'd524,32'd-615,32'd-1024,32'd977,32'd-7553,32'd1234,32'd9882,32'd7983,32'd-5000,32'd4611,32'd-3706,32'd1235,32'd-5278,32'd-8481,32'd-1820,32'd-249,32'd-508,32'd6040,32'd-117,32'd-3728,32'd3422,32'd-7543,32'd-1329,32'd4497,32'd-7045,32'd2565,32'd720,32'd5541,32'd-8027,32'd-588,32'd-8813,32'd4929,32'd-309,32'd1638,32'd1160,32'd-1282,32'd-372,32'd3598,32'd728,32'd6972,32'd-5742,32'd3527,32'd-8544,32'd-1152,32'd-5981,32'd2398,32'd2117,32'd-27,32'd-4011,32'd10166,32'd2712,32'd3066,32'd-4599,32'd4799,32'd-6723,32'd4074};
    Wh[94]='{32'd-445,32'd-4970,32'd173,32'd2902,32'd-1522,32'd-68,32'd-1712,32'd-3845,32'd6635,32'd3471,32'd1616,32'd2322,32'd-2346,32'd-101,32'd-6938,32'd-386,32'd-7075,32'd-250,32'd-208,32'd1866,32'd37,32'd6137,32'd3654,32'd2415,32'd244,32'd-409,32'd1677,32'd112,32'd4201,32'd850,32'd3334,32'd1591,32'd-7656,32'd4294,32'd-458,32'd1302,32'd-3498,32'd-2489,32'd-4272,32'd2369,32'd1231,32'd-1302,32'd-1028,32'd-718,32'd-231,32'd-4206,32'd1973,32'd2873,32'd-2047,32'd-1542,32'd7060,32'd139,32'd-5288,32'd2371,32'd1861,32'd-2934,32'd342,32'd-1226,32'd2406,32'd1140,32'd4294,32'd-2464,32'd-2551,32'd4448,32'd993,32'd5405,32'd-2210,32'd3684,32'd-263,32'd-227,32'd-3903,32'd-6591,32'd-587,32'd-2756,32'd-710,32'd1751,32'd-2897,32'd2208,32'd-3459,32'd3078,32'd2998,32'd-7421,32'd2036,32'd54,32'd4057,32'd-2912,32'd-2851,32'd1679,32'd1068,32'd706,32'd-462,32'd6635,32'd-636,32'd1058,32'd-5288,32'd395,32'd1308,32'd878,32'd-4711,32'd2073,32'd-2006,32'd9277,32'd3698,32'd-16386,32'd2004,32'd907,32'd-2482,32'd5688,32'd10273,32'd-5991,32'd-92,32'd-4379,32'd12666,32'd-7973,32'd5830,32'd2081,32'd1318,32'd5517,32'd-3249,32'd8364,32'd-3068,32'd2714,32'd-11826,32'd-12324,32'd737,32'd6176,32'd-3830,32'd3786,32'd4892,32'd-6313,32'd-1829,32'd1000,32'd8623,32'd-12744,32'd837,32'd645,32'd-1184,32'd3811,32'd2092,32'd1904,32'd4682,32'd-225,32'd7602,32'd-1940,32'd1713,32'd-10869,32'd7797,32'd-10234,32'd2697,32'd-3583,32'd-3398,32'd-4562,32'd-10078,32'd2504,32'd-2260,32'd-7060,32'd-8901,32'd-5581,32'd-2109,32'd-12246,32'd11074,32'd-1915,32'd-95,32'd-5209,32'd2805,32'd-4194,32'd1473,32'd-3051,32'd1890,32'd-5585,32'd4763,32'd1154,32'd-2479,32'd-5786,32'd-3264,32'd678,32'd2854,32'd2683,32'd5947,32'd-2678,32'd2061,32'd-6254,32'd-183,32'd1519,32'd-439,32'd376,32'd-783,32'd732,32'd14189,32'd877,32'd-4926,32'd-6801,32'd-8339,32'd1777,32'd1334,32'd7456,32'd-3562,32'd3562,32'd-3493,32'd1909,32'd166,32'd-84,32'd-3891,32'd5747,32'd-4101,32'd-451,32'd-6586,32'd-3750,32'd-4409,32'd3317,32'd-5854,32'd-8056,32'd3173,32'd4311,32'd-419,32'd6787,32'd-5615,32'd-6767,32'd-2410,32'd8535,32'd-677,32'd5742,32'd-237,32'd-6225,32'd4140,32'd6240,32'd3842,32'd318,32'd1754,32'd-2604,32'd-332,32'd-4934,32'd1335,32'd1069,32'd-8056,32'd-1713,32'd-2822,32'd-5161,32'd-1794,32'd3649,32'd-4167,32'd1833,32'd1737,32'd-7094,32'd-1895,32'd-1335,32'd-4814,32'd-2066,32'd-485,32'd2106,32'd-1507,32'd-2832,32'd365,32'd1798,32'd2243,32'd-2103,32'd-4682,32'd1021,32'd-2254,32'd-12050,32'd3725,32'd-2325,32'd3454,32'd63,32'd2136,32'd-1219,32'd-4218,32'd-11416,32'd-267,32'd-503,32'd-684,32'd6840,32'd-2995,32'd1169,32'd2751,32'd-5751,32'd-2203,32'd-342,32'd1188,32'd4057,32'd-3547,32'd-3935,32'd-1632,32'd3603,32'd-115,32'd-7460,32'd-5771,32'd-7202,32'd-3876,32'd-1238,32'd3842,32'd-7973,32'd-4843,32'd-3911,32'd4125,32'd-11650,32'd-3388,32'd-2199,32'd-5581,32'd5927,32'd171,32'd-7456,32'd-41,32'd-406,32'd-1785,32'd-2558,32'd2285,32'd4479,32'd5361,32'd4675,32'd-5126,32'd-1926,32'd-1030,32'd3659,32'd-3256,32'd-6118,32'd4826,32'd806,32'd-7231,32'd-2006,32'd5258,32'd10791,32'd-4094,32'd849,32'd3144,32'd3037,32'd4201,32'd2310,32'd-1228,32'd1585,32'd3098,32'd5400,32'd-7558,32'd-1341,32'd57,32'd4033,32'd-3850,32'd-6513,32'd-2036,32'd-3383,32'd158,32'd-3430,32'd-646,32'd-5878,32'd-2387,32'd3623,32'd6225,32'd513,32'd1943,32'd-1790,32'd-1926,32'd-548,32'd-3994,32'd1326,32'd8330,32'd4213,32'd-911,32'd-2017,32'd4125,32'd5605,32'd6181,32'd-7519,32'd-2413,32'd7275,32'd-1638,32'd1513,32'd-2712,32'd2279,32'd-1408,32'd-431,32'd2683,32'd4128,32'd-508,32'd-1896,32'd-2465,32'd-5351,32'd5454,32'd-194,32'd21,32'd9384,32'd1242,32'd6308,32'd-3505,32'd894,32'd-4599,32'd-3281,32'd-3176,32'd-3479,32'd785,32'd7211,32'd3186,32'd2875,32'd-4091,32'd2856,32'd1851,32'd-4870,32'd4003,32'd3393,32'd-4406,32'd1495};
    Wh[95]='{32'd-239,32'd-5756,32'd2705,32'd-4116,32'd330,32'd-1119,32'd-5161,32'd-3032,32'd5585,32'd1517,32'd-1752,32'd1511,32'd-419,32'd-7739,32'd-4201,32'd-2827,32'd-3710,32'd498,32'd-172,32'd939,32'd193,32'd-2144,32'd6206,32'd-2119,32'd-1385,32'd2734,32'd-3176,32'd1524,32'd-1751,32'd1562,32'd-2597,32'd-623,32'd-5029,32'd1676,32'd-5078,32'd323,32'd-347,32'd-2263,32'd534,32'd-3110,32'd-7197,32'd-3251,32'd-7827,32'd87,32'd725,32'd-5541,32'd-3105,32'd1684,32'd-5141,32'd-490,32'd-7548,32'd1034,32'd2563,32'd-689,32'd4370,32'd-11289,32'd-2225,32'd-1540,32'd-4145,32'd-4799,32'd-1285,32'd-2973,32'd-2963,32'd6962,32'd-3215,32'd-641,32'd-888,32'd1557,32'd1250,32'd405,32'd1027,32'd5576,32'd-1357,32'd3901,32'd296,32'd-2827,32'd-5922,32'd3889,32'd-3906,32'd2288,32'd988,32'd-5444,32'd-709,32'd934,32'd4777,32'd-5532,32'd90,32'd-3154,32'd-2335,32'd3652,32'd-1477,32'd-4025,32'd-1038,32'd3361,32'd2269,32'd-1423,32'd-2868,32'd3012,32'd576,32'd-5698,32'd-2321,32'd-716,32'd-3793,32'd2617,32'd-192,32'd1411,32'd1651,32'd1381,32'd-3405,32'd2636,32'd-4587,32'd3408,32'd-6328,32'd-1003,32'd-3754,32'd-982,32'd-2314,32'd1342,32'd1645,32'd81,32'd-3134,32'd-2355,32'd4189,32'd-1155,32'd-5083,32'd-3818,32'd6879,32'd-2429,32'd7290,32'd-1614,32'd1040,32'd49,32'd-2504,32'd935,32'd-1074,32'd-2956,32'd-6396,32'd2028,32'd415,32'd-847,32'd3569,32'd-376,32'd4301,32'd1206,32'd-2169,32'd-729,32'd-26,32'd-764,32'd1809,32'd1833,32'd-2078,32'd2246,32'd-380,32'd-3327,32'd-7343,32'd5454,32'd-1850,32'd-2707,32'd3386,32'd-4682,32'd-4887,32'd-5288,32'd359,32'd-3022,32'd-5156,32'd1499,32'd2875,32'd3928,32'd-858,32'd-401,32'd773,32'd-1885,32'd4792,32'd-207,32'd1143,32'd-1140,32'd1536,32'd4282,32'd1121,32'd102,32'd-2344,32'd5258,32'd-4282,32'd4885,32'd1071,32'd-1994,32'd-3974,32'd-253,32'd8608,32'd-2349,32'd1324,32'd4113,32'd4868,32'd3674,32'd-2326,32'd-5610,32'd1418,32'd-1142,32'd3920,32'd-1168,32'd2705,32'd4589,32'd4377,32'd-2059,32'd-3808,32'd-1313,32'd2822,32'd885,32'd-235,32'd-3920,32'd-5527,32'd2592,32'd-3542,32'd-2563,32'd3676,32'd-290,32'd812,32'd-7788,32'd5200,32'd1130,32'd933,32'd4211,32'd5380,32'd-830,32'd-7954,32'd1074,32'd-1879,32'd2231,32'd-2174,32'd391,32'd20,32'd-1112,32'd79,32'd703,32'd1347,32'd-2580,32'd1175,32'd2153,32'd6196,32'd219,32'd1669,32'd4509,32'd-10468,32'd4741,32'd-3022,32'd-928,32'd-2310,32'd-3200,32'd4084,32'd-4157,32'd-1789,32'd3576,32'd-2885,32'd-664,32'd-4670,32'd-4113,32'd374,32'd106,32'd-1121,32'd5864,32'd-1483,32'd1594,32'd-4638,32'd1855,32'd1391,32'd781,32'd-6015,32'd317,32'd2370,32'd1994,32'd-3122,32'd-78,32'd-1362,32'd855,32'd1185,32'd-3203,32'd3635,32'd1546,32'd-2939,32'd1506,32'd-5703,32'd-625,32'd2731,32'd6015,32'd2041,32'd-3530,32'd2678,32'd523,32'd499,32'd-3476,32'd1090,32'd6093,32'd-1239,32'd7324,32'd2222,32'd-2717,32'd3710,32'd-1937,32'd1824,32'd1634,32'd2280,32'd-2346,32'd-1146,32'd-5327,32'd-3908,32'd-5444,32'd2078,32'd792,32'd-1071,32'd-6274,32'd4782,32'd-672,32'd-738,32'd-4086,32'd1623,32'd-2440,32'd2304,32'd-1013,32'd2325,32'd715,32'd-1159,32'd-2445,32'd2141,32'd-889,32'd-2895,32'd3303,32'd1329,32'd-970,32'd1934,32'd997,32'd-2680,32'd-5161,32'd703,32'd1056,32'd2322,32'd-4008,32'd-1638,32'd-5434,32'd423,32'd3779,32'd-4650,32'd1910,32'd-4787,32'd1348,32'd3647,32'd-2529,32'd-356,32'd3986,32'd1839,32'd-3159,32'd-4428,32'd2044,32'd-1390,32'd429,32'd2034,32'd-1591,32'd3020,32'd-4873,32'd163,32'd-5327,32'd-915,32'd164,32'd162,32'd-4794,32'd-2169,32'd-5029,32'd-4526,32'd3374,32'd-631,32'd2119,32'd1265,32'd-2402,32'd-1237,32'd-3562,32'd-9624,32'd3706,32'd-819,32'd942,32'd-1256,32'd4038,32'd-4641,32'd-2714,32'd-59,32'd-1822,32'd-1040,32'd1315,32'd3188,32'd56,32'd314,32'd-2636,32'd-1566,32'd2078,32'd-3688,32'd-1312,32'd2247,32'd4885,32'd-816,32'd-2988,32'd-177,32'd-2132};
    Wh[96]='{32'd-159,32'd-3730,32'd-986,32'd-4277,32'd-1562,32'd1226,32'd-1132,32'd619,32'd-4331,32'd-267,32'd-3281,32'd-662,32'd-7,32'd-702,32'd1325,32'd-3247,32'd-3015,32'd574,32'd569,32'd-2702,32'd-1877,32'd-2250,32'd2010,32'd-1441,32'd493,32'd-2204,32'd-3186,32'd-1650,32'd1885,32'd-306,32'd-819,32'd-305,32'd-1104,32'd1058,32'd322,32'd142,32'd697,32'd2264,32'd-704,32'd-4572,32'd1632,32'd-3342,32'd2399,32'd-3942,32'd824,32'd852,32'd464,32'd-2780,32'd791,32'd434,32'd2414,32'd-1170,32'd-4338,32'd2814,32'd1560,32'd-639,32'd283,32'd580,32'd-2744,32'd-1464,32'd-335,32'd-2041,32'd1339,32'd-7172,32'd-975,32'd-2357,32'd144,32'd-5112,32'd2023,32'd-698,32'd3454,32'd480,32'd-2792,32'd-5957,32'd-847,32'd-4035,32'd260,32'd-4919,32'd-850,32'd-3195,32'd2418,32'd-4260,32'd-4047,32'd1650,32'd191,32'd-3784,32'd1237,32'd-552,32'd-5439,32'd2147,32'd-1862,32'd-8911,32'd-3356,32'd1514,32'd-5400,32'd-2475,32'd2502,32'd-2369,32'd-1730,32'd-494,32'd2973,32'd-71,32'd-4069,32'd-4770,32'd5405,32'd-2958,32'd-2893,32'd-4020,32'd-1002,32'd770,32'd10,32'd6523,32'd5097,32'd-38,32'd-4145,32'd822,32'd174,32'd1956,32'd-4145,32'd-3571,32'd3955,32'd3769,32'd2270,32'd-2241,32'd3591,32'd-3146,32'd-279,32'd139,32'd2656,32'd522,32'd3364,32'd510,32'd-99,32'd653,32'd6787,32'd-4367,32'd-6884,32'd3037,32'd-8364,32'd3288,32'd-1940,32'd1423,32'd2233,32'd1693,32'd-4523,32'd3859,32'd571,32'd3273,32'd-9116,32'd2822,32'd-953,32'd-60,32'd88,32'd-563,32'd-4416,32'd-3142,32'd3276,32'd-1458,32'd1922,32'd-6811,32'd3032,32'd-704,32'd-1599,32'd3151,32'd1608,32'd792,32'd-624,32'd-504,32'd-1175,32'd4484,32'd2049,32'd-3256,32'd-4904,32'd-3376,32'd-1149,32'd2161,32'd448,32'd-2106,32'd1232,32'd-4890,32'd895,32'd-4631,32'd-1934,32'd3928,32'd393,32'd780,32'd-8325,32'd-3701,32'd-2308,32'd7954,32'd-168,32'd-1106,32'd-1281,32'd4492,32'd543,32'd33,32'd1235,32'd-1217,32'd-1750,32'd3217,32'd-1196,32'd-2714,32'd-525,32'd265,32'd-2286,32'd905,32'd2624,32'd-1911,32'd775,32'd-2836,32'd517,32'd-2561,32'd-7431,32'd4946,32'd-2301,32'd637,32'd2578,32'd5688,32'd908,32'd-2998,32'd360,32'd-554,32'd-1430,32'd1149,32'd636,32'd-773,32'd17,32'd908,32'd-129,32'd-3305,32'd-1137,32'd-6508,32'd-4333,32'd638,32'd-239,32'd1789,32'd-77,32'd808,32'd-1189,32'd-1800,32'd-1442,32'd-2712,32'd946,32'd-879,32'd3046,32'd1026,32'd2773,32'd702,32'd-4245,32'd214,32'd-2575,32'd-991,32'd-3679,32'd-613,32'd-134,32'd-2252,32'd3657,32'd2491,32'd-345,32'd5605,32'd541,32'd2070,32'd-3598,32'd-1802,32'd-1039,32'd2858,32'd-1569,32'd446,32'd-372,32'd3159,32'd-5302,32'd952,32'd3317,32'd94,32'd-1436,32'd4216,32'd2604,32'd54,32'd-2159,32'd-1121,32'd-3281,32'd-3684,32'd-3017,32'd470,32'd1918,32'd3278,32'd683,32'd-4289,32'd-1181,32'd4282,32'd1452,32'd4465,32'd-3227,32'd-1046,32'd-2770,32'd-3889,32'd-3242,32'd-1566,32'd-852,32'd3808,32'd-2502,32'd2192,32'd-2761,32'd-752,32'd-1203,32'd-6347,32'd-1225,32'd-6030,32'd-1457,32'd-4497,32'd-1369,32'd-4785,32'd-3024,32'd-4074,32'd-1005,32'd-9082,32'd1304,32'd-158,32'd1271,32'd-9174,32'd-886,32'd-2636,32'd-3676,32'd-1628,32'd3488,32'd-2888,32'd-4965,32'd3051,32'd305,32'd657,32'd-3845,32'd-762,32'd-5800,32'd2988,32'd162,32'd-1506,32'd4248,32'd-5297,32'd2011,32'd310,32'd2332,32'd1113,32'd91,32'd-6098,32'd1922,32'd-1290,32'd7851,32'd-721,32'd-9941,32'd2536,32'd2785,32'd-2888,32'd989,32'd1968,32'd5229,32'd1749,32'd1760,32'd-755,32'd4169,32'd-5019,32'd-1053,32'd-1856,32'd-2478,32'd-4318,32'd5405,32'd1032,32'd-1678,32'd300,32'd-1021,32'd3356,32'd-3044,32'd-1129,32'd-346,32'd3232,32'd-2128,32'd-3283,32'd2668,32'd3200,32'd138,32'd-397,32'd-4272,32'd3935,32'd-2056,32'd271,32'd-4936,32'd659,32'd-1303,32'd-2337,32'd-2692,32'd-5302,32'd1241,32'd-4372,32'd720,32'd-143,32'd480,32'd3854,32'd11835,32'd-1016,32'd-2498,32'd1826};
    Wh[97]='{32'd2137,32'd767,32'd-653,32'd-2775,32'd1867,32'd1445,32'd-5009,32'd-6166,32'd-847,32'd3520,32'd-914,32'd-2416,32'd2868,32'd1164,32'd-2902,32'd4665,32'd7446,32'd6440,32'd-3569,32'd2783,32'd1365,32'd-987,32'd3122,32'd1437,32'd-617,32'd-1849,32'd3979,32'd1949,32'd303,32'd3435,32'd-264,32'd-282,32'd1035,32'd-3066,32'd5034,32'd711,32'd2247,32'd-1685,32'd-2304,32'd2452,32'd-107,32'd10,32'd-6943,32'd-6840,32'd-186,32'd-1390,32'd-2993,32'd-6782,32'd-1921,32'd1589,32'd1301,32'd-485,32'd-3803,32'd3500,32'd596,32'd-2343,32'd1558,32'd-94,32'd-736,32'd13300,32'd-1655,32'd-2915,32'd-5043,32'd2805,32'd2413,32'd518,32'd-925,32'd-1545,32'd2108,32'd-2614,32'd1270,32'd-92,32'd3095,32'd-4348,32'd-1583,32'd4143,32'd-393,32'd3098,32'd422,32'd5356,32'd-4255,32'd-12812,32'd-2558,32'd-2060,32'd256,32'd3666,32'd-872,32'd-542,32'd1633,32'd5288,32'd-2917,32'd4726,32'd-540,32'd-5273,32'd-9272,32'd-574,32'd-2292,32'd-286,32'd-2423,32'd-3903,32'd-10615,32'd-1218,32'd908,32'd-3896,32'd491,32'd-1943,32'd4753,32'd-3100,32'd1205,32'd-2941,32'd738,32'd-1065,32'd-3547,32'd-1335,32'd-3193,32'd-3750,32'd3200,32'd4699,32'd7104,32'd7973,32'd783,32'd1194,32'd3903,32'd5766,32'd-8452,32'd-4372,32'd3696,32'd4699,32'd2102,32'd2971,32'd-5058,32'd-4323,32'd-4665,32'd4123,32'd-6972,32'd5429,32'd-108,32'd-4829,32'd3896,32'd-5629,32'd12109,32'd-1213,32'd-1701,32'd-6235,32'd853,32'd-7885,32'd-194,32'd-10009,32'd298,32'd-2230,32'd2469,32'd-4436,32'd2995,32'd-7065,32'd-1147,32'd-1993,32'd-266,32'd-1207,32'd2175,32'd1222,32'd13291,32'd-2482,32'd1453,32'd-10371,32'd-1473,32'd2229,32'd994,32'd3278,32'd2292,32'd-2233,32'd-3947,32'd3432,32'd-5073,32'd-8432,32'd-2330,32'd4750,32'd-3469,32'd-882,32'd-881,32'd-509,32'd-2108,32'd1937,32'd-4565,32'd-299,32'd1583,32'd3205,32'd2719,32'd-3798,32'd13154,32'd4709,32'd1964,32'd1563,32'd-3635,32'd-3151,32'd-1528,32'd-4782,32'd-2137,32'd4116,32'd1369,32'd-2381,32'd-335,32'd2880,32'd1799,32'd2568,32'd-2012,32'd764,32'd5078,32'd-2203,32'd-6191,32'd4699,32'd3300,32'd-869,32'd5712,32'd-6406,32'd3486,32'd2113,32'd-2192,32'd-4809,32'd-1632,32'd1851,32'd3579,32'd1729,32'd1948,32'd995,32'd3276,32'd1088,32'd-595,32'd1948,32'd-897,32'd1931,32'd-3298,32'd-2841,32'd5781,32'd-1771,32'd495,32'd-7006,32'd-980,32'd-407,32'd-223,32'd-2702,32'd2165,32'd-588,32'd551,32'd5336,32'd-2541,32'd889,32'd601,32'd2873,32'd231,32'd-4948,32'd-4,32'd1953,32'd2167,32'd4318,32'd1884,32'd992,32'd2448,32'd3471,32'd2226,32'd-4782,32'd-1412,32'd8242,32'd6381,32'd-1212,32'd-3078,32'd0,32'd-2539,32'd2978,32'd2247,32'd-3129,32'd-1896,32'd-3283,32'd-2592,32'd6010,32'd-704,32'd-1012,32'd7758,32'd-1951,32'd3723,32'd-3037,32'd-2709,32'd-1488,32'd8955,32'd3803,32'd2250,32'd3122,32'd-1875,32'd-2248,32'd5170,32'd3044,32'd-4423,32'd11904,32'd-1356,32'd-2785,32'd-82,32'd-5029,32'd3688,32'd-1429,32'd1228,32'd3547,32'd-1695,32'd-628,32'd-1262,32'd-2937,32'd1665,32'd-118,32'd-3613,32'd-2427,32'd-886,32'd673,32'd3574,32'd-2624,32'd1278,32'd-828,32'd251,32'd150,32'd-7451,32'd3120,32'd-3552,32'd-2902,32'd52,32'd3281,32'd3049,32'd3198,32'd-240,32'd321,32'd3903,32'd435,32'd3479,32'd4104,32'd-1534,32'd447,32'd-4709,32'd2416,32'd451,32'd2912,32'd-1450,32'd-4177,32'd2727,32'd1766,32'd2868,32'd6123,32'd-564,32'd1495,32'd1695,32'd6943,32'd-5908,32'd8168,32'd6318,32'd-17,32'd3693,32'd2481,32'd-4360,32'd2432,32'd-863,32'd-589,32'd12587,32'd-5932,32'd-3989,32'd5986,32'd-6074,32'd5761,32'd-4753,32'd4265,32'd3452,32'd2644,32'd-6855,32'd2563,32'd-7622,32'd-2958,32'd2734,32'd5097,32'd3391,32'd-4497,32'd684,32'd-608,32'd3588,32'd1895,32'd-1711,32'd1530,32'd-1956,32'd60,32'd-2275,32'd1424,32'd5356,32'd-6230,32'd1000,32'd-1719,32'd6445,32'd-3666,32'd-7026,32'd-2481,32'd-1442,32'd-4946,32'd-575,32'd-4819,32'd-8481,32'd4943,32'd1614,32'd-984};
    Wh[98]='{32'd4829,32'd-2001,32'd1375,32'd-2736,32'd-1259,32'd886,32'd-8310,32'd-2558,32'd2924,32'd-1724,32'd-12343,32'd-6572,32'd-855,32'd-3244,32'd4030,32'd-5273,32'd-3767,32'd-3308,32'd-4926,32'd4675,32'd480,32'd623,32'd-3483,32'd-4853,32'd419,32'd4155,32'd-4489,32'd-103,32'd-2785,32'd3105,32'd-275,32'd-5375,32'd-4240,32'd-4833,32'd2536,32'd-2634,32'd2958,32'd-1508,32'd-8515,32'd-2658,32'd-1494,32'd-137,32'd1955,32'd-1746,32'd2792,32'd-1071,32'd-2247,32'd-5087,32'd-783,32'd1568,32'd-8383,32'd-3720,32'd-75,32'd513,32'd1611,32'd3059,32'd-492,32'd7509,32'd-755,32'd-3444,32'd4411,32'd4099,32'd-2958,32'd-3417,32'd822,32'd5312,32'd-2731,32'd-5781,32'd2792,32'd3898,32'd7,32'd-876,32'd-1932,32'd-4423,32'd-1063,32'd-6972,32'd-4741,32'd-2,32'd5292,32'd-1030,32'd-4416,32'd-1049,32'd632,32'd3332,32'd1156,32'd1434,32'd-4199,32'd1160,32'd-3674,32'd7905,32'd-1788,32'd-1408,32'd3713,32'd2912,32'd-1401,32'd-3395,32'd6450,32'd-2268,32'd-4846,32'd888,32'd-3510,32'd2436,32'd-828,32'd-4382,32'd5263,32'd266,32'd-3737,32'd3232,32'd-1773,32'd482,32'd-361,32'd3728,32'd-6811,32'd-349,32'd3300,32'd-1975,32'd-3850,32'd320,32'd1777,32'd-615,32'd4536,32'd-3454,32'd-4123,32'd-3872,32'd-5864,32'd-14453,32'd3168,32'd429,32'd4592,32'd-8066,32'd5888,32'd-3320,32'd-2030,32'd-2032,32'd3173,32'd-1771,32'd8330,32'd1789,32'd-4521,32'd78,32'd-522,32'd4340,32'd4309,32'd-552,32'd2313,32'd2451,32'd3879,32'd-2266,32'd3249,32'd2175,32'd6420,32'd2636,32'd1800,32'd-5219,32'd-1223,32'd3906,32'd8994,32'd-279,32'd-95,32'd-6191,32'd2644,32'd1452,32'd-6611,32'd-4401,32'd1210,32'd-4218,32'd-2342,32'd-3405,32'd294,32'd2495,32'd2421,32'd4096,32'd2651,32'd-1389,32'd-386,32'd-5976,32'd-4187,32'd6264,32'd-3813,32'd-1172,32'd744,32'd-2751,32'd-2080,32'd876,32'd2663,32'd2863,32'd-5551,32'd3139,32'd5092,32'd11162,32'd1890,32'd1718,32'd-4570,32'd2592,32'd-1320,32'd-5126,32'd-5004,32'd-6401,32'd419,32'd266,32'd-493,32'd6171,32'd1250,32'd1233,32'd1754,32'd1211,32'd4978,32'd668,32'd-3862,32'd316,32'd-272,32'd-2321,32'd3601,32'd3232,32'd5190,32'd-1359,32'd2050,32'd-2900,32'd-4040,32'd-1419,32'd1383,32'd-577,32'd2575,32'd7543,32'd-733,32'd6142,32'd661,32'd3559,32'd4621,32'd-2270,32'd1756,32'd-6640,32'd-4384,32'd2961,32'd-3552,32'd548,32'd-5512,32'd-1103,32'd3261,32'd-864,32'd-497,32'd-2230,32'd-5131,32'd2297,32'd1155,32'd1862,32'd5283,32'd-4291,32'd3085,32'd-2800,32'd4018,32'd1473,32'd-3815,32'd1313,32'd-5351,32'd-1635,32'd4912,32'd7397,32'd-1981,32'd4257,32'd313,32'd2077,32'd6010,32'd2744,32'd-5834,32'd4858,32'd-1711,32'd997,32'd-1033,32'd60,32'd7158,32'd8325,32'd-1914,32'd1060,32'd-2702,32'd4531,32'd3779,32'd1507,32'd-1811,32'd765,32'd-4392,32'd-5322,32'd2109,32'd-5371,32'd-2448,32'd1185,32'd-2917,32'd1071,32'd2175,32'd3525,32'd1643,32'd3664,32'd2309,32'd717,32'd152,32'd3388,32'd-961,32'd-191,32'd5566,32'd-3735,32'd-795,32'd1813,32'd-3076,32'd971,32'd-1323,32'd-3347,32'd2163,32'd-8222,32'd-282,32'd-2036,32'd2553,32'd-4672,32'd905,32'd-3754,32'd11054,32'd-3593,32'd4223,32'd-885,32'd559,32'd-992,32'd1004,32'd-2766,32'd-241,32'd348,32'd-1156,32'd2442,32'd2646,32'd-650,32'd4531,32'd-853,32'd-2236,32'd5317,32'd-183,32'd820,32'd1293,32'd2381,32'd-3208,32'd-1729,32'd-905,32'd3444,32'd1409,32'd-2578,32'd3034,32'd-5996,32'd5268,32'd-3198,32'd6567,32'd217,32'd8295,32'd-2658,32'd-3867,32'd2214,32'd-6694,32'd-1668,32'd994,32'd903,32'd1868,32'd3510,32'd-2421,32'd-1599,32'd2241,32'd1096,32'd1171,32'd517,32'd2238,32'd6186,32'd-2802,32'd4091,32'd3771,32'd-2397,32'd-5307,32'd1211,32'd-858,32'd-529,32'd-4382,32'd-4714,32'd3767,32'd1193,32'd689,32'd4223,32'd-1634,32'd-1520,32'd5351,32'd-8457,32'd-1907,32'd9252,32'd-5234,32'd2868,32'd1418,32'd2866,32'd1784,32'd-2766,32'd3239,32'd-6562,32'd-1049,32'd-3918,32'd-438,32'd-4501,32'd2215,32'd-687};
    Wh[99]='{32'd2485,32'd-4499,32'd272,32'd-1187,32'd-1330,32'd976,32'd-268,32'd-75,32'd-7495,32'd456,32'd4,32'd-4267,32'd-4423,32'd4475,32'd-2697,32'd659,32'd-3386,32'd378,32'd-4489,32'd2929,32'd-960,32'd-1336,32'd-2641,32'd-26,32'd157,32'd2225,32'd-5263,32'd-1008,32'd-1827,32'd-9218,32'd3095,32'd1143,32'd-2150,32'd1105,32'd3867,32'd2283,32'd-3730,32'd2398,32'd1427,32'd-5112,32'd-2714,32'd-1105,32'd1981,32'd-5717,32'd2115,32'd-3017,32'd-3,32'd-5087,32'd-5517,32'd391,32'd-1262,32'd-2937,32'd-1800,32'd1972,32'd3537,32'd-311,32'd-4816,32'd5366,32'd-1511,32'd2807,32'd1446,32'd903,32'd-3222,32'd-1370,32'd-906,32'd7036,32'd137,32'd899,32'd3271,32'd-2600,32'd-2814,32'd-1978,32'd-5712,32'd-4089,32'd-2191,32'd-6391,32'd917,32'd-1270,32'd-949,32'd-1221,32'd1184,32'd2303,32'd5058,32'd-4377,32'd2414,32'd4431,32'd-3486,32'd4479,32'd-988,32'd-85,32'd-1348,32'd1002,32'd764,32'd323,32'd-1246,32'd-4042,32'd3154,32'd-1580,32'd-168,32'd-5830,32'd-10292,32'd-798,32'd-1522,32'd7939,32'd5810,32'd1793,32'd-1988,32'd5336,32'd-348,32'd-3757,32'd-3244,32'd1379,32'd-5371,32'd1205,32'd2414,32'd-2932,32'd-309,32'd-729,32'd-2205,32'd5400,32'd2489,32'd3347,32'd-2587,32'd-4199,32'd-1571,32'd-7436,32'd8017,32'd1119,32'd3383,32'd-418,32'd-979,32'd1693,32'd2158,32'd-797,32'd2592,32'd-256,32'd1403,32'd-1802,32'd-469,32'd-70,32'd-4658,32'd1319,32'd5942,32'd1492,32'd-925,32'd3068,32'd577,32'd-4494,32'd1330,32'd-7749,32'd795,32'd5029,32'd-7451,32'd-2268,32'd-4995,32'd-4143,32'd-3122,32'd-1905,32'd1992,32'd-3334,32'd-2214,32'd1054,32'd1716,32'd-1061,32'd5727,32'd2196,32'd2445,32'd-5507,32'd-754,32'd-3395,32'd-5024,32'd2587,32'd-12353,32'd-4990,32'd6723,32'd-2302,32'd-3613,32'd-2709,32'd-4475,32'd-397,32'd6132,32'd-2320,32'd-5107,32'd888,32'd-903,32'd1286,32'd-1245,32'd-7407,32'd-4184,32'd3322,32'd512,32'd1486,32'd1049,32'd802,32'd2819,32'd-4721,32'd4304,32'd899,32'd6303,32'd-2626,32'd-2064,32'd-1428,32'd5249,32'd-4199,32'd-3437,32'd534,32'd-452,32'd159,32'd-1752,32'd-897,32'd-3090,32'd-5659,32'd4443,32'd-1246,32'd1455,32'd-44,32'd2731,32'd-420,32'd-946,32'd-2761,32'd-273,32'd-3457,32'd-1329,32'd1596,32'd-588,32'd-3537,32'd-2939,32'd-3603,32'd-3186,32'd-1463,32'd1910,32'd-3969,32'd565,32'd-944,32'd-1184,32'd3911,32'd990,32'd-2504,32'd1676,32'd-3530,32'd512,32'd3354,32'd1105,32'd-2702,32'd-3037,32'd-3796,32'd-4184,32'd-1041,32'd-1621,32'd1588,32'd-3200,32'd-136,32'd5214,32'd-3796,32'd1771,32'd-3249,32'd28,32'd6103,32'd-3132,32'd-1439,32'd-2218,32'd-1920,32'd-3151,32'd1013,32'd179,32'd-2822,32'd-5634,32'd-5698,32'd-2305,32'd921,32'd413,32'd5874,32'd-2366,32'd1126,32'd-1805,32'd-235,32'd-1837,32'd-437,32'd2971,32'd-4221,32'd-1188,32'd241,32'd-3835,32'd-8378,32'd-5766,32'd-7998,32'd-2968,32'd-7968,32'd-3791,32'd1888,32'd-1510,32'd-10419,32'd-2354,32'd-427,32'd6645,32'd-1700,32'd-2543,32'd-1080,32'd101,32'd-1423,32'd-4890,32'd626,32'd5932,32'd-2780,32'd225,32'd-1505,32'd-2402,32'd-2119,32'd853,32'd-4565,32'd3991,32'd-5483,32'd2299,32'd-5322,32'd-5341,32'd-502,32'd1737,32'd-390,32'd-3334,32'd-1877,32'd-1098,32'd2220,32'd1043,32'd4406,32'd203,32'd-2322,32'd-2805,32'd-2158,32'd4272,32'd-792,32'd317,32'd-1834,32'd-4252,32'd-1340,32'd2883,32'd1503,32'd-1357,32'd-6733,32'd773,32'd1729,32'd-2661,32'd-711,32'd1555,32'd-2971,32'd1604,32'd677,32'd2695,32'd-6586,32'd3354,32'd2156,32'd1069,32'd-9174,32'd-3886,32'd1231,32'd4924,32'd7866,32'd1040,32'd7080,32'd5747,32'd2712,32'd-3249,32'd-588,32'd-3654,32'd-2807,32'd3933,32'd-8657,32'd-2768,32'd2247,32'd2012,32'd-1687,32'd-2612,32'd3596,32'd-3449,32'd-4724,32'd-4130,32'd1898,32'd4875,32'd317,32'd1350,32'd1716,32'd-3583,32'd-2159,32'd-252,32'd-5664,32'd-2050,32'd6713,32'd-2541,32'd-5634,32'd-7011,32'd-3852,32'd4138,32'd2272,32'd2739,32'd1417,32'd5932,32'd2758,32'd1944,32'd-158,32'd597,32'd-1636};

    #10$display("EOF");
    #10$finish;
    end
    endmodule
    